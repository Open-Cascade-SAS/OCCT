-- Created on: 1995-01-27
-- Created by: Marie Jose MARTZ
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class BRShell from BRepToIGES inherits BREntity from BRepToIGES

    ---Purpose: This class implements the transfer of Shape Entities from Geom
    --          To IGES. These can be :
    --            . Vertex
    --            . Edge
    --            . Wire
  

uses

    Shape                from TopoDS,
    Face                 from TopoDS,
    Shell                from TopoDS,
    IGESEntity           from IGESData,
    BREntity             from BRepToIGES    
    
is 
    
    Create 
    	returns BRShell from BRepToIGES;
    
    Create (BR : BREntity from BRepToIGES)
    	returns BRShell from BRepToIGES;    


    TransferShell (me    : in out;
                   start : Shape from TopoDS)
    	returns mutable IGESEntity from IGESData;
    ---Purpose :  Transfert an Shape entity from TopoDS to IGES
    --            This entity must be a Face or a Shell.
    --            If this Entity could not be converted, this member returns a NullEntity.


    TransferShell (me    : in out;
                   start : Shell from TopoDS)
    	returns mutable IGESEntity from IGESData;
    ---Purpose :  Transfert an Shell entity from TopoDS to IGES
    --            If this Entity could not be converted, this member returns a NullEntity.


    TransferFace (me    : in out;
                  start : Face from TopoDS)
    	returns mutable IGESEntity from IGESData;
    ---Purpose :  Transfert a Face entity from TopoDS to IGES
    --            If this Entity could not be converted, this member returns a NullEntity.


end BRShell;
