-- Created on: 1993-04-13
-- Created by: Gerard GRAS
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class SetOfSegments from Graphic2d inherits Line from Graphic2d

	---Version:

	---Purpose: The primitive SetOfSegments
        --  Warning: This primitive must be use as possible for performance
        --         improvment but is drawn with a global line attributes 
        --         for all the set. 
	--	    But when the set contains a lot of contigous segments
	--	   with a line attrib different to the default,it's
	--	   more preferable to use a SetOfPolylines for to insure
	--	   a better quality.
        --         NOTE: than the method PickedIndex() permits to known 
        --              the last picked segment in the set. 
	---References:

uses
	Drawer			from Graphic2d,
	GraphicObject		from Graphic2d,
	Length			from Quantity,
	SequenceOfShortReal	from TShort,
	FStream			from Aspect,
	IFStream		from Aspect

raises
	SegmentDefinitionError	from Graphic2d,
	OutOfRange from Standard

is
	-------------------------
	-- Category: Constructors
	-------------------------

	Create (aGraphicObject: GraphicObject from Graphic2d)
	returns mutable SetOfSegments from Graphic2d;
	---Level: Public
	---Purpose: Creates an empty set of segments in the graphic 
	--         object <aGraphicObject>.
	---Category: Constructors

	Add(me : mutable; X1, Y1, X2, Y2: Length from Quantity)
	---Level: Public
	---Purpose: Add a segment in the set 
	--	    The first point is <X1>, <Y1>.
	--	    The second point is <X2>, <Y2>.
	--  Trigger: Raises SegmentDefinitionError if the
	--          first point and the second point are identical.
	raises SegmentDefinitionError from Graphic2d;
	---Category: Update method

	Length(me) returns Integer from Standard;
	---Level: Public
	---Purpose: Returns the number of segments in the set.
	---Category: Inquiry method

	Values( me; 
            aRank: Integer from Standard;
		    X1, Y1, X2, Y2: out Length from Quantity )
	---Level: Public
	---Purpose: Returns the segment of rank <aRank> from the set.
	--  Trigger: Raises OutOfRange if <aRank> is <1 or >Length()
	raises OutOfRange from Standard;
	---Category: Inquiry method

	--------------------------
	-- Category: Draw and Pick
	--------------------------

	Draw (me : mutable; aDrawer: Drawer from Graphic2d)
	is static protected;
	---Level: Internal
	---Purpose: Draws the set of segments <me>.

    DrawElement( me : mutable; aDrawer: Drawer from Graphic2d;
                 anIndex: Integer from Standard)
        is redefined protected;
    	---Level: Internal
    	---Purpose: Draws element <anIndex> of the set <me>.

    DrawVertex( me : mutable; aDrawer: Drawer from Graphic2d;
                anIndex: Integer from Standard)
        is redefined protected;
    	---Level: Internal
    	---Purpose: Draws vertex <anIndex> of the set <me>.

	Pick (me : mutable; X, Y: ShortReal from Standard;
		aPrecision: ShortReal from Standard;
		aDrawer: Drawer from Graphic2d)
	returns Boolean from Standard
	is static protected;
	---Level: Internal
        ---Purpose: Returns Standard_True if one segment of the set <me> 
	--	    is picked, Standard_False if not.
	--  Warning: The PickIndex() method returns the rank of the picked
	--	    segment if any.

	----------------------------------------------------------------------

	Save( me; aFStream: in out FStream from Aspect ) is virtual;
--	Retrieve( me; aIFStream: in out IFStream from AIS2D ) is virtual;

fields

	myX1:	SequenceOfShortReal from TShort;
	myY1:	SequenceOfShortReal from TShort;
	myX2:	SequenceOfShortReal from TShort;
	myY2:	SequenceOfShortReal from TShort;

end SetOfSegments from Graphic2d;
