-- Created on: 1992-06-22
-- Created by: Gilles DEBARBOUILLE
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Lexicon from Units 

inherits

    TShared from MMgt 

	---Purpose: This class defines a lexicon useful to analyse and
	--          recognize the  different key words  included  in a
	--          sentence.  The lexicon is stored  in a sequence of
	--          tokens.

uses

    HAsciiString   from TCollection,
    AsciiString    from TCollection,
    TokensSequence from Units

is

    Create returns mutable Lexicon from Units;
    
    ---Level: Internal 
    
    ---Purpose: Creates an empty instance of Lexicon.
    
    Creates(me : mutable ; afilename : CString)
    
    ---Level: Internal 
    
    ---Purpose: Reads the file <afilename> to create a sequence  of tokens
    --          stored in <thesequenceoftokens>.
    
    is static;
    
    Sequence(me) returns any TokensSequence from Units
    
    ---Level: Internal 
    
    ---C++: inline
    
    ---Purpose: Returns the first item of the sequence of tokens.
    
    is static;
    
    FileName(me) returns AsciiString from TCollection
    
    ---Level: Internal 
    
    ---Purpose: Returns in a AsciiString from TCollection the name of the file.
    
    is static;
    
    UpToDate(me) returns Boolean
    
    ---Level: Internal 
    
    ---Purpose: Returns true if  the  file has not  changed  since the
    --          creation   of   the  Lexicon   object.   Returns false
    --          otherwise.

    is virtual;
    
    AddToken(me : mutable ; aword , amean : CString ; avalue : Real)
    
    ---Level: Internal 
    
    ---Purpose: Adds to the lexicon a new token with <aword>, <amean>,
    --          <avalue>  as  arguments.  If there is  already a token
    --          with   the  field  <theword>  equal    to <aword>, the
    --          existing token is updated.
    
    is static;
    
    Dump(me)
    
    ---Level: Internal 
    
    ---C++: inline
    ---Purpose: Useful for debugging.

    is virtual;
    
fields

    thefilename         : HAsciiString from TCollection;
    thetime             : Time from Standard;
    thesequenceoftokens : TokensSequence from Units;

end Lexicon;
