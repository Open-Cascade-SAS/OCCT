-- File:	Image_BilinearPixelInterpolation.cdl
-- Created:	Tue Jul 27 18:47:06 1993
-- Author:	Jean Louis FRENKEL
--		<jlf@sparc3>
---Copyright:	 Matra Datavision 1993

class BilinearPixelInterpolation from Image inherits PixelInterpolation from Image

	---Purpose: The class BilinearPixelInterpolation is used to compute a  
	--            SubPixel value on non integer Image coordinate
	--          BilinearPixelInterpolation redefined a new method to compute
	--	      a SubPixel value .
	--	    The value is the bilinear interpolation of the 
	--	      four nearest Image Pixel.
	--	    If V1, V2, V3, V4 is the value  and (X1,Y1) , (X2,Y2), 
	--              (X3,Y3), (X4,Y4) the coordinates of the four nearest 
	--		Image Pixel then first we solve :
	--		V1 = a*X1 + b*Y1 + c*X1*Y1 + d 
	--		V2 = a*X2 + b*Y2 + c*X2*Y2 + d 
	--		V3 = a*X3 + b*Y3 + c*X3*Y3 + d 
	--		V1 = a*X4 + b*Y4 + c*X4*Y4 + d 
	--
	--	      and V = a*FX + b*XY + c*FX*FY + d
	--	      is the Image SubPixel value on non integer 
	--	      coordinate (FX,FY).


uses

    Image 		from Image,
    Pixel       	from Aspect,
    ColorPixel       	from Aspect,
    IndexPixel       	from Aspect,
    DColorImage 	from Image,
    DIndexedImage 	from Image

is

    	Create returns BilinearPixelInterpolation from Image ;
	---Level: Public
    	---Purpose: Create a BilinearPixelInterpolation  object.

	Interpolate( me ; aImage   : Image from Image ;
		          FX,FY      : Real  from Standard ;
			  LowerX,LowerY,UpperX,UpperY : Integer from Standard ;
		          RetPixel : in out Pixel from Aspect ) 
		returns Boolean from Standard is redefined ;
	---Level: Public
    	---Purpose: Redefined the method to compute SubPixel's value 
	--	      on non integer Image coordinate.
	--	    LowerX,LowerY,UpperX,UpperY is the Image Min Max, it's used
	--	      to check if the SubPixel coordinate FX,FY is outside of 
	--	      image.
	--          Return True  if Interpolation Succes.
	--	    Return False if the SubPixel is out from Image.

	Interpolate( me ; aImage   : DColorImage from Image ;
		          FX,FY      : Real  from Standard ;
			  LowerX,LowerY,UpperX,UpperY : Integer from Standard ;
		          RetPixel : in out ColorPixel from Aspect ) 
		returns Boolean from Standard  is redefined;
	---Level: Public
    	---Purpose: Compute SubPixel's value on non integer Image coordinate for
	--	      DColorImage and ColorPixel.
	--	    LowerX,LowerY,UpperX,UpperY is the Image Min Max, it's used
	--	      to check if the SubPixel coordinate FX,FY is outside of 
	--	      image.
	--          Return True  if Interpolation Succes.
	--	    Return False if the SubPixel is out from Image.

	Interpolate( me ; aImage   : DIndexedImage from Image ;
		          FX,FY      : Real  from Standard ;
			  LowerX,LowerY,UpperX,UpperY : Integer from Standard ;
		          RetPixel : in out IndexPixel from Aspect ) 
		returns Boolean from Standard  is redefined;
	---Level: Public
    	---Purpose: Compute SubPixel's value on non integer Image coordinate for
	--	      DIndexedImage and IndexPixel.
	--	    LowerX,LowerY,UpperX,UpperY is the Image Min Max, it's used
	--	      to check if the SubPixel coordinate X,Y is outside of 
	--	      image.
	--          Return True  if Interpolation Succes.
	--	    Return False if the SubPixel is out from Image.

end BilinearPixelInterpolation from Image;
