-- Created on: 2003-06-04
-- Created by: Galina KULIKOVA
-- Copyright (c) 2003-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package RWStepDimTol 

	---Purpose: Packsge contains tools for parsing and formatting GD&T entities.

    uses
    	TCollection,
    	RWStepRepr, 
    	RWStepShape,
    	RWStepVisual,
    	RWStepBasic,
    	TColStd,
	StepData,
    	Interface, 
	StepDimTol,
    	MMgt

    is
    	class RWAngularityTolerance;
    	class RWCircularRunoutTolerance;
    	class RWConcentricityTolerance;
    	class RWCylindricityTolerance;
    	class RWCoaxialityTolerance;
    	class RWFlatnessTolerance;
    	class RWLineProfileTolerance;
    	class RWParallelismTolerance;
    	class RWPerpendicularityTolerance;
    	class RWPositionTolerance;
    	class RWRoundnessTolerance;
    	class RWStraightnessTolerance;
    	class RWSurfaceProfileTolerance;
    	class RWSymmetryTolerance;
    	class RWTotalRunoutTolerance;
    
    	class RWGeometricTolerance;
    	class RWGeometricToleranceRelationship;
    	class RWGeometricToleranceWithDatumReference;
    	class RWModifiedGeometricTolerance;
     
    	class RWDatum;
    	class RWDatumFeature;
    	class RWDatumReference;
    	class RWCommonDatum;
    	class RWDatumTarget;
    	class RWPlacedDatumTargetFeature;
    	
	class RWGeoTolAndGeoTolWthDatRefAndModGeoTolAndPosTol;


end RWStepDimTol;
