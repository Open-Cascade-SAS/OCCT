-- Created on: 1995-03-21
-- Created by: Laurent BOURESCHE
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Regul from ChFiDS 

	---Purpose: Storage of  a curve  and its 2 faces or surfaces of  support.

is

    Create returns Regul from ChFiDS;
    
    SetCurve(me : in out; IC : Integer from Standard)
    is static;
    
    SetS1(me     : in out; 
    	  IS1    : Integer from Standard;
	  IsFace : Boolean from Standard = Standard_True)
    is static;
	  
    SetS2(me     : in out; 
    	  IS2    : Integer from Standard;
	  IsFace : Boolean from Standard = Standard_True)
    is static;
	  
    IsSurface1(me) returns Boolean from Standard is static;

    IsSurface2(me) returns Boolean from Standard is static;
    
    Curve(me) returns Integer from Standard is static;

    S1(me) returns Integer from Standard is static;

    S2(me) returns Integer from Standard is static;

fields

    icurv : Integer from Standard;
    is1   : Integer from Standard;
    is2   : Integer from Standard;

end Regul;
