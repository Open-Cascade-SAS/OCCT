-- Created on: 1993-10-20
-- Created by: Bruno DUMORTIER
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class CompBezierCurvesToBSplineCurve from ShapeConstruct 

	---Purpose: Converts a list  of connecting Bezier Curves to  a
	--          BSplineCurve.
	--          if possible, the continuity of the BSpline will be 
	--          increased to more than C0.

uses
    Array1OfReal            from TColStd,
    SequenceOfReal          from TColStd,
    SequenceOfInteger       from TColStd,
    Array1OfInteger         from TColStd,
    Array1OfPnt             from TColgp,
    SequenceOfPnt           from TColgp,
    SequenceOfArray1OfPoles from Convert

    -------------------------------------------------------------------------
    --- Don't forget to use the method Perform before accessing the Result.
    -------------------------------------------------------------------------

raises
    ConstructionError from Standard

is
    Create ( AngularTolerance : Real = 1.0e-4 )
    returns CompBezierCurvesToBSplineCurve from ShapeConstruct;

    AddCurve( me    : in out;
              Poles : Array1OfPnt from TColgp)
    is static;


    Perform(me: in out)
    	---Purpose: Computes the algorithm.
    is static;
    
    
    Degree(me) returns Integer from Standard
    is static;
    
    NbPoles(me) returns Integer from Standard
    is static;
    
    Poles(me; Poles : in out Array1OfPnt from TColgp)
    is static;
    
    NbKnots(me) returns Integer from Standard
    is static;
    
    KnotsAndMults(me;
                  Knots : in out Array1OfReal    from TColStd;
		  Mults : in out Array1OfInteger from TColStd)
    is static;
    
    
fields
    mySequence          : SequenceOfArray1OfPoles from Convert;
    CurvePoles          : SequenceOfPnt           from TColgp;
    CurveKnots          : SequenceOfReal          from TColStd;
    KnotsMultiplicities : SequenceOfInteger       from TColStd;
    myDegree            : Integer                 from Standard;
    myAngular           : Real                    from Standard;   
    myDone              : Boolean                 from Standard;

end CompBezierCurvesToBSplineCurve;
