-- Created on: 2002-12-12
-- Created by: data exchange team
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class CurveElementEndRelease from StepFEA
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity CurveElementEndRelease

uses
    CurveElementEndCoordinateSystem from StepFEA,
    HArray1OfCurveElementEndReleasePacket from StepElement

is
    Create returns CurveElementEndRelease from StepFEA;
	---Purpose: Empty constructor

    Init (me: mutable; aCoordinateSystem: CurveElementEndCoordinateSystem from StepFEA;
                       aReleases: HArray1OfCurveElementEndReleasePacket from StepElement);
	---Purpose: Initialize all fields (own and inherited)

    CoordinateSystem (me) returns CurveElementEndCoordinateSystem from StepFEA;
	---Purpose: Returns field CoordinateSystem
    SetCoordinateSystem (me: mutable; CoordinateSystem: CurveElementEndCoordinateSystem from StepFEA);
	---Purpose: Set field CoordinateSystem

    Releases (me) returns HArray1OfCurveElementEndReleasePacket from StepElement;
	---Purpose: Returns field Releases
    SetReleases (me: mutable; Releases: HArray1OfCurveElementEndReleasePacket from StepElement);
	---Purpose: Set field Releases

fields
    theCoordinateSystem: CurveElementEndCoordinateSystem from StepFEA;
    theReleases: HArray1OfCurveElementEndReleasePacket from StepElement;

end CurveElementEndRelease;
