-- Created on: 1997-04-21
-- Created by: Denis PASCAL
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Distance from DrawDim inherits Dimension from DrawDim

	---Purpose: 

uses Face    from TopoDS,
     Display from Draw

is

    Create (plane1 : Face from TopoDS; plane2 : Face from TopoDS)
    returns mutable Distance from DrawDim;

    Create (plane1 : Face from TopoDS)
    returns mutable Distance from DrawDim;
    
    Plane1 (me) returns Face from TopoDS;
	---C++: return const&

    Plane1 (me : mutable; face : Face from TopoDS);    

    Plane2 (me) returns Face from TopoDS;
	---C++: return const&

    Plane2 (me : mutable; face : Face from TopoDS);
    
    DrawOn (me; dis : in out Display);
    
fields

    myPlane1 : Face  from TopoDS;
    myPlane2 : Face  from TopoDS;
    
end Distance;
