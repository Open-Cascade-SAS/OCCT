-- Created on: 2002-10-29
-- Created by: Michael SAZONOV
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package BinObjMgt 

---Purpose: This package defines services to manage the storage
--          grain of data produced by applications.

uses
    TDF,
    Standard,
    TCollection,
    TColStd

is

        -- Storage Relocation Table
    alias SRelocationTable is IndexedMapOfTransient from TColStd;

        -- Retrieval Relocation Table
    alias RRelocationTable is DataMapOfIntegerTransient from TColStd;

    primitive PChar;            -- pointer to Character from Standard;
    primitive PByte;            -- pointer to Byte from Standard;
    primitive PExtChar;         -- pointer to ExtCharacter from Standard;
    primitive PInteger;         -- pointer to Integer from Standard;
    primitive PReal;            -- pointer to Real from Standard;
    primitive PShortReal;       -- pointer to ShortReal from Standard;

    class Persistent;

end BinObjMgt;
