-- Created on: 2006-08-08
-- Created by: Galina KULIKOVA
-- Copyright (c) 2006-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class ShapeDivideArea from ShapeUpgrade  inherits ShapeDivide from ShapeUpgrade

	---Purpose: Divides faces from sprcified shape  by max area criterium.

uses

    Shape from TopoDS,
    FaceDivide from ShapeUpgrade

is
     Create returns ShapeDivideArea from ShapeUpgrade;
    	---Purpose:
    
    Create (S: Shape from TopoDS)
    returns ShapeDivideArea from ShapeUpgrade;
    	---Purpose: Initialize by a Shape.
	
    GetSplitFaceTool (me) returns FaceDivide from ShapeUpgrade
    is redefined protected;
    	---Purpose: Returns the tool for splitting faces. 
	

     MaxArea(me: in out) returns Real;
    ---C++: inline
    ---C++: return &
    ---Purpose:Set max area allowed for faces 	

    
fields

    myMaxArea : Real;

end ShapeDivideArea;
