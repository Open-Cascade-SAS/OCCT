-- Created on: 2008-08-15
-- Created by: Sergey ZARITCHNY <szy@opencascade.com>
-- Copyright (c) 2008-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Name_2 from PNaming inherits Persistent from Standard

	---Purpose: 
uses
   NamedShape          from PNaming,
   HArray1OfNamedShape from PNaming, 
   HAsciiString        from PCollection

is
    Create returns Name_2 from PNaming;
    
    Type      (me : mutable; T : Integer from Standard);
    ---C++: inline
    
    ShapeType (me : mutable; T : Integer from Standard);
    ---C++: inline
    
    Arguments (me :mutable ; Args : HArray1OfNamedShape from PNaming);
    ---C++: inline

    StopNamedShape (me : mutable; arg : NamedShape  from PNaming);
    ---C++: inline

    Orientation (me : mutable; Or : Integer from Standard);
    ---C++: inline
 
    Type      (me) returns Integer from Standard;
    ---C++: inline
    
    ShapeType (me) returns Integer from Standard;
    ---C++: inline

    Arguments (me) returns HArray1OfNamedShape from PNaming;
    ---C++: inline

    StopNamedShape (me) returns NamedShape  from PNaming;
     ---C++: inline

    Index(me : mutable; I : Integer from Standard);
    ---C++: inline

    Index(me) returns Integer from Standard;
    ---C++: inline

    ContextLabel   (me) returns HAsciiString from PCollection;
    ---C++: return const&
    ---C++: inline 
    
    ContextLabel   (me : mutable; theLab : HAsciiString from PCollection);
    ---C++: inline
	
    Orientation(me) returns Integer from Standard; 
    ---C++: inline

fields 

    myType         : Integer             from Standard;
    myShapeType    : Integer             from Standard;
    myArgs         : HArray1OfNamedShape from PNaming;
    myStop         : NamedShape          from PNaming;
    myIndex        : Integer             from Standard;
    myContextLabel : HAsciiString        from PCollection;
    myOrientation  : Integer             from Standard;
end Name_2;
