-- Created on: 2009-04-06
-- Created by: Sergey ZARITCHNY
-- Copyright (c) 2009-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Position from TDataXtd inherits Attribute from TDF

	---Purpose: Position of a Label

uses
    RelocationTable     from TDF,
    GUID                from Standard,
    Attribute           from TDF,
    Pnt                 from gp,
    Label               from TDF
    


is

    Set(myclass; aLabel: Label from TDF; aPos : Pnt from gp);
    ---Purpose: Create if not found the TDataXtd_Position attribute set its position to <aPos>
    
    Set (myclass; aLabel : Label from TDF)  
    ---Purpose: Find an existing, or create an empty, Position.
    --            the Position attribute is returned.
    returns Position from TDataXtd;
    
    Get(myclass; aLabel: Label from TDF; aPos : in out Pnt from gp)
    ---Purpose: Search label <aLabel) for the TDataXtd_Position attribute and get its position
    --          if found returns True
    returns Boolean from Standard;
    
    Create 
    returns Position from TDataXtd;
    
    ID(me) returns GUID from Standard
    is redefined static;
	---Purpose: Returns the ID of the attribute.
	---C++: return const &
    
    GetID(myclass) returns GUID from Standard;
	---Purpose: Returns the ID of the attribute.
	---C++: return const &


    Restore(me: mutable; anAttribute : Attribute from TDF)
    is redefined;
	---Purpose: Restores the contents from <anAttribute> into this
	--          one. It is used when aborting a transaction.
	--          
 
    -- Copy use methods
    -- ----------------

    NewEmpty(me)
    returns Attribute from TDF
    is redefined;
    ---Purpose: Returns an new empty attribute from the good end
    --          type. It is used by the copy algorithm.

    Paste(me; intoAttribute    : Attribute from TDF;
    	      aRelocTationable : RelocationTable from TDF)
    is redefined;
	---Purpose: This method is different from the "Copy" one,
	--          because it is used when copying an attribute from
	--          a source structure into a target structure. This
	--          method pastes the current attribute to the label
	--          corresponding to the insertor. The pasted
	--          attribute may be a brand new one or a new version
	--          of the previous one.


    GetPosition (me)
    ---C++: return const &
    returns Pnt from gp;
    
    SetPosition (me: mutable ; aPos : Pnt from gp);

fields

    myPosition : Pnt from gp;	
    
end Position;



