-- Created on: 1992-04-06
-- Created by: Christophe MARION
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class WiresBlock from HLRAlgo inherits TShared from MMgt

	---Purpose: A WiresBlock is a set of Blocks. It is used by the
	--          DataStructure to structure the Edges.
	--          
	--          A WiresBlock contains :
	--          
	--          * An Array  of Blocks.

uses
    Address           from Standard,
    Boolean           from Standard,
    Integer           from Standard,
    EdgesBlock        from HLRAlgo,
    Array1OfTransient from TColStd
    
is
    Create(NbWires : Integer from Standard)
	---Purpose: Create a Block of Blocks.
    returns mutable WiresBlock from HLRAlgo;

    NbWires(me) returns Integer from Standard
    is static;
    
    Set(me : mutable; I  : Integer     from Standard;
		      W  : EdgesBlock  from HLRAlgo)
    is static;		   

    Wire(me : mutable; I : Integer from Standard)
    returns any EdgesBlock from HLRAlgo
	---C++: return &
    is static;
    
    UpdateMinMax(me : mutable; TotMinMax : Address from Standard)
    is static;

    MinMax(me) returns Address from Standard
	---C++: inline
    is static;

fields
    myWires  : Array1OfTransient from TColStd;
    myMinMax : Integer           from Standard[16];

end WiresBlock;
