-- Created on: 2003-09-29
-- Created by: Alexander SOLOVYOV and Sergey LITONIN
-- Copyright (c) 2003-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SensitiveFace from MeshVS inherits SensitiveFace from Select3D

	---Purpose: This class provides custom sensitive face, which will be selected if it center is in rectangle.

uses
  EntityOwner from SelectBasics,

  Array1OfPnt from TColgp,

  TypeOfSensitivity from Select3D,
  Projector         from Select3D,

  Pnt   from gp,
  Pnt2d from gp,

  Array1OfPnt2d from TColgp,

  Box2d from Bnd

is

  Create ( theOwner    : EntityOwner from SelectBasics;
           thePoints   : Array1OfPnt from TColgp;
           theSensType : TypeOfSensitivity from Select3D = Select3D_TOS_INTERIOR )
    returns SensitiveFace from MeshVS;

  Project( me: mutable; aProjector : Projector from Select3D ) is redefined;

  Matches  ( me: mutable; XMin, YMin, XMax, YMax: Real;
             aTol: Real ) returns Boolean is redefined;

  Matches  ( me: mutable; Polyline: Array1OfPnt2d from TColgp;
              aBox:Box2d; aTol: Real ) returns Boolean is redefined;

fields
  myCentre      : Pnt   from gp is protected;
  myProjCentre  : Pnt2d from gp is protected;

end SensitiveFace;
