-- File:        Face.cdl
-- Created:     Mon Dec  4 12:02:26 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWFace from RWStepShape

	---Purpose : Read & Write Module for Face

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     Face from StepShape,
     EntityIterator from Interface

is

	Create returns RWFace;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable Face from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : Face from StepShape);

	Share(me; ent : Face from StepShape; iter : in out EntityIterator);

end RWFace;
