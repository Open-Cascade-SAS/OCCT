-- Created on: 1995-03-10
-- Created by: Laurent PAINNOT
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Polygon2D from DrawTrSurf inherits Drawable2D from Draw

    	---Purpose: Used to display a 2d polygon.
    	--          
    	--          Optional display of nodes.


uses Polygon2D   from Poly,
     Display     from Draw,
     Drawable3D  from Draw,
     Interpretor from Draw,
     OStream
is

    Create(P: Polygon2D from Poly)
    returns Polygon2D from DrawTrSurf;
    
    Polygon2D(me) returns Polygon2D from Poly;
    
    ShowNodes(me: mutable; B: Boolean);
    
    ShowNodes(me) returns Boolean;
    
    DrawOn(me; dis: in out Display);
    
    Copy(me) returns Drawable3D from Draw
    is redefined;
	---Purpose: For variable copy.


    Dump(me; S : in out OStream)
    is redefined;
	---Purpose: For variable dump.

    Whatis(me; I : in out Interpretor from Draw)
    is redefined;
	---Purpose: For variable whatis command. Set  as a result  the
	--          type of the variable.


fields

    myPolygon2D:  Polygon2D from Poly;
    myNodes:      Boolean;

end Polygon2D;
