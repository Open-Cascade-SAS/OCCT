-- File:        ShapeRepresentationRelationshipWithTransformation.cdl
-- Created:     Mon Dec  4 12:02:31 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWShapeRepresentationRelationshipWithTransformation from RWStepRepr

	---Purpose : Read & Write Module for ShapeRepresentationRelationshipWithTransformation

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     ShapeRepresentationRelationshipWithTransformation from StepRepr,
     EntityIterator from Interface

is

	Create returns RWShapeRepresentationRelationshipWithTransformation;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable ShapeRepresentationRelationshipWithTransformation from StepRepr);

	WriteStep (me; SW : in out StepWriter; ent : ShapeRepresentationRelationshipWithTransformation from StepRepr);

	Share(me; ent : ShapeRepresentationRelationshipWithTransformation from StepRepr; iter : in out EntityIterator);

end RWShapeRepresentationRelationshipWithTransformation;
