-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class UncertaintyMeasureWithUnit from StepBasic 

inherits MeasureWithUnit from StepBasic 

uses

	HAsciiString from TCollection, 
	MeasureValueMember from StepBasic,
	Unit from StepBasic
is

	Create returns mutable UncertaintyMeasureWithUnit;
	---Purpose: Returns a UncertaintyMeasureWithUnit


	Init (me : mutable;
	      aValueComponent : MeasureValueMember from StepBasic;
	      aUnitComponent : Unit from StepBasic) is redefined;

	Init (me : mutable;
	      aValueComponent : MeasureValueMember from StepBasic;
	      aUnitComponent : Unit from StepBasic;
	      aName : HAsciiString from TCollection;
	      aDescription : HAsciiString from TCollection) is virtual;

	-- Specific Methods for Field Data Access --

	SetName(me : mutable; aName : HAsciiString);
	Name (me) returns HAsciiString;
	SetDescription(me : mutable; aDescription : HAsciiString);
	Description (me) returns HAsciiString;

fields

	name : HAsciiString from TCollection;
	description : HAsciiString from TCollection;

end UncertaintyMeasureWithUnit;
