-- Created on: 2014-03-15
-- Created by: Laurent PAINNOT
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class FunctionRoot from math
     ---Purpose:
     -- This class implements the computation of a root of a function of
     -- a single variable which is near an initial guess using a minimization 
     -- algorithm.Knowledge of the derivative is required. The
     -- algorithm used is the same as in

uses Vector from math, Matrix from math, 
     FunctionWithDerivative from math,
     OStream from Standard
     
raises NotDone from StdFail

is

    Create(F: in out FunctionWithDerivative;
           Guess, Tolerance: Real;
	   NbIterations: Integer = 100)
    ---Purpose:
    -- The Newton-Raphson method is done to find the root of the function F 
    -- from the initial guess Guess.The tolerance required on
    -- the root is given by Tolerance. Iterations are stopped if
    -- the expected solution does not stay in the range A..B.
    -- The solution is found when abs(Xi - Xi-1) <= Tolerance;
    -- The maximum number of iterations allowed is given by NbIterations.

    returns FunctionRoot;

    
    Create(F: in out FunctionWithDerivative;
           Guess, Tolerance,A,B: Real;
	   NbIterations: Integer = 100)
    ---Purpose:
    -- The Newton-Raphson method is done to find the root of the function F 
    -- from the initial guess Guess.
    -- The tolerance required on the root is given by Tolerance.
    -- Iterations are stopped if the expected solution does not stay in the
    -- range A..B
    -- The solution is found when abs(Xi - Xi-1) <= Tolerance;
    -- The maximum number of iterations allowed is given by NbIterations.

    returns FunctionRoot;
    
    
    IsDone(me)
      ---Purpose: Returns true if the computations are successful, otherwise returns false.
      ---C++: inline
    returns Boolean
    is static;
    
    
    Root(me)
       ---Purpose: returns the value of the root.
       -- Exception NotDone is raised if the root was not found.
      ---C++: inline

    returns Real
    raises NotDone
    is static;


    Derivative(me)
    ---Purpose: returns the value of the derivative at the root.
    -- Exception NotDone is raised if the root was not found.
      ---C++: inline

    returns Real
    raises NotDone
    is static;
    
    
    Value(me)
    	---Purpose: returns the value of the function at the root.
    -- Exception NotDone is raised if the root was not found.
      ---C++: inline

    returns Real
    raises NotDone
    is static;
    
    
    NbIterations(me)
    	---Purpose: returns the number of iterations really done on the 
    	-- computation of the Root.
        -- Exception NotDone is raised if the root was not found.
      ---C++: inline

    returns Integer
    raises NotDone
    is static;


    Dump(me; o: in out OStream)
	---Purpose: Prints on the stream o information on the current state 
    	--          of the object.
    	--          Is used to redefine the operator <<.

    is static;
    
	
fields

Done:           Boolean;
TheRoot:        Real ;
TheError:       Real ;
TheDerivative:  Real ;
NbIter:         Integer;

end FunctionRoot;
