-- Created on: 1993-03-02
-- Created by: Philippe DAUTRY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class SweptSurface from PGeom inherits Surface from PGeom

        ---Purpose : A  swept surface  is  one that is constructed  by
        --         sweeping a curve by another curve.
        --         
	---See Also : SweptSurface from Geom.


uses Dir         from gp,
     Curve       from PGeom,
     SurfaceForm from GeomAbs, 
     Shape       from GeomAbs

is


    Initialize;
	---Purpose: Initializes the field(s) with default value(s).
    	---Level: Internal 


    Initialize(aBasisCurve: Curve from PGeom;
    	       aDirection: Dir from gp);
	---Purpose: Initialize the fields with these values.
    	---Level: Internal 


  BasisCurve (me: mutable; aBasisCurve: Curve from PGeom);
        ---Purpose : Set the value of the field basisCurve with <aBasisCurve>.
    	---Level: Internal 


  BasisCurve (me) returns Curve from PGeom;
        ---Purpose : Returns the value of the field basisCurve.
    	---Level: Internal 


  Direction (me: mutable; aDirection: Dir from gp);
        ---Purpose : Set the value of the field direction with <aDirection>.
    	---Level: Internal 


  Direction (me) returns Dir from gp;
        ---Purpose : Returns the value of the field direction.
    	---Level: Internal 


fields

  basisCurve : Curve       from PGeom   is protected;
  direction  : Dir         from gp      is protected;

end;
