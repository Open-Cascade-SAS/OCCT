-- Created by: DAUTRY Philippe
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

--      	--------------------

---Version:	0.0
--Version	Date		Purpose
--		0.0	Oct 10 1997	Creation


deferred class DeltaOnRemoval from TDF
    inherits AttributeDelta from TDF

	---Purpose: This class provides default services for an
	--          AttributeDelta on a REMOVAL action.
	--          
	--          Applying this AttributeDelta means ADDING its
	--          attribute.

uses

    Attribute from TDF

-- raises

is

    Initialize(anAtt : Attribute from TDF);
	---Purpose: Initializes a TDF_DeltaOnRemoval.

end DeltaOnRemoval;
