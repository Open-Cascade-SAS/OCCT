-- Created on: 1993-07-01
-- Created by: Jean Louis FRENKEL
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Modified: TCL G002A, 28-11-00, new method GeomCurve(...)


class Curve from GGraphic2d inherits Line from Graphic2d

	---Version:

	---Purpose: The primitive Curve

	---Keywords: Primitive, Curve
	---Warning:
	---References:

uses
	Drawer		from Graphic2d,
	Curve		from Geom2d,
	GraphicObject	from Graphic2d,
	FStream		from Aspect,
	IFStream	from Aspect
is
	--------------------------------------
	-- Category: Constructors
	--------------------------------------

	Create (aGraphicObject: GraphicObject from Graphic2d;
		aCurve: Curve from Geom2d)
	returns mutable Curve from GGraphic2d;
	---Level: Public
	---Purpose: Creates a curve.
	---Category: Constructors

	--------------------------------------
	-- Category: Inquire methods
	--------------------------------------

	GeomCurve( me ) returns Curve from Geom2d;
	---Level: Internal
	---Purpose: returns the geometric curve

	--------------------------------------
	-- Category: Draw and Pick
	--------------------------------------

	Draw (me : mutable; aDrawer: Drawer from Graphic2d)
	is static protected;
	---Level: Internal
	---Purpose: Draws the curve <me>.

	Pick (me : mutable; X, Y: ShortReal from Standard;
		aPrecision: ShortReal from Standard;
		aDrawer: Drawer from Graphic2d)
	returns Boolean from Standard is static protected;
	---Level: Internal
	---Purpose: Returns Standard_True if the curve <me> is picked,
	--	    Standard_False if not.

	----------------------------------------------------------------

	Save( me; aFStream: in out FStream from Aspect ) is virtual protected;
	Retrieve(myclass; anIFStream: in out IFStream from Aspect;
		aGraphicObject: GraphicObject from Graphic2d);

fields
	myCurve:	Curve from Geom2d;

end Curve from GGraphic2d;
