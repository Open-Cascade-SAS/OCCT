-- Created on: 1992-08-18
-- Created by: Arnaud BOUZY
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class GenRel from ExprIntrp inherits Generator from ExprIntrp

	---Purpose: Implements an interpreter for equations or system 
	--          of equations made of expressions of package Expr.

uses GeneralRelation from Expr,
    AsciiString from TCollection

raises NoSuchObject

is

    Create
    ---Purpose: Creates an empty generator
    ---Level: Advanced
    returns mutable GenRel is private;

    Create( myclass ) returns GenRel;
    
    Process(me : mutable; str : AsciiString)
    ---Purpose: Processes given string.
    ---Level: Advanced 
    is static;

    IsDone(me)
    ---Purpose: Returns false if any syntax error has occurred during 
    --          process. 
    ---Level: Advanced 
    returns Boolean
    is static;
	    
    Relation(me)
    ---Purpose: Returns relation generated. Raises an exception if 
    --          IsDone answers false.
    ---Level: Advanced 
    returns mutable GeneralRelation
    raises NoSuchObject
    is static;
    
fields

    done : Boolean;
    myRelation : GeneralRelation;
    
end GenRel;
