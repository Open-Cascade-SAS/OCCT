-- Created on: 1997-10-29
-- Created by: Roman BORISOV
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package FEmTool 

	---Purpose: Tool to Finite Element methods
	
	---Level: Advanced
uses  
    TCollection, 
    TColStd, 
    math, 
    PLib,
    GeomAbs 
is  
                   
    class  Assembly; 
      
    ---Purpose: To define Criterium (or  Energy) on finite element   
    deferred  class  ElementaryCriterion;     
    class  LinearTension;      
    class  LinearFlexion;      
    class  LinearJerk;
      
    ---Purpose: To define sparse Matrix          
    deferred  class  SparseMatrix; 
    class  ProfileMatrix;

    ---Purpose: Do define one curves with Finite Element
    class  Curve;   
    
    ---Purpose:  To  define  set  of  functions  for  calculating  matrix 
    --	         elements  of  RefMatrix  by  Gauss  integration. 
    class  ElementsOfRefMatrix; 
     
    --  instantiate  classes  
      
    ---Purpose:  To define the  table  [Freedom's degree] [Dimension,Element]
    --           which gives Index  of Freedom's degree in the
    --           assembly problem.
   
    class  AssemblyTable
    instantiates Array2 from TCollection (HArray1OfInteger from  TColStd);     
    class  HAssemblyTable   
    instantiates HArray2 from TCollection (HArray1OfInteger from  TColStd,
    	    	    	                   AssemblyTable  from  FEmTool); 
					    
    ---Purpose:  To  define  list  of  segments with  non-zero  coefficients   
    --           of constraint 
        
    class  ListOfVectors  
    instantiates  List  from  TCollection  (HArray1OfReal  from  TColStd); 

    ---Purpose:  To  define  sequence  of  constraints 
    
    class  SeqOfLinConstr  
    instantiates  Sequence  from  TCollection  (ListOfVectors  from  FEmTool); 
      
     
end FEmTool;
