-- Created on: 1998-03-23
-- Created by: # Andre LIEUTIER
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class LinearScalarConstraint from Plate
---Purpose : define on or several constraints  as linear combination of
--         the X,Y and Z components of a set of PinPointConstraint
--         
uses 
   XY from gp, 
   XYZ from gp, 
   PinpointConstraint  from  Plate,
   HArray1OfPinpointConstraint  from  Plate,
   HArray2OfXYZ from TColgp,
   Array1OfPinpointConstraint  from  Plate,
   Array2OfXYZ from TColgp,
   Array1OfXYZ from TColgp 
   
raises
    DimensionMismatch from Standard,
    OutOfRange from Standard
   
is
    Create
         returns LinearScalarConstraint;

    Create  (PPC1  :  PinpointConstraint; coeff  :  XYZ ) 
           returns LinearScalarConstraint; 

    Create  (PPC  :  Array1OfPinpointConstraint; coeff  :  Array1OfXYZ ) 
           returns LinearScalarConstraint
	   raises DimensionMismatch from Standard;
    -- PPC and coeff have to be of the same length

    Create  (PPC  :  Array1OfPinpointConstraint; coeff  :  Array2OfXYZ )
           returns LinearScalarConstraint
	   raises DimensionMismatch from Standard;
    --  the length of PPC  have to be the  Row lentgth of  coeff

    Create  (ColLen,RowLen  :  Integer ) 
    -- initialize with 0 valued PPC and Coeffs
           returns LinearScalarConstraint;

    -- Accessors :
    GetPPC(me) returns Array1OfPinpointConstraint;
    ---C++: inline 
    ---C++: return const &

    Coeff(me) returns Array2OfXYZ;
    ---C++: inline 
    ---C++: return const &

    SetPPC (me : in out;  
    	Index: Integer from Standard;  
    	Value: PinpointConstraint) 
    	---Purpose:  Sets   the PinPointConstraint of   index Index to
    	--          Value raise if Index is greater than the length of
    	--          PPC or the Row length of coeff or lower  than 1
    	raises OutOfRange from Standard;

    SetCoeff (me : in out;  
    	Row, Col: Integer from Standard;  
    	Value: XYZ) 
    	---Purpose:  Sets the coeff  of index (Row,Col)  to Value 
    	--           raise if  Row (respectively Col)  is greater than the
    	--          Row (respectively Column) length of coeff
    	raises OutOfRange from Standard;

fields
    
    myPPC  :  HArray1OfPinpointConstraint;
    myCoef :  HArray2OfXYZ;

end;
