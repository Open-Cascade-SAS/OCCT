-- Created on: 2002-12-10
-- Created by: data exchange team
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V2.0

class ElementAspect from StepElement
inherits SelectType from StepData

    ---Purpose: Representation of STEP SELECT type ElementAspect

uses
    SelectMember from StepData,
    ElementVolume from StepElement,
    CurveEdge from StepElement

is
    Create returns ElementAspect from StepElement;
	---Purpose: Empty constructor

    CaseNum (me; ent: Transient) returns Integer;
	---Purpose: Recognizes a kind of ElementAspect select type
	--          return 0 

    CaseMem (me; ent: SelectMember from StepData) returns Integer is redefined;
	---Purpose: Recognizes a items of select member ElementAspectMember
	--          1 -> ElementVolume
	--          2 -> Volume3dFace
	--          3 -> Volume2dFace
	--          4 -> Volume3dEdge
	--          5 -> Volume2dEdge
	--          6 -> Surface3dFace
	--          7 -> Surface2dFace
	--          8 -> Surface3dEdge
	--          9 -> Surface2dEdge
	--          10 -> CurveEdge
	--          0 else


     NewMember(me) returns SelectMember from StepData is redefined;
	---Purpose: Returns a new select member the type ElementAspectMember

    SetElementVolume(me: in out; aVal :ElementVolume from StepElement);
	---Purpose: Set Value for ElementVolume

    ElementVolume (me) returns ElementVolume from StepElement;
	---Purpose: Returns Value as ElementVolume (or Null if another type)

    SetVolume3dFace(me: in out; aVal :Integer);
	---Purpose: Set Value for Volume3dFace

    Volume3dFace (me) returns Integer;
	---Purpose: Returns Value as Volume3dFace (or Null if another type)

    SetVolume2dFace(me: in out; aVal :Integer);
	---Purpose: Set Value for Volume2dFace

    Volume2dFace (me) returns Integer;
	---Purpose: Returns Value as Volume2dFace (or Null if another type)

    SetVolume3dEdge(me: in out; aVal :Integer);
	---Purpose: Set Value for Volume3dEdge

    Volume3dEdge (me) returns Integer;
	---Purpose: Returns Value as Volume3dEdge (or Null if another type)

    SetVolume2dEdge(me: in out; aVal :Integer);
	---Purpose: Set Value for Volume2dEdge

    Volume2dEdge (me) returns Integer;
	---Purpose: Returns Value as Volume2dEdge (or Null if another type)

    SetSurface3dFace(me: in out; aVal :Integer);
	---Purpose: Set Value for Surface3dFace

    Surface3dFace (me) returns Integer;
	---Purpose: Returns Value as Surface3dFace (or Null if another type)

    SetSurface2dFace(me: in out; aVal :Integer);
	---Purpose: Set Value for Surface2dFace

    Surface2dFace (me) returns Integer;
	---Purpose: Returns Value as Surface2dFace (or Null if another type)

    SetSurface3dEdge(me: in out; aVal :Integer);
	---Purpose: Set Value for Surface3dEdge

    Surface3dEdge (me) returns Integer;
	---Purpose: Returns Value as Surface3dEdge (or Null if another type)

    SetSurface2dEdge(me: in out; aVal :Integer);
	---Purpose: Set Value for Surface2dEdge

    Surface2dEdge (me) returns Integer;
	---Purpose: Returns Value as Surface2dEdge (or Null if another type)

    SetCurveEdge(me: in out; aVal :CurveEdge from StepElement);
	---Purpose: Set Value for CurveEdge

    CurveEdge (me) returns CurveEdge from StepElement;
	---Purpose: Returns Value as CurveEdge (or Null if another type)

end ElementAspect;
