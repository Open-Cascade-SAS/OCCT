-- File:        ReparametrisedCompositeCurveSegment.cdl
-- Created:     Mon Dec  4 12:02:31 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWReparametrisedCompositeCurveSegment from RWStepGeom

	---Purpose : Read & Write Module for ReparametrisedCompositeCurveSegment

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     ReparametrisedCompositeCurveSegment from StepGeom,
     EntityIterator from Interface

is

	Create returns RWReparametrisedCompositeCurveSegment;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable ReparametrisedCompositeCurveSegment from StepGeom);

	WriteStep (me; SW : in out StepWriter; ent : ReparametrisedCompositeCurveSegment from StepGeom);

	Share(me; ent : ReparametrisedCompositeCurveSegment from StepGeom; iter : in out EntityIterator);

end RWReparametrisedCompositeCurveSegment;
