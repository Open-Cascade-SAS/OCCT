-- Created on: 1992-03-26
-- Created by: Herve LEGRAND
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


package GeomLProp

    ---Purpose: These global functions compute the degree of
    --          continuity of a 3D curve built by concatenation of two
    --          other curves (or portions of curves) at their junction point.

uses Standard, gp, Geom, GeomAbs, LProp

is
    
    private  class CurveTool; 
    private  class SurfaceTool;
					    
    class CLProps from GeomLProp 
            instantiates CLProps from LProp(Curve      from Geom,
	                                    Vec        from gp,
					    Pnt        from gp,
					    Dir        from gp,
					    CurveTool  from GeomLProp); 
					     

    class SLProps from GeomLProp 
            instantiates SLProps from LProp(Surface     from Geom,
	                                    SurfaceTool from GeomLProp); 

    
    Continuity(C1,C2 : Curve from Geom;
    	       u1,u2 : Real from Standard;
    	       r1,r2 : Boolean from Standard;
               tl,ta : Real from Standard) 
    ---Purpose: Computes the regularity at the junction between C1 and
    --          C2. The booleans r1 and r2 are true if the curves must
    --          be taken reversed.  The point u1 on C1 and the point
    --          u2 on C2 must be confused.
    --          tl and ta are the linear and angular tolerance used two
    --          compare the derivative.
    returns Shape from GeomAbs;

    
    Continuity(C1,C2 : Curve from Geom;
    	       u1,u2 : Real from Standard;
    	       r1,r2 : Boolean from Standard) 
    ---Purpose: The  same  as  preciding   but   using  the   standard
    --          tolerances from package Precision.
    returns Shape from GeomAbs;

end GeomLProp;    




