-- Created on: 1993-06-14
-- Created by: Martine LANGLOIS
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class MakeDirection from GeomToStep inherits Root from GeomToStep

    ---Purpose: This class implements the mapping between classes 
    --          Direction from Geom, Geom2d and Dir, Dir2d from gp, and the
    --          class Direction from StepGeom which describes a direction
    --          from Prostep. 
  
uses Dir from gp,
     Dir2d from gp,
     Direction from Geom,
     Direction from Geom2d,
     Direction from StepGeom
     
raises NotDone from StdFail
     
is 

Create ( D : Dir from gp ) returns MakeDirection;

Create ( D : Dir2d from gp ) returns MakeDirection;

Create ( D : Direction from Geom ) returns MakeDirection;

Create ( D : Direction from Geom2d ) returns MakeDirection;

Value (me) returns Direction from StepGeom
    raises NotDone
    is static;
    ---C++: return const&
    
fields

    theDirection : Direction from StepGeom;
    	-- The solution from StepGeom
    	
end MakeDirection;


