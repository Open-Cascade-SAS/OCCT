-- Created on: 1997-03-28
-- Created by: Christian CAILLET
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MeasureValueMember  from StepBasic    inherits  SelectReal  from StepData

    ---Purpose : for Select MeasureValue, i.e. :
    --         length_measure,time_measure,plane_angle_measure,
    --         solid_angle_measure,ratio_measure,parameter_value,
    --         context_dependent_measure,positive_length_measure,
    --         positive_plane_angle_measure,positive_ratio_measure,
    --	       area_measure,volume_measure

uses CString

is

    Create returns mutable MeasureValueMember;
    -- starts as case null (no name)

    HasName (me) returns Boolean  is redefined;
    -- returns True is case not null

    Name    (me) returns CString  is redefined;
    --  returns a name according to the case
    --  0 -> void
    --  1 -> LENGTH_MEASURE
    --  2 -> TIME_MEASURE
    --  3 -> PLANE_ANGLE_MEASURE
    --  4 -> SOLID_ANGLE_MEASURE
    --  5 -> RATIO_MEASURE
    --  6 -> PARAMETER_VALUE
    --  7 -> CONTEXT_DEPENDANT_MEASURE
    --  8 -> POSITIVE_LENGTH_MEASURE
    --  9 -> POSITIVE_PLANE_ANGLE_MEASURE
    --  10 -> POSITIVE_RATIO_MEASURE
    --  11 -> AREA_MEASURE
    --  12 ->VOLUME_MEASURE
    --  13 ->MASS_MEASURE
    --  14 ->THERMODYNAMIC_TEMPERATURE_MEASURE
    
    SetName (me : mutable; name : CString)  returns Boolean  is redefined;
    -- checks for one of the names above, and sets the case number
    -- accepts a void name (case 0)

fields

    thecase : Integer;

end MeasureValueMember;
