-- File:    QATelco_MyText.cdl
-- Created: Wed Apr 10 10:30:17 2002
-- Author:  QA Admin
--      <qa@umnox.nnov.matra-dtv.fr>
---Copyright:    Matra Datavision 2002

class  MyText  from  QATelco  inherits  InteractiveObject  from  AIS 
uses 
    ExtendedString from TCollection, 
    Pnt from gp, 
    PresentationManager3d from PrsMgr, 
    Presentation from Prs3d,
    NameOfColor  from  Quantity,
    Selection from SelectMgr
is 
    Create(aText  :ExtendedString  from  TCollection;aPosition  : Pnt  from  gp)
    returns mutable MyText from QATelco;
    Create(aText  :ExtendedString  from  TCollection;aPosition  : Pnt  from  gp;aFont :  CString from Standard; aColor : NameOfColor  from  Quantity; aHeight :Real  from  Standard)
    returns mutable MyText from QATelco;

    NbPossibleSelection(me)
    returns Integer from Standard
    is redefined virtual protected;
    
    Compute(me:mutable;
            aPresentationManager: PresentationManager3d from PrsMgr;
            aPresentation: mutable Presentation from Prs3d;
            aMode: Integer from Standard = 0)
    is redefined virtual protected;

    ComputeSelection(me:mutable; aSelection :mutable Selection from SelectMgr;
                                 aMode      : Integer) is redefined virtual protected;

fields
        myPosition                   : Pnt from gp;
        myText                       : ExtendedString from TCollection;
        myNameOfColor                : NameOfColor from Quantity;
        myNameOfFont                 : CString from Standard;
        myHeight                     : Real from Standard;
end MyText;
    
