-- Created on: 1999-10-14
-- Created by: VKH
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Updated:     GG IMP100701 Add the "depth" field and method
--              to the pixmap object.

class PixMap from Xw

    ---Version:

    ---Purpose: This class defines a X11 pixmap

    ---Keywords: Bitmap, Pixmap, X11

inherits
    Transient             from Standard
uses
    Handle                from Aspect,
    Color                 from Quantity,
    Window                from Aspect,
    Window                from Xw
raises
    PixmapDefinitionError from Aspect,
    PixmapError           from Aspect
is
    Create ( aWindow          : Window from Aspect;
             aWidth, anHeight : Integer from Standard;
             aDepth           : Integer from Standard = 0 )
    returns mutable PixMap from Xw
    raises PixmapDefinitionError from Aspect;
    ---Level: Public
    ---Purpose:  Warning! When <aDepth> is NULL , the pixmap is created
    -- with the SAME depth than the window <aWindow>

    ---------------------------------------------------
    -- Category: Methods to modify the class definition
    ---------------------------------------------------

    Destroy ( me : mutable )
    ---Level: Advanced
    ---Purpose: Destroies the Pixmap
    --  Trigger: Raises if Pixmap is not defined properly
    raises PixmapError from Aspect is virtual;

    Dump ( me ; aFilename : CString from Standard;
           aGammaValue: Real from Standard = 1.0 )
    returns Boolean
    is virtual;
    ---Level: Advanced
    ---Purpose:
    -- Dumps the Bitmap to an image file with
    -- an optional gamma correction value
    -- and returns TRUE if the dump occurs normaly.
    ---Category: Methods to modify the class definition

    PixelColor ( me         : in;
                 theX, theY : in Integer from Standard )
    returns Color from Quantity
    is virtual;
    ---Purpose:
    -- Returns the pixel color.

    ----------------------------
    -- Category: Inquire methods
    ----------------------------

    PixmapID ( me ) returns Handle from Aspect is virtual;
    ---Level: Advanced
    ---Purpose: Returns the ID of the just created pixmap
    ---Category: Inquire methods

    ----------------------------
    -- Category: Private methods
    ----------------------------

    PreferedDepth( me ; aWindow : Window from Aspect;
                   aDepth : Integer from Standard)
    returns Integer from Standard is private;

fields
    myPixmap : Handle from Aspect is protected;
    myWindow : Window from Xw;
    myWidth  : Integer from Standard is protected;
    myHeight : Integer from Standard is protected;
    myDepth	 : Integer from Standard is protected;
end PixMap;
