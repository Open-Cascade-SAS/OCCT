-- Created on: 1996-02-16
-- Created by: Philippe MANGIN
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Batten from DrawFairCurve inherits  BSplineCurve2d from DrawTrSurf

	---Purpose: Interactive Draw object of type "Batten"

uses Batten from FairCurve, 
     BSplineCurve2d from DrawTrSurf,
     Pnt2d from gp

is
   Create(TheBatten : Address)
   returns mutable Batten from DrawFairCurve;
   Compute(me:mutable);
   SetPoint(me: mutable; Side : Integer; Point : Pnt2d);
   SetAngle(me: mutable; Side : Integer; Angle : Real);
   SetSliding(me: mutable; Length : Real);
   SetHeight(me: mutable; Heigth : Real);
   SetSlope(me: mutable; Slope : Real);
   GetAngle(me; Side : Integer) returns Real;
   GetSliding(me) returns Real;
   FreeSliding(me:mutable);
   FreeAngle(me:mutable; Side : Integer);
   Dump(me; S : in out OStream)
	---Purpose: For variable dump.
  is redefined;
   
fields
 MyBatten : Address is protected;
end Batten;
