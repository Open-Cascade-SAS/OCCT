-- Created on: 1992-05-22
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

generic class IntCurveCurveGen from IntCurve (
    TheCurve         as any;
    TheCurveTool     as any) -- as CurveTool from IntCurve(TheCurve)

	---Purpose: Provides the algorithm to intersect two 2D-curves.
	--          The curves may be parametric curves or Conic (see
	--          the template class CurveTool).
	--
	-- Note: The  exception  ConstructionError  is   raised  in
	--          constructors  or in Perform  methods when a domain
	--          (Domain from IntRes2d)  is not  correct, i-e  when
	--          the method  TheType  returns GeomAbs_Circle     or
	--          GeomAbs_Ellipsei   and the corresponding domain is
	--          not  closed (use the SetEquivalentParameters for a
	--          domain on  a circle  or an  ellipse)  or  when the
	--          method  TheType   returns  GeomAbs_Other and   the
	--          domain     of  the   curve   is    not     bounded
	--          (HasFirstPoint() && HasLastPoint() return True).
        ---Level: Advanced
        
inherits Intersection from IntRes2d

uses Domain        from IntRes2d,
     IntConicConic from IntCurve,
     IConicTool    from IntCurve,
     Array1OfReal  from TColStd
 
raises ConstructionError from Standard

		      
    	class TheProjPCur instantiates ProjPCurGen from IntCurve(
	    	        TheCurve,
    	    	        TheCurveTool);
		       
        class TheIntConicCurve instantiates IntConicCurveGen from IntCurve
	                (IConicTool      from  IntCurve,
                         TheCurve,
			 TheCurveTool,
                         TheProjPCur);

        class IntConicCurve instantiates UserIntConicCurveGen from IntCurve
	                (IConicTool      from  IntCurve,
                         TheCurve,
			 TheCurveTool,
                         TheIntConicCurve);

    	class TheIntPCurvePCurve  instantiates IntPolyPolyGen from IntCurve
	                (TheCurve,
			 TheCurveTool,
                         TheProjPCur);
is

    Create
    
	---Purpose: Empty constructor.
    	returns IntCurveCurveGen from IntCurve;
    	---C++: inline


    Create (C:  TheCurve; TolConf,Tol: Real from Standard)
    
    	---Purpose: Self Intersection of a curve
    	---C++: inline
    	returns IntCurveCurveGen from IntCurve
	raises ConstructionError from Standard;


    Create (C:  TheCurve; D: Domain from IntRes2d;
    	    TolConf,Tol: Real from Standard)
	    
        ---Purpose: Self Intersection of a curve with a domain.
    	---C++: inline
    	returns IntCurveCurveGen from IntCurve
	raises ConstructionError from Standard;
	    

    Create (C1:  TheCurve; C2:  TheCurve;
    	    TolConf,Tol: Real from Standard)

	---Purpose: Intersection between 2 curves.
    	---C++: inline 
    	returns IntCurveCurveGen from IntCurve
	raises ConstructionError from Standard;


    Create (C1:  TheCurve; D1: Domain from IntRes2d;
            C2:  TheCurve; 
    	    TolConf,Tol: Real from Standard)

	---Purpose: Intersection between 2 curves.
    	---C++: inline
    	returns IntCurveCurveGen from IntCurve
	raises ConstructionError from Standard;
	
	
    Create (C1:  TheCurve; 
            C2:  TheCurve; D2: Domain from IntRes2d;
    	    TolConf,Tol: Real from Standard)
    
	---Purpose: Intersection between 2 curves.
    	---C++: inline
    	returns IntCurveCurveGen from IntCurve
	raises ConstructionError from Standard;



    Create (C1:  TheCurve; D1: Domain from IntRes2d;
            C2:  TheCurve; D2: Domain from IntRes2d;
    	    TolConf,Tol: Real from Standard)

	---Purpose: Intersection between 2 curves.
    	---C++: inline
    	returns IntCurveCurveGen from IntCurve
	raises ConstructionError from Standard;



    Perform (me: in out;
             C1:  TheCurve; D1: Domain from IntRes2d;
             C2:  TheCurve; D2: Domain from IntRes2d;
    	     TolConf,Tol: Real from Standard)
	---Purpose: Intersection between 2 curves.

    	raises ConstructionError from Standard
    	is static;

    Perform (me: in out;
             C1:  TheCurve; 
             C2:  TheCurve; 
    	     TolConf,Tol: Real from Standard)
    	
	---Purpose: Intersection between 2 curves.
    	---C++: inline
    	raises ConstructionError from Standard
    	is static;

    Perform (me: in out;
             C1:  TheCurve; D1: Domain from IntRes2d;
    	     TolConf,Tol: Real from Standard)

	---Purpose: Intersection between 2 curves.
    	raises ConstructionError from Standard
    	is static;

    Perform (me: in out;
             C1:  TheCurve; 
    	     TolConf,Tol: Real from Standard)

	---Purpose: Intersection between 2 curves.

    	raises ConstructionError from Standard
    	is static;

    Perform (me: in out;
             C1:  TheCurve; D1: Domain from IntRes2d;
             C2:  TheCurve; 
    	     TolConf,Tol: Real from Standard)
    	---C++: inline
	---Purpose: Intersection between 2 curves.

    	raises ConstructionError from Standard
    	is static;

    Perform (me: in out;
             C1:  TheCurve; 
             C2:  TheCurve; D2: Domain from IntRes2d;
    	     TolConf,Tol: Real from Standard)
    	---C++: inline
	---Purpose: Intersection between 2 curves.

    	raises ConstructionError from Standard
    	is static;


    ComputeDomain(me;  C1: TheCurve; TolDomain: Real from Standard)
    
    	---Purpose: Create a domain from a curve
        returns Domain from IntRes2d
        is static;
	
    
    
    InternalPerform(me: in out;
             C1:  TheCurve; D1: Domain from IntRes2d;
             C2:  TheCurve; D2: Domain from IntRes2d;
    	     TolConf,Tol: Real from Standard;
    	     Composite: Boolean from Standard)

	---Purpose: Intersection between 2 curves.

    	raises ConstructionError from Standard
    	is static private;
	
	
	
    InternalCompositePerform_noRecurs(me: in out;
    	    NbInterC1: Integer from Standard;
	    C1:  TheCurve;
    	    NumInterC1: Integer from Standard;
	    Tab1: Array1OfReal from TColStd;
            D1: Domain from IntRes2d;          
	    NbInterC2: Integer from Standard;
	    C2:  TheCurve;
	    NumInterC2: Integer from Standard;
	    Tab2: Array1OfReal from TColStd;
	    D2: Domain from IntRes2d;
    	    TolConf,Tol: Real from Standard)
	
     	---Purpose: Part of InternalCompositePerform function
     
     	raises ConstructionError from Standard
    	is static private;
    	
  

    InternalCompositePerform(me: in out;
             C1:  TheCurve; D1: Domain from IntRes2d;
	     N1,NB1: Integer from Standard;
	     Tab1: Array1OfReal from TColStd;
             C2:  TheCurve; D2: Domain from IntRes2d;
	     N2,NB2: Integer from Standard;
	     Tab2: Array1OfReal from TColStd;
    	     TolConf,Tol: Real from Standard;
    	     Composite: Boolean from Standard)

	---Purpose: Intersection between 2 curves.

    	raises ConstructionError from Standard
    	is static private;


fields

    param1inf     : Real              from Standard;
    param1sup     : Real              from Standard;
    param2inf     : Real              from Standard;
    param2sup     : Real              from Standard;
    intconiconi   : IntConicConic     from IntCurve;
    intconicurv   : TheIntConicCurve;
    intcurvcurv   : TheIntPCurvePCurve;

end IntCurveCurveGen;





