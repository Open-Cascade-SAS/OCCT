-- Created on: 1993-01-11
-- Created by: CKY / Contract Toubro-Larsen ( Kiran )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package IGESGeom


        ---Purpose : This package consists of B-Rep and CSG Solid entities

uses

        Standard,
        TCollection,
	TColgp,
	TColStd,
        gp,
	Message,
        Interface,
        IGESBasic,
        IGESData

is

        class CircularArc;

        class CompositeCurve;

        class ConicArc;

        class CopiousData;

        class Plane;

        class Line;

        class SplineCurve;

        class SplineSurface;

        class Point;

        class RuledSurface;

        class SurfaceOfRevolution;

        class TabulatedCylinder;

        class Direction;

        class TransformationMatrix;

        class Flash;

        class BSplineCurve;

        class BSplineSurface;

        class OffsetCurve;

        class OffsetSurface;

        class Boundary;

        class CurveOnSurface;

        class BoundedSurface;

        class TrimmedSurface;

    	--    Tools for Entities    --

        class ToolCircularArc;
        class ToolCompositeCurve;
        class ToolConicArc;
        class ToolCopiousData;
        class ToolPlane;
        class ToolLine;
        class ToolSplineCurve;
        class ToolSplineSurface;
        class ToolPoint;
        class ToolRuledSurface;
        class ToolSurfaceOfRevolution;
        class ToolTabulatedCylinder;
        class ToolDirection;
        class ToolTransformationMatrix;
        class ToolFlash;
        class ToolBSplineCurve;
        class ToolBSplineSurface;
        class ToolOffsetCurve;
        class ToolOffsetSurface;
        class ToolBoundary;
        class ToolCurveOnSurface;
        class ToolBoundedSurface;
        class ToolTrimmedSurface;

    -- Definition and Exploitation of Entities defined in this Package

    class Protocol;
    class ReadWriteModule;
    class GeneralModule;
    class SpecificModule;

    -- Instantiations :

    class  Array1OfBoundary instantiates  Array1 from TCollection (Boundary);
    class  Array1OfCurveOnSurface        instantiates
	  Array1 from TCollection (CurveOnSurface);
    class  Array1OfTransformationMatrix  instantiates
    	  Array1 from TCollection (TransformationMatrix);

    class HArray1OfBoundary instantiates HArray1 from TCollection
    	 (Boundary,Array1OfBoundary);
    class HArray1OfCurveOnSurface        instantiates HArray1 from TCollection
    	 (CurveOnSurface,Array1OfCurveOnSurface);
    class HArray1OfTransformationMatrix  instantiates HArray1 from TCollection
    	 (TransformationMatrix,Array1OfTransformationMatrix);

    -- Package Methods

    Init;
    ---Purpose : Prepares dymanic data (Protocol, Modules) for this package

    Protocol  returns Protocol from IGESGeom;
    ---Purpose : Returns the Protocol for this Package

end IGESGeom;
