-- Created on: 1998-10-29
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Hctxee2d from TopOpeBRep inherits TShared from  MMgt

uses

    Shape from TopoDS,
    Edge from TopoDS,
    Surface from BRepAdaptor,
    Face from TopoDS,
    Curve from Geom2dAdaptor,
    CurveType from GeomAbs,
    Domain from IntRes2d
    
is

    Create returns Hctxee2d from TopOpeBRep;
    SetEdges(me:mutable;E1,E2:Edge;BAS1,BAS2:Surface from BRepAdaptor);
    Edge(me;I:Integer) returns Shape;---C++ : return const &
    Curve(me;I:Integer) returns Curve from Geom2dAdaptor; ---C++ : return const &
    Domain(me;I:Integer) returns Domain from IntRes2d; ---C++ : return const &

fields

    myEdge1 : Edge from TopoDS;
    myCurve1 : Curve from Geom2dAdaptor;
    myDomain1 : Domain from IntRes2d;

    myEdge2 : Edge from TopoDS;
    myCurve2 : Curve from Geom2dAdaptor;
    myDomain2 : Domain from IntRes2d;

end Hctxee2d from TopOpeBRep;
