-- Created by: Peter KURNEV
-- Copyright (c) 2010-2012 OPEN CASCADE SAS
-- Copyright (c) 2007-2010 CEA/DEN, EDF R&D, OPEN CASCADE
-- Copyright (c) 2003-2007 OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN, CEDRAT,
--                         EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

deferred class BuilderArea from BOPAlgo 
    	inherits Algo from BOPAlgo 
	 
	---Purpose: The root class for algorithms to build  
    	--          faces/solids from set of edges/faces  

uses 
    Shape from TopoDS, 
    BaseAllocator from BOPCol, 
    ListOfShape from BOPCol,
    MapOfOrientedShape from BOPCol, 
    Context  from BOPInt 
    
--raises

is 
    Initialize  
    	returns BuilderArea from BOPAlgo; 
    ---C++: alias "Standard_EXPORT virtual ~BOPAlgo_BuilderArea();"  
     
    Initialize(theAllocator: BaseAllocator from BOPCol)   
    	returns BuilderArea from BOPAlgo; 
     
    SetContext(me:out; 
    	    theContext:Context from BOPInt);  
    	
    Shapes(me) 
    	returns ListOfShape from BOPCol;   
    ---C++:  return const &   
    ---C++: alias "Standard_EXPORT void SetShapes(const BOPCol_ListOfShape& theLS);"  
    
    Loops(me)  
    	returns ListOfShape from BOPCol; 
    ---C++:  return const &   
     
    Areas(me) 
    	returns ListOfShape from BOPCol; 
    ---C++:  return const &     
     
    PerformShapesToAvoid(me:out) 
    	is deferred protected; 
	 
    PerformLoops(me:out) 
    	is deferred protected;  
	 
    PerformAreas(me:out)   
    	is deferred protected;  

    PerformInternalShapes(me:out)   
    	is deferred protected;  

fields  
    myContext        :  Context from BOPInt is protected; 
    myShapes         :  ListOfShape from BOPCol is protected;  
    myLoops          :  ListOfShape from BOPCol is protected;  
    myLoopsInternal  :  ListOfShape from BOPCol is protected;
    
    myAreas          :  ListOfShape from BOPCol is protected;  
    myShapesToAvoid  :  MapOfOrientedShape from BOPCol is protected;  
    --
       	 

end BuilderArea; 

