-- File:	DNaming_Line3DDriver.cdl
-- Created:	Fri Feb 26 15:51:03 2010
-- Author:	Sergey ZARITCHNY <sergey.zaritchny@opencascade.com> 
--		<szy@petrox.nnov.matra-dtv.fr>
---Copyright:	Open CasCade SA 2010 

class Line3DDriver from DNaming inherits Driver from TFunction

	---Purpose: Computes Line 3D function

uses
     Label            from TDF, 
     Logbook          from TFunction,
     Function         from TFunction,
     Wire             from TopoDS,
     Array1OfShape    from TopTools
is
  Create returns mutable Line3DDriver from DNaming;
    ---Purpose: Constructor

    ---Purpose: validation
    --          ==========

    Validate(me; theLog : in out Logbook from TFunction)
    is redefined;
    ---Purpose: Validates labels of a function in <log>.
    --          In regeneration mode this method must be called (by the
    --          solver) even if the function is not executed, to build
    --          the valid label scope.

    ---Purpose: execution of function
    --          ======================

    MustExecute (me; theLog : Logbook from TFunction)
    ---Purpose: Analyse in <log> if the loaded function must be executed
    --          (i.e.arguments are modified) or not.
    --          If the Function label itself is modified, the function must
    --          be executed.
    returns Boolean from Standard
    is redefined;

    Execute (me; theLog : in out Logbook from TFunction)
    ---Purpose: Execute the function and push in <log> the impacted
    --          labels (see method SetImpacted).
    returns Integer from Standard
    is redefined;
      
    LoadNamingDS(me; theResultLabel : Label from TDF; theWire :  Wire from TopoDS;  
    	    	     theVertexes :  Array1OfShape from TopTools; 
    	    	     isClosed : Boolean from Standard = Standard_False)  is private; 
    ---Purpose: Loads a Line3D in a data framework  
    
end Line3DDriver;

