-- Created on: 1994-02-21
-- Created by: Laurent PAINNOT
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MCurvesToBSpCurve from Approx



uses MultiBSpCurve        from AppParCurves,
     MultiCurve           from AppParCurves,
     SequenceOfMultiCurve from AppParCurves

is


    Create returns MCurvesToBSpCurve;
    
    Reset(me: in out) 
    	--- Clear the internal Sequence Of MultiCurve
    is static;
    
    Append(me: in out; MC: MultiCurve from AppParCurves)
    is static;


    Perform(me: in out)
    is static;
    
    Perform(me: in out; TheSeq: SequenceOfMultiCurve from AppParCurves)
    is static;
    
    
    Value(me)
    	---Purpose: return the composite MultiCurves as a MultiBSpCurve.
    	---C++: return const&

    returns MultiBSpCurve
    is static;


    ChangeValue(me: in out)
    	---Purpose: return the composite MultiCurves as a MultiBSpCurve.
    	---C++: return const&

    returns MultiBSpCurve
    is static;


fields


mySpline: MultiBSpCurve           from AppParCurves;
myDone  : Boolean                 from Standard;
myCurves: SequenceOfMultiCurve    from AppParCurves; 

end MCurvesToBSpCurve;
