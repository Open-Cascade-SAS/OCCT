-- Created on: 1999-11-26
-- Created by: Andrey BETENEV
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0

class SurfaceBoundary from StepGeom
inherits SelectType from StepData

    ---Purpose: Representation of STEP SELECT type SurfaceBoundary

uses
    BoundaryCurve from StepGeom,
    DegeneratePcurve from StepGeom

is
    Create returns SurfaceBoundary from StepGeom;
	---Purpose: Empty constructor

    CaseNum (me; ent: Transient) returns Integer;
	---Purpose: Recognizes a kind of SurfaceBoundary select type
	--          1 -> BoundaryCurve from StepGeom
	--          2 -> DegeneratePcurve from StepGeom
	--          0 else

    BoundaryCurve (me) returns BoundaryCurve from StepGeom;
	---Purpose: Returns Value as BoundaryCurve (or Null if another type)

    DegeneratePcurve (me) returns DegeneratePcurve from StepGeom;
	---Purpose: Returns Value as DegeneratePcurve (or Null if another type)

end SurfaceBoundary;
