-- Created on: 1995-11-03
-- Created by: Laurent BOURESCHE
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SimpleBound from GeomFill inherits Boundary from GeomFill 

	---Purpose: Defines a 3d curve as a boundary for a
    	-- GeomFill_ConstrainedFilling algorithm.
    	-- This curve is unattached to an existing surface.D
      -- Contains fields to allow a reparametrization of curve.

uses
    Pnt            from gp,
    Vec            from gp,
    Function       from Law,
    HCurve         from Adaptor3d

is

    Create(Curve  : HCurve from Adaptor3d;
           Tol3d  : Real from Standard;
    	   Tolang : Real from Standard)
    returns SimpleBound from GeomFill;

    	--- Purpose:
    	-- Constructs the boundary object defined by the 3d curve.
    	-- The surface to be built along this boundary will be in the
    	-- tolerance range defined by Tol3d.
    	-- This object is to be used as a boundary for a
    	-- GeomFill_ConstrainedFilling framework.
    	-- Dummy is initialized but has no function in this class.
    	-- Warning
    	-- Curve is an adapted curve, that is, an object which is an interface between:
    	-- -   the services provided by a 3D curve from the package Geom
    	-- -   and those required of the curve by the computation
    	--   algorithm which uses it.
    	-- The adapted curve is created in one of the following ways:
    	-- -   First sequence:
    	-- Handle(Geom_Curve) myCurve = ... ;
    	-- Handle(GeomAdaptor_HCurve)
    	--     Curve = new
    	-- GeomAdaptor_HCurve(myCurve);
    	-- -   Second sequence:
    	-- // Step 1
    	-- Handle(Geom_Curve) myCurve = ... ;
    	-- GeomAdaptor_Curve Crv (myCurve);
    	-- // Step 2
    	-- Handle(GeomAdaptor_HCurve)
    	--     Curve = new
    	-- GeomAdaptor_HCurve(Crv);
    	-- You use the second part of this sequence if you already
    	-- have the adapted curve Crv.
    	-- The boundary is then constructed with the Curve object:
    	-- Standard_Real Tol = ... ;
    	-- Standard_Real dummy = 0. ;
    	-- myBoundary = GeomFill_SimpleBound
    	-- (Curve,Tol,dummy);
    
    Value(me; 
          U : Real from Standard) 
    returns Pnt from gp;

    D1(me; 
       U : Real from Standard; 
       P : out Pnt from gp; 
       V : out Vec from gp) ;

    Reparametrize(me           : mutable;
    	    	  First, Last  : Real from Standard;
                  HasDF, HasDL : Boolean from Standard;
                  DF, DL       : Real from Standard;
                  Rev          : Boolean from Standard);
		  
    Bounds(me; First, Last : out Real from Standard);

    IsDegenerated(me) returns Boolean from Standard;

fields

    myC3d  : HCurve         from Adaptor3d;
    myPar  : Function       from Law;

end SimpleBound;
