-- Created by: Peter Kurnev
-- Copyright (c) 2010-2012 OPEN CASCADE SAS
-- Copyright (c) 2007-2010 CEA/DEN, EDF R&D, OPEN CASCADE
-- Copyright (c) 2003-2007 OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN, CEDRAT,
--                         EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.
--
class CheckerSI from BOPAlgo 
    inherits PaveFiller from BOPAlgo  
    
    ---Purpose: Checks shape on self-interference.

is
    Create 
    returns CheckerSI from BOPAlgo;  
    ---C++: alias "Standard_EXPORT virtual ~BOPAlgo_CheckerSI();" 
 
    Init  (me:out) 
    is redefined protected;

    SetLevelOfCheck(me:out; 
      theLevel: Integer from Standard); 
    ---Purpose:  Sets the level of checking shape on self-interference.
    --           It defines which interferferences will be checked: 
    --           0 - only V/V; 
    --           1 - V/V and V/E; 
    --           2 - V/V, V/E and E/E; 
    --           3 - V/V, V/E, E/E and V/F;
    --           4 - V/V, V/E, E/E, V/F and E/F; 
    --           5 - all interferences, default value.
 
fields
    myLevelOfCheck: Integer from Standard is protected;
  
end CheckerSI;
