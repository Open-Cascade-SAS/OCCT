-- Created on: 1992-09-28
-- Created by: Ramin BARRETO
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class ErrorHandler from Standard

uses 
    Failure from Standard,
    Boolean from Standard,
    Address from Standard,
    PErrorHandler from Standard,
    Type from Standard
is
    Create returns ErrorHandler;
    	--- Purpose: Create a ErrorHandler (to be used with try{}catch(){}).
    	--           It uses the "setjmp" and "longjmp" routines. 
    	---Level: Advanced
    
    Destroy(me: in out);
    	---Purpose: Unlinks and checks if there is a raised exception.
    	---C++: alias ~
    	---Level: Advanced
        
    Unlink(me: in out);
    	---Purpose: Removes handler from the handlers list
	---Level: Advanced
    
    Catches(me: in out; aType: Type) returns Boolean;
    	---Purpose: Returns "True" if the caught exception has the same type 
    	--          or inherits from "aType"
    	---Level: Advanced
    
    Label(me: in out) returns JmpBuf from Standard;
    	---Purpose: Returns label for jump
    	---C++: inline
    	---C++: return &
    	---Level: Advanced

    Abort(myclass; theError : Failure) is private;
    ---Purpose: A exception is raised but it is not yet caught.
    --          So Abort the current function and transmit the exception
    --          to "calling routines".
    -- Warning: If no catch is prepared for this exception, it displays the
    --          exception name and calls "exit(1)".
    ---Level: Internal

    Error(me) returns Failure;
    	---Purpose: Returns the current Error.

    LastCaughtError(myclass) returns Failure;
    	---Purpose: Returns the caught exception.
    	--    
    	---Level: Advanced
    
    Error(myclass; aError: Failure) is private;
    	---Purpose: Set the Error which will be transmitted to "calling routines".
    	---Level: Advanced
    
    IsInTryBlock(myclass) returns Boolean from  Standard;
    	---Purpose: Test if the code is currently running in a try block
    	---Level: Internal
	
    FindHandler(myclass; theStatus: HandlerStatus from Standard;
    	    	    	 theUnlink: Boolean       from Standard) 
    returns PErrorHandler from Standard is private;
    	---Purpose: Returns the current handler (Top in former implemntations)
    
fields

    myPrevious    : PErrorHandler from Standard;
    myCaughtError : Failure from Standard;
    myLabel       : JmpBuf from Standard;
    myStatus      : HandlerStatus from Standard;
    myThread      : ThreadId from Standard; 
    myCallbackPtr : Address from Standard;

friends
    class Failure,
    class ErrorHandlerCallback
    
end ErrorHandler from Standard;
