-- Created on: 1999-05-06
-- Created by: data exchange team
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SplitSurfaceAngle from ShapeUpgrade inherits SplitSurface from ShapeUpgrade

	---Purpose: Splits a surfaces of revolution, cylindrical, toroidal, 
    	--          conical, spherical so that each resulting segment covers 
	--          not more than defined number of degrees. 

is

    Create (MaxAngle: Real)  returns mutable SplitSurfaceAngle from ShapeUpgrade;
    	---Purpose: Empty constructor.
    
    SetMaxAngle (me: mutable; MaxAngle: Real);
    	---Purpose: Set maximal angle 
    
    MaxAngle (me) returns Real;
    	---Purpose: Returns maximal angle 
    
    Compute(me: mutable; Segment: Boolean) is redefined;
    	---Purpose: Performs splitting of the supporting surface(s).
	---         First defines splitting values, then calls inherited method.

fields

    myMaxAngle: Real;

end SplitSurfaceAngle;
