-- File:        ViewVolume.cdl
-- Created:     Mon Dec  4 12:02:33 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWViewVolume from RWStepVisual

	---Purpose : Read & Write Module for ViewVolume

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     ViewVolume from StepVisual,
     EntityIterator from Interface

is

	Create returns RWViewVolume;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable ViewVolume from StepVisual);

	WriteStep (me; SW : in out StepWriter; ent : ViewVolume from StepVisual);

	Share(me; ent : ViewVolume from StepVisual; iter : in out EntityIterator);

end RWViewVolume;
