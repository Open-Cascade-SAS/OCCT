-- Created on: 1995-03-27
-- Created by: Christophe MARION
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class FaceData from HLRTopoBRep

	---Purpose: Contains the  3 ListOfShape of  a Face  ( Internal
	--          OutLines, OutLines on restriction and IsoLines ).

uses
    Shape       from TopoDS,
    ListOfShape from TopTools

is
    Create returns FaceData from HLRTopoBRep;

    FaceIntL(me) 
    returns ListOfShape from TopTools
	---C++: inline
	---C++: return const &
    is static;

    FaceOutL(me) 
    returns ListOfShape from TopTools
	---C++: inline
	---C++: return const &
    is static;

    FaceIsoL(me) 
    returns ListOfShape from TopTools
	---C++: inline
	---C++: return const &
    is static;

    AddIntL(me : in out) 
    returns ListOfShape from TopTools
	---C++: inline
	---C++: return &
    is static;

    AddOutL(me : in out) 
    returns ListOfShape from TopTools
	---C++: inline
	---C++: return &
    is static;

    AddIsoL(me : in out) 
    returns ListOfShape from TopTools
	---C++: inline
	---C++: return &
    is static;

fields

    myIntL : ListOfShape from TopTools;
    -- For a face the list of internal OutLines.

    myOutL : ListOfShape from TopTools;
    -- For a face the list of not OutLines on restriction.

    myIsoL : ListOfShape from TopTools;
    -- For a face the list of IsoLines.

end FaceData;
