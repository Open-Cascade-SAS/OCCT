-- Created on: 1991-04-15
-- Created by: Philippe DAUTRY
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

generic class QualifiedCurv from GccEnt (TheCurve as any)

	---Purpose: Creates a qualified 2d line.

uses Position from GccEnt

is

Create(Curve     : TheCurve                ;
       Qualifier : Position from GccEnt ) 
returns QualifiedCurv from GccEnt;
-- is private;

Qualified(me) returns TheCurve
is static;

Qualifier(me) returns Position from GccEnt
is static;

IsUnqualified(me) returns Boolean from Standard
is static;
    	---Purpose: Returns true if the solution is unqualified and false in the 
    	--          other cases.

IsEnclosing(me) returns Boolean from Standard
is static;
    	---Purpose: Returns true if the solution is Enclosing the Curv and false in 
    	--          the other cases.

IsEnclosed(me) returns Boolean from Standard
is static;
    	---Purpose: Returns true if the solution is Enclosed in the Curv and false in 
    	--          the other cases.

IsOutside(me) returns Boolean from Standard
is static;
    	---Purpose: Returns true if the solution is Outside the Curv and false in 
    	--          the other cases.

fields

TheQualifier : Position from GccEnt;
TheQualified : TheCurve;

-- friends

-- Unqualified(Obj : Curv2d) from GccEnt,
-- Enclosing  (Obj : Curv2d) from GccEnt,
-- Enclosed   (Obj : Curv2d) from GccEnt,
-- Outside    (Obj : Curv2d) from GccEnt

end QualifiedCurv;


