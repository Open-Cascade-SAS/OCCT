-- File:	GeomAbs.cdl
-- Created:	Mon Feb 22 15:03:40 1993
-- Author:	Modelistation
--		<model@sdsun2>
---Copyright:	 Matra Datavision 1993



package GeomAbs 

	---Purpose: This package gives resources for Geometric applications
	--         
	-- it contains :
	--          CurveType enumeration to describe the different type of 
	--          curves 
	--          
	--          SurfaceType enumeration to describe the different type of
	--          surfaces
	--          
	--          Shape enumeration to  describe the continuity of curve
	--           or surface
	--           
	--          CurveForm enumeration to describe the specific form of
	--          curve 
	--           
	--          SurfaceForm enumeration to describe the specific form of
	--          surface
	--          
	--           BSplKnotDistribution enumeration to describe the 
	--           repartition of set of knots
	--           
	--           UVSense enumeration to describe the orientation of 
	--           the parametric surface 
uses Standard 

is

enumeration CurveType 
       is  Line, Circle, Ellipse, Hyperbola, Parabola,
           BezierCurve, BSplineCurve,OtherCurve end;
    	---Purpose:
    	-- Identifies the type of a curve.
enumeration SurfaceType 
       is  Plane, Cylinder, Cone ,Sphere ,Torus, BezierSurface, 
           BSplineSurface, SurfaceOfRevolution , SurfaceOfExtrusion,
	   OffsetSurface,OtherSurface end;

enumeration Shape is C0, G1, C1, G2, C2, C3, CN;
        --- Purpose :
        -- Provides information about the continuity of a curve:
    	-- -   C0: only geometric continuity.
    	-- -   G1: for each point on the curve, the tangent vectors
    	--   "on the right" and "on the left" are collinear with the same orientation.
    	-- -   C1: continuity of the first derivative. The "C1" curve is
    	--   also "G1" but, in addition, the tangent vectors " on the
    	--   right" and "on the left" are equal.
    	-- -   G2: for each point on the curve, the normalized
    	-- normal vectors "on the right" and "on the left" are equal.
    	-- -   C2: continuity of the second derivative.
    	-- -   C3: continuity of the third derivative.
    	-- -   CN: continuity of the N-th derivative, whatever is the
    	--   value given for N (infinite order of continuity).
    	-- Also provides information about the continuity of a surface:
    	-- -   C0: only geometric continuity.
    	-- -   C1: continuity of the first derivatives; any
    	--   isoparametric (in U or V) of a surface "C1" is also "C1".
    	-- -   G2: for BSpline curves only; "on the right" and "on the
    	--   left" of a knot the computation of the "main curvature
    	-- radii" and the "main directions" (when they exist) gives the same result.
    	-- -   C2: continuity of the second derivative.
    	-- -   C3: continuity of the third derivative.
    	-- -   CN: continuity of any N-th derivative, whatever is the
    	--   value given for N (infinite order of continuity).
    	-- We may also say that a surface is "Ci" in u, and "Cj" in v
    	-- to indicate the continuity of its derivatives up to the order
    	-- i in the u parametric direction, and j in the v parametric direction.


enumeration SurfaceForm is

PlanarForm, ConicalForm, CylindricalForm, ToroidalForm, SphericalForm,
RevolutionForm, RuledForm, QuadricForm, OtherSurfaceForm;
        --- Purpose :
        --  This enumeration is used to note specific surface form.



enumeration CurveForm is

PolylineForm, CircularForm, EllipticForm, HyperbolicForm, ParabolicForm,
OtherCurveForm;
        --- Purpose :
        --  This enumeration is used to note specific curve form.


enumeration BSplKnotDistribution is
NonUniform, Uniform, QuasiUniform, PiecewiseBezier;
        --- Purpose :
        --  This enumeration is used in the classes BSplineCurve and
        --  BSplineSurface to describe the repartition of set of knots.
        --  (comments in classes BSplineCurve and BSplineSurface)


enumeration UVSense is SameUV, SameU, SameV, OppositeUV;
        --- Purpose :
        --  This enumeration is used in the class RectangularTrimmedSurface
        --  to compare the orientation of the basic surface and the orientation
        --  of the trimmed surface and in the class ElementarySurface to know 
        --  the direction of parametrization by comparison with the default
        --  construction mode.

enumeration IsoType is IsoU,IsoV,NoneIso;
	---Purpose: this enumeration describes if a curve is an U isoparaetric
	--          or V isoparametric


enumeration JoinType is Arc, Tangent, Intersection;
	---Purpose: Characterizes the type of a join, built by an algorithm for
    	-- constructing parallel curves, between two consecutive
    	-- arcs of a contour parallel to a given contour.

end GeomAbs;
