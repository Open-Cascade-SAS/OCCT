-- Created on: 2001-06-25
-- Created by: Michael KLOKOV
-- Copyright (c) 2001-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Area3dBuilder from BOP inherits AreaBuilder from BOP

    ---Purpose: 
    	
    -- The algorithm is used to construct Solids from a LoopSet,
    -- where the Loop is the composite topological object of the boundary,
    -- here it is a Shell(s) or block(s) of Faces.
    -- The LoopSet gives an iteration on Loops.
    -- For each Loop  it indicates if it is on the boundary (shell) or if it
    -- results from  an interference (block of faces).
    -- The result of the algorithm is an iteration on areas.
    -- An area is described by a set of Loops. 
    
uses
    LoopSet from BOP,
    LoopClassifier from BOP

is

    Create returns Area3dBuilder from BOP;
    	---Purpose:  
    	--- Empty  Constructor 
    	---
    Create(LS:out LoopSet from BOP;
    	   LC:out LoopClassifier from BOP;
    	   ForceClass: Boolean from Standard = Standard_False)
    	returns Area3dBuilder from BOP;
    	---Purpose:  
    	--- Creates an  object to build solids on
    	--- the (shells,  blocks of faces) of <LS>,  
    	--- using the classifier <LC>. 
	---
    
    InitAreaBuilder(me:                in out;
    	    	    LS:out LoopSet from BOP;
	    	    LC:out LoopClassifier from BOP;
    	    	    ForceClass: Boolean from Standard)
    	is redefined;
    	---Purpose:  
    	--- Initialize the object to find the areas of
    	--- the shapes described by <LS>, 
    	--- using the classifier <LC>. 
	---
    
end Area3dBuilder from BOP;
