-- Created on: 1993-08-10
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class PointsOnSurface from BRep inherits PointRepresentation from BRep

	---Purpose: 

uses

    Surface  from Geom,
    Location from TopLoc

is
    Initialize (P : Real;
    	    	S : Surface  from Geom;
    	        L : Location from TopLoc);
		

    Surface(me) returns any Surface from Geom
	---C++: return const &
    is redefined;
    
    Surface(me : mutable; S : Surface from Geom)
    is redefined;    

fields

    mySurface : Surface from Geom;

end PointsOnSurface;
