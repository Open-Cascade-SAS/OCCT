-- Created on: 1994-12-16
-- Created by: Laurent BUCHARD
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Modified by skv - Fri Jul 14 16:46:18 2006 OCC12627


class Elements from Geom2dHatch


uses 
    Orientation      from TopAbs,
    Lin2d            from gp,
    Pnt2d            from gp,
    Integer          from Standard,
    Element          from Geom2dHatch,
    MapIntegerHasher from TColStd,
    Curve            from Geom2dAdaptor,
    MapOfElements    from Geom2dHatch,
    DataMapIteratorOfMapOfElements from Geom2dHatch

raises         
    DomainError  from Standard,
    NoSuchObject from Standard


is 

    Create
    returns Elements from Geom2dHatch;

    Create(Other : Elements from Geom2dHatch)
    returns Elements from Geom2dHatch;

        

----------------------------------------------------------------------
--               E m u l a t i o n   o f   D a t a M a p  
--               
--                  f r o m  T C o l l e c t  i o n                                                                          
----------------------------------------------------------------------
    Clear(me : in out)
	---C++: alias ~
    is static;

    Bind(me : in out; K : Integer from Standard; I : Element from Geom2dHatch) returns Boolean
    is static;

    IsBound(me; K : Integer from Standard) returns Boolean
    is static;
    
    UnBind(me : in out; K : Integer from Standard) returns Boolean
    is static;
    
    Find(me; K : Integer from Standard) returns any Element from Geom2dHatch
    raises NoSuchObject from Standard  -- when <K> is not in the map.
	---C++: alias operator()
	---C++: return const &
    is static;
    
    ChangeFind(me : in out; K : Integer from Standard) returns any Element from Geom2dHatch
    raises NoSuchObject from Standard  -- when <K> is not in the map.
	---C++: alias operator()
	---C++: return &
    is static;

----------------------------------------------------------------------
--      M e t h o d s   u s e d   b y   t h e   C l a s s i f i e r 
--      
--      see BRepClass_FaceExplorer for the Purposes
----------------------------------------------------------------------

    Reject(me;  P : Pnt2d from gp) 
        returns Boolean from Standard
    is static;
    
-- Modified by skv - Fri Jul 14 16:46:18 2006 OCC12627 Begin
    Segment(me: in out;  P   :     Pnt2d from gp;
    	                 L   : out Lin2d from gp; 
                         Par : out Real)
    returns  Boolean from Standard
    is static;
    
    OtherSegment(me: in out;  P   :     Pnt2d from gp;
    	                      L   : out Lin2d from gp; 
                              Par : out Real)
    returns Boolean from Standard
    is static;
    
-- Modified by skv - Fri Jul 14 16:46:18 2006 OCC12627 End

    InitWires(me : in out)
    is static;
    
    MoreWires(me) returns
       Boolean from Standard
    is static;
    	
    NextWire(me : in out)
    is static;
    
    RejectWire(me; L : Lin2d from gp; 
                 Par : Real  from Standard) 
    	returns Boolean from Standard
    is static;
    
    InitEdges(me : in out)
    is static;
    
    MoreEdges(me) 
       returns Boolean from Standard
    is static;
    
    NextEdge(me  : in out) 
    is static;

    RejectEdge(me; L : Lin2d from gp; 
                 Par : Real  from Standard) 
    	returns Boolean from Standard
    is static;
    
    CurrentEdge(me; E : out Curve  from Geom2dAdaptor;
    	           Or : out Orientation from TopAbs)
    is static;
    

fields 

    myMap    : MapOfElements from Geom2dHatch; 
    Iter     : DataMapIteratorOfMapOfElements;
    NumWire  : Integer from Standard;
    NumEdge  : Integer from Standard;
    myCurEdge: Integer from Standard;
    
end Elements from Geom2dHatch; 
