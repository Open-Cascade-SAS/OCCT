-- Created by: Peter KURNEV
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Set from BOPTools 

	---Purpose: 

uses  
    ShapeEnum from TopAbs,
    Shape from TopoDS,
    ListOfShape from BOPCol,
    BaseAllocator from BOPCol 
    
--raises

is 
    Create 
    	returns Set from BOPTools;  
    ---C++: alias "virtual ~BOPTools_Set();"  
    ---C++: inline 
    
    Create (theAllocator: BaseAllocator from BOPCol)
    	returns Set from BOPTools; 
    ---C++: inline
     
    Assign(me:out;  
    	    Other : Set from BOPTools) 
    	returns Set from BOPTools; 
    ---C++: alias operator =
    ---C++: return &   
    ---C++: inline 
    
    Clear(me:out) 
    	is protected; 
    ---C++: inline
     
    Shape(me) 
    	 returns Shape from TopoDS; 
    ---C++: return const & 
    ---C++: inline 
     
    Add(me:out; 
    	    theS:Shape from TopoDS; 
    	    theType: ShapeEnum from TopAbs);  
    ---C++: inline 
     
    AddEdges(me:out; 
    	    theS:Shape from TopoDS);  
    ---C++: inline 
     
    NbShapes(me) 
    	    returns Integer from Standard; 
    ---C++: inline 
     
    IsEqual(me; 
    	    aOther:Set from BOPTools) 
	returns Boolean from Standard;   
    ---C++: inline 
     
    HashCode(me; 
	    Upper : Integer  from Standard)  
    	returns Integer from Standard;   	 
    ---C++: inline 
    
fields   
    myAllocator : BaseAllocator from BOPCol is protected; 
    myShapes    : ListOfShape from BOPCol is protected;   
    myShape     : Shape from TopoDS is protected; 
    myNbShapes  : Integer from Standard is protected;
    mySum       : Integer from Standard is protected; 
    myUpper     : Integer from Standard is protected; 
    
end Set;
