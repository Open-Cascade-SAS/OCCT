-- Created on: 1991-02-20
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class AnaIntersection from IntAna2d

    ---Purpose: Implementation of the analytical intersection between:
    --          - two Lin2d,
    --          - two Circ2d,
    --          - a Lin2d and a Circ2d,
    --          - an element of gp (Lin2d, Circ2d, Elips2d, Parab2d, Hypr2d)
    --          and another conic.
    --          No tolerance is given for all the intersections: the tolerance
    --          will be the "precision machine".


uses Vec2d            from gp,
     Lin2d            from gp,
     Circ2d           from gp,
     Elips2d          from gp,
     Parab2d          from gp,
     Hypr2d           from gp,
     Conic            from IntAna2d,
     IntPoint         from IntAna2d

raises NotDone    from StdFail,
       OutOfRange from Standard

is

    Create
    
	---Purpose: Empty constructor. IsDone returns False.

    	returns AnaIntersection;


    Create( L1,L2: Lin2d from gp)
    
    	---Purpose: Intersection between two lines.
    
    	returns AnaIntersection
	
	raises NotDone from StdFail;


    Create( C1,C2: Circ2d from gp)
    
    	---Purpose: Intersection between two circles.
    
    	returns AnaIntersection
	
	raises NotDone from StdFail;


    Create( L: Lin2d from gp; C: Circ2d from gp)
    
    	---Purpose: Intersection between a line and a circle.
    
    	returns AnaIntersection
	
	raises NotDone from StdFail;


    Create(L: Lin2d from gp; C: Conic from IntAna2d)
    
    	---Purpose: Intersection between a line and a conic.
    
    	returns AnaIntersection
	
	raises NotDone from StdFail;


    Create(C: Circ2d from gp; Co: Conic from IntAna2d)
    
    	---Purpose: Intersection between a circle and another conic.
    
    	returns AnaIntersection
	
	raises NotDone from StdFail;


    Create(E: Elips2d from gp; C: Conic from IntAna2d)
    
    	---Purpose: Intersection between an ellipse and another conic.
    
    	returns AnaIntersection
	
	raises NotDone from StdFail;


    Create(P: Parab2d from gp; C: Conic from IntAna2d)
    
    	---Purpose: Intersection between a parabola and another conic.
    
    	returns AnaIntersection
	
	raises NotDone from StdFail;


    Create(H: Hypr2d from gp; C: Conic from IntAna2d)
    
    	---Purpose: Intersection between an hyperbola and another conic.
    
    	returns AnaIntersection
	
	raises NotDone from StdFail;


    Perform(me: in out; L1,L2: Lin2d from gp)
    
    	---Purpose: Intersection between two lines.
    
	raises NotDone from StdFail
	
	is static;


    Perform(me: in out; C1,C2: Circ2d from gp)
    
    	---Purpose: Intersection between two circles.
    
	raises NotDone from StdFail
	
	is static;


    Perform(me: in out; L: Lin2d from gp; C: Circ2d from gp)
    
    	---Purpose: Intersection between a line and a circle.
    
	raises NotDone from StdFail
	
	is static;


    Perform(me: in out; L: Lin2d from gp; C: Conic from IntAna2d)
    
    	---Purpose: Intersection between a line and a conic.
    
	raises NotDone from StdFail
	
	is static;


    Perform(me: in out; C: Circ2d from gp; Co: Conic from IntAna2d)
    
    	---Purpose: Intersection between a circle and another conic.
    
	raises NotDone from StdFail
	
	is static;


    Perform(me: in out; E: Elips2d from gp; C: Conic from IntAna2d)
    
    	---Purpose: Intersection between an ellipse and another conic.
    
	raises NotDone from StdFail
	
	is static;


    Perform(me: in out; P: Parab2d from gp; C: Conic from IntAna2d)
    
    	---Purpose: Intersection between a parabola and another conic.
    
	raises NotDone from StdFail
	
	is static;


    Perform(me: in out; H: Hypr2d from gp; C: Conic from IntAna2d)
    
    	---Purpose: Intersection between an hyperbola and another conic.
    
	raises NotDone from StdFail
	
	is static;


    IsDone(me)
    
	---Purpose: Returns TRUE if the computation was succesfull.
    
    	returns Boolean
	---C++: inline
	is static;


    IsEmpty(me)
    
	---Purpose: Returns TRUE when there is no intersection, i-e
	--           - no intersection point
	--           - the elements are not identical.
	--          The element may be parallel in this case.
    
    	returns Boolean
	
	raises NotDone from StdFail
	---C++:inline
	is static;


    IdenticalElements(me)
    
    	---Purpose: For the intersection between an element of gp and a conic
    	--          known by an implicit equation, the result will be TRUE
    	--          if the element of gp verifies the implicit equation.
    	--          For the intersection between two Lin2d or two Circ2d, the
    	--          result will be TRUE if the elements are identical.
    	--          The function returns FALSE in all the other cases.

    	returns Boolean
	
	raises NotDone from StdFail
	---C++:inline
	is static;


    ParallelElements(me)
    
    	---Purpose: For the intersection between two Lin2d or two Circ2d,
    	--          the function returns TRUE if the elements are parallel.
    	--          The function returns FALSE in all the other cases.
    	
	returns Boolean
	
	raises NotDone from StdFail
	---C++:inline
	is static;
    

    NbPoints(me)
    
    	---Purpose: returns the number of IntPoint between the 2 curves.

    	returns Integer
	
	raises NotDone from StdFail
	---C++:inline
	is static;


    Point(me; N: Integer)
    
    	---Purpose: returns the intersection point of range N;
    	--          If (N<=0) or (N>NbPoints), an exception is raised.

    	returns IntPoint from IntAna2d

    	raises NotDone from StdFail,
               OutOfRange from Standard
	---C++:return const &
	---C++:inline
	is static;
	

fields

    done        : Boolean from Standard;
    para        : Boolean from Standard;
    iden        : Boolean from Standard;
    empt        : Boolean from Standard;
    nbp         : Integer from Standard;
    lpnt        : IntPoint from IntAna2d [4];

end AnaIntersection;
