-- Created on: 1990-12-13
-- Created by: Remi Lequette
-- Copyright (c) 1990-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Update:      Frederic Maupas


deferred class TShape from PTopoDS inherits Persistent from Standard

	---Purpose: A TShape  is a topological  structure describing a
	--          set of points in a 2D or 3D space.
	--          

    	--  All the information stored are potentially frozen.  So has
    	--  the "free"  information no  sense in  the D.B. context.  A
    	--  Shape from PTopoDS translated in  a Shape from TopoDS will
    	--  be automatically frozen (not free).

uses
    HArray1OfHShape from PTopoDS,
    HShape          from PTopoDS,
    ShapeEnum       from TopAbs

is
    Initialize;
	---Level: Internal 
	
    ShapeType(me) returns ShapeEnum from TopAbs
	---Purpose: Returns the type as a term of the ShapeEnum enum :
	--          VERTEX, EDGE, WIRE, FACE, ....
    	---Level: Internal 
    is deferred;

    Modified(me) returns Boolean
	---Purpose: Returns the modification flag.
    	---Level: Internal 
    is static;
    
    Modified(me : mutable; M : Boolean)
	---Purpose: Sets the modification flag.
    	---Level: Internal 
    is static;
    
    Checked(me) returns Boolean
       ---Purpose: Returns the checked flag.
    	---Level: Internal 
    is static;
        
    Checked(me : mutable; C : Boolean)
       ---Purpose: Sets the checked flag.
    	---Level: Internal 
    is static;
        
    Orientable(me) returns Boolean
       ---Purpose: Returns the orientability flag.
    	---Level: Internal 
    is static;
    
    Orientable(me : mutable; C : Boolean)
       ---Purpose: Sets the orientability flag.
    	---Level: Internal 
    is static;
    
    Closed(me) returns Boolean
       ---Purpose: Returns the closedness flag.
    	---Level: Internal 
    is static;
    
    Closed(me : mutable; C : Boolean)
       ---Purpose: Sets the closedness flag.
    	---Level: Internal 
    is static;
    
    Infinite(me) returns Boolean
       ---Purpose: Returns the infinity flag.
    	---Level: Internal 
    is static;
    
    Infinite(me : mutable; C : Boolean)
       ---Purpose: Sets the infinity flag.
    	---Level: Internal 
    is static;
    
    Convex(me) returns Boolean
       ---Purpose: Returns the convexness flag.
    	---Level: Internal 
    is static;
    
    Convex(me : mutable; C : Boolean)
       ---Purpose: Sets the convexness flag.
    	---Level: Internal 
    is static;
    
    
    Shapes(me) returns HArray1OfHShape from PTopoDS
       ---Purpose: Sets the hshape list
    	---Level: Internal 
    is static;
    
    Shapes(me; I : Integer from Standard) returns HShape from PTopoDS
       ---Purpose: Sets the i th element of the HShape list
       ---Level: Internal 
    is static;

    Shapes(me: mutable; S : HArray1OfHShape from PTopoDS)
       ---Purpose: Returns the HShape list
        ---Level: Internal 
    is static;
    
    Shapes(me: mutable; I : Integer from Standard; S : HShape from PTopoDS)
       ---Purpose: Returns the i th element of the hshape list
        ---Level: Internal 
    is static;
    
    
fields

    myShapes  : HArray1OfHShape from PTopoDS;
    myFlags   : Integer         from Standard;

end TShape;

