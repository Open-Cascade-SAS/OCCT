-- Created on: 1995-12-04
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package RWStepShape 

uses

	StepData, Interface, TCollection, TColStd, StepShape

is


--class ReadWriteModule;

--class GeneralModule;

class RWAdvancedBrepShapeRepresentation;
class RWAdvancedFace;
class RWBlock;
class RWBooleanResult;
class RWBoxDomain;
class RWBoxedHalfSpace;
class RWBrepWithVoids;
class RWClosedShell;
class RWCompoundShapeRepresentation;
class RWConnectedEdgeSet;
class RWConnectedFaceShapeRepresentation;
class RWConnectedFaceSet;
-- Removed from Rev2 to Rev4 : class RWCsgRepresentation;
class RWCsgShapeRepresentation;
class RWCsgSolid;
class RWDefinitionalRepresentationAndShapeRepresentation; -- abv CAX-IF TRJ4 k1_geo-ac
class RWEdge;
class RWEdgeBasedWireframeModel;
class RWEdgeBasedWireframeShapeRepresentation;
class RWEdgeCurve;
class RWEdgeLoop;
class RWExtrudedAreaSolid;
class RWFace;
class RWFaceBasedSurfaceModel;
class RWFaceBound;
class RWFaceOuterBound;
class RWFaceSurface;
class RWFacetedBrep;
class RWFacetedBrepAndBrepWithVoids; -- Added by FMA
class RWFacetedBrepShapeRepresentation;
class RWGeometricCurveSet;
class RWGeometricSet;
class RWGeometricallyBoundedSurfaceShapeRepresentation;
class RWGeometricallyBoundedWireframeShapeRepresentation;
class RWHalfSpaceSolid;
class RWLoop;
class RWManifoldSolidBrep;
class RWManifoldSurfaceShapeRepresentation;
class RWNonManifoldSurfaceShapeRepresentation;
class RWOpenShell;
class RWOrientedClosedShell;
class RWOrientedEdge;
class RWOrientedFace;
class RWOrientedOpenShell;
class RWOrientedPath;
class RWPath;
class RWPolyLoop;
class RWRevolvedAreaSolid;
class RWRightAngularWedge;
class RWRightCircularCone;
class RWRightCircularCylinder;
class RWShapeRepresentation;
class RWShellBasedSurfaceModel;
class RWSolidModel;
class RWSolidReplica;
class RWSphere;
class RWSweptAreaSolid;
class RWTopologicalRepresentationItem;
class RWTorus;
class RWTransitionalShapeRepresentation;
class RWVertex;
class RWVertexLoop;
class RWVertexPoint;
class RWLoopAndPath;

    --  Added from AP214 CC1 to CC2

class RWContextDependentShapeRepresentation;
class RWShapeDefinitionRepresentation;  -- moved from StepRepr

-- Added from CC2 to DIS
class RWSweptFaceSolid;
class RWExtrudedFaceSolid;
class RWRevolvedFaceSolid;

    -- ABV 18 Apr 00: for dimensions and tolerances (Part 47)
    class RWAngularLocation;
    class RWAngularSize;
    class RWDimensionalCharacteristicRepresentation;
    class RWDimensionalLocation;
    class RWDimensionalLocationWithPath;
    class RWDimensionalSize;
    class RWDimensionalSizeWithPath;
    class RWShapeDimensionRepresentation;

    -- CKY 25 APR 2001 : dim.tol, continued (TR7J)
    class RWLimitsAndFits;
    class RWToleranceValue;
    class RWMeasureQualification;
    class RWPlusMinusTolerance;
    class RWPrecisionQualifier;
    class RWTypeQualifier;

    class RWQualifiedRepresentationItem;
    class RWMeasureRepresentationItemAndQualifiedRepresentationItem;
    
--  Added from AP214 IS to DIS
    
    class RWConnectedFaceSubSet;
    class RWSeamEdge;
    class RWSubedge;
    class RWSubface;
    
--- Added for AP209
    class RWPointRepresentation;

--- added for TR12J (GD&T) 
    class RWShapeRepresentationWithParameters;

	---Package Method ---

--	Init;
	---Purpose: enforced the initialisation of the  libraries

end RWStepShape;
