-- Created on: 1994-02-24
-- Created by: Laurent BOURESCHE
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package BRepLProp

    ---Purpose: These global functions compute the degree of
-- continuity of a curve built by concatenation of two
-- edges at their junction point.

uses Standard, gp, BRepAdaptor, GeomAbs, LProp

is
    
    class CurveTool;
    class SurfaceTool;
    
					    
    class CLProps from BRepLProp 
            instantiates CLProps from LProp(Curve      from BRepAdaptor,
	                                    Vec        from gp,
					    Pnt        from gp,
					    Dir        from gp,
					    CurveTool  from BRepLProp);

    class SLProps from BRepLProp 
            instantiates SLProps from LProp(Surface     from BRepAdaptor,
	                                    SurfaceTool from BRepLProp);

    
    Continuity(C1,C2 : Curve from BRepAdaptor;
    	       u1,u2 : Real from Standard;
               tl,ta : Real from Standard) 
    ---Purpose: Computes the regularity at the junction between C1 and
    --          C2. The point u1 on C1 and the point u2 on  C2 must be
    --          confused.   tl  and ta  are  the  linear  and  angular
    --          tolerance used two compare the derivative.
    returns Shape from GeomAbs;

    
    Continuity(C1,C2 : Curve from BRepAdaptor;
    	       u1,u2 : Real from Standard)
    ---Purpose: The  same  as  preciding   but   using  the   standard
    --          tolerances from package Precision.
    returns Shape from GeomAbs;

end BRepLProp;    
