-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DegenerateToroidalSurface from StepGeom 

inherits ToroidalSurface from StepGeom 

uses

	Boolean from Standard, 
	HAsciiString from TCollection, 
	Axis2Placement3d from StepGeom, 
	Real from Standard
is

	Create returns mutable DegenerateToroidalSurface;
	---Purpose: Returns a DegenerateToroidalSurface


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aPosition : mutable Axis2Placement3d from StepGeom;
	      aMajorRadius : Real from Standard;
	      aMinorRadius : Real from Standard) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aPosition : mutable Axis2Placement3d from StepGeom;
	      aMajorRadius : Real from Standard;
	      aMinorRadius : Real from Standard;
	      aSelectOuter : Boolean from Standard) is virtual;

	-- Specific Methods for Field Data Access --

	SetSelectOuter(me : mutable; aSelectOuter : Boolean);
	SelectOuter (me) returns Boolean;

fields

	selectOuter : Boolean from Standard;

end DegenerateToroidalSurface;
