-- Created on: 1993-11-16
-- Created by: Laurent BOURESCHE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class FaceInterference from ChFiDS 

	---Purpose: interference face/fillet

uses Curve from Geom2d,
     Orientation from TopAbs

is
    Create returns FaceInterference from ChFiDS;
    
    SetInterference(me             : in out; 
    	    	    LineIndex      : Integer from Standard;
		    Trans          : Orientation from TopAbs; 
    	    	    PCurv1 ,PCurv2 : Curve from Geom2d )is static;
    ---C++: inline
    	    	
    SetTransition(me : in out; Trans : Orientation from TopAbs) is static;
    
    SetFirstParameter(me : in out; U1 : Real)    is static;
    ---C++: inline
    	    	
    SetLastParameter(me : in out; U1 : Real)     is static;
    ---C++: inline
    	    	
    SetParameter(me      : in out; 
    	    	 U1      : Real from Standard;
                 IsFirst : Boolean from Standard)
    is static;
  
    LineIndex(me) returns Integer from Standard;
    ---C++: inline
    	    	
    SetLineIndex(me : in out; I : Integer from Standard);
    ---C++: inline
    	    	
    Transition(me) returns Orientation from TopAbs is static;
    ---C++: inline

    PCurveOnFace(me) returns Curve from Geom2d is static;
    ---C++: inline
    ---C++: return const &

    PCurveOnSurf(me) returns Curve from Geom2d is static;
    ---C++: inline
    ---C++: return const &

    ChangePCurveOnFace(me : in out) returns Curve from Geom2d is static;
    ---C++: inline
    ---C++: return &

    ChangePCurveOnSurf(me : in out) returns Curve from Geom2d is static;
    ---C++: inline
    ---C++: return &

    FirstParameter(me) returns Real from Standard is static ;
    ---C++: inline

    LastParameter(me) returns Real from Standard is static;
    ---C++: inline

    Parameter(me; IsFirst : Boolean from Standard) 
    returns Real from Standard is static;

fields

firstParam     : Real        from Standard;
lastParam      : Real        from Standard;
pCurveOnFace   : Curve       from Geom2d;
pCurveOnSurf   : Curve       from Geom2d; 
lineindex      : Integer     from Standard;
LineTransition : Orientation from TopAbs;
end FaceInterference;
