-- Created on: 2004-09-03
-- Created by: Oleg FEDYAEV
-- Copyright (c) 2004-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class CheckResult from BOP
    ---Purpose: contains information about faulty shapes and faulty types
    ---         can't be processed by Boolean Operations

uses

    Shape       from TopoDS,
    ListOfShape from TopTools,
    CheckStatus from BOP

is

    Create
    	returns CheckResult;
    ---Purpose: empty constructor
    
    SetShape1(me: in out; TheShape : Shape from TopoDS);
    ---Purpose: sets ancestor shape (object) for faulty sub-shapes
    
    AddFaultyShape1(me: in out; TheShape: Shape from TopoDS);
    ---Purpose: adds faulty sub-shapes from object to a list
    
    SetShape2(me: in out; TheShape: Shape from TopoDS);
    ---Purpose: sets ancestor shape (tool) for faulty sub-shapes
    
    AddFaultyShape2(me: in out; TheShape: Shape from TopoDS);
    ---Purpose: adds faulty sub-shapes from tool to a list
    
    GetShape1(me)
    	returns Shape from TopoDS;
	---C++: return const &
	---Purpose: returns ancestor shape (object) for faulties

    GetShape2(me)
    	returns Shape from TopoDS;
	---C++: return const &
	---Purpose: returns ancestor shape (tool) for faulties
	
    GetFaultyShapes1(me)
    	returns ListOfShape from TopTools;
	---C++: return const &
	---Purpose: returns list of faulty shapes for object
	
    GetFaultyShapes2(me)
    	returns ListOfShape from TopTools;
	---C++: return const &
	---Purpose: returns list of faulty shapes for tool

    SetCheckStatus(me: in out; TheStatus: CheckStatus from BOP);
    ---Purpose: set status of faulty
    
    GetCheckStatus(me)
    	returns CheckStatus from BOP;
	---Purpose: gets status of faulty
	
fields

    myShape1 : Shape from TopoDS;
    myShape2 : Shape from TopoDS;
    myStatus : CheckStatus from BOP;
    myFaulty1 : ListOfShape from TopTools;
    myFaulty2 : ListOfShape from TopTools;

end CheckResult;
