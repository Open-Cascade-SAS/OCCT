-- Created on: 1995-01-04
-- Created by: Bruno DUMORTIER
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MakeSolid from BRepLib  inherits MakeShape from BRepLib

	---Purpose: Makes a solid from compsolid  or  shells.

uses
    Solid             from TopoDS,
    CompSolid         from TopoDS,
    Shell             from TopoDS, 
    Face              from TopoDS,
    ListOfShape       from TopTools,
    ShapeModification from BRepLib

raises
    NotDone from StdFail
    
is

    Create
	---Level: Public
	---Purpose: Solid covers whole space.
    returns MakeSolid from BRepLib;

    ----------------------------------------------
    -- From CompSolid
    ----------------------------------------------

    Create(S : CompSolid from TopoDS)
	---Purpose: Make a solid from a CompSolid.
	---Level: Public
    returns MakeSolid from BRepLib;

    

    ----------------------------------------------
    -- From shells
    ----------------------------------------------

    Create(S : Shell from TopoDS)
	---Purpose: Make a solid from a shell.
	---Level: Public
    returns MakeSolid from BRepLib;

    
    Create(S1,S2 : Shell from TopoDS)
	---Purpose: Make a solid from two shells.
	---Level: Public
    returns MakeSolid from BRepLib;
    
    Create(S1,S2,S3 : Shell from TopoDS)
	---Purpose: Make a solid from three shells.
	---Level: Public
    returns MakeSolid from BRepLib;
    

    ----------------------------------------------
    -- From solid and shells
    ----------------------------------------------

    Create(So : Solid from TopoDS)
	---Purpose: Make a solid from a solid. Usefull for adding later.
	---Level: Public
    returns MakeSolid from BRepLib;
    
    Create(So : Solid from TopoDS; S : Shell from TopoDS)
	---Purpose: Add a shell to a solid.
	---Level: Public
    returns MakeSolid from BRepLib;
    
	
    ----------------------------------------------
    -- Auxiliary methods
    ----------------------------------------------

    Add(me : in out; S : Shell from TopoDS)
	---Purpose: Add the shell to the current solid.
	---Level: Public
    is static;
    
    ----------------------------------------------
    -- Results
    ----------------------------------------------

    Solid(me) returns Solid from TopoDS
	---Purpose: Returns the new Solid.
	--          
	---C++: return const &
	---C++: alias "Standard_EXPORT operator TopoDS_Solid() const;"
 	---Level: Public
    raises
    	NotDone from StdFail
    is static;

    FaceStatus(me; F: Face from TopoDS) 
    	---Purpose: returns the status of the Face after
    	--          the shape creation. 
	---Level: Public
    returns ShapeModification from BRepLib
    is redefined;
 
fields  

    myDeletedFaces: ListOfShape   from TopTools is protected;

end MakeSolid;
