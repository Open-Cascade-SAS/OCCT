--
-- File:        AlienImage_X11XWDAlienData.cdl
-- Created:     23/03/93
-- Author:      BBL
--
---Copyright:   Matravision 1993
--

class X11XWDAlienData from AlienImage inherits AlienImageData from AlienImage

        ---Version: 0.0

        ---Purpose: This class defines a X11 Alien image.
        ---Keywords:
        ---Warning:
        ---References:

uses
        File                    from OSD,
        AsciiString             from TCollection,
        ColorImage              from Image,
        PseudoColorImage        from Image,
        Image                   from Image,
        X11XColor               from AlienImage,
        X11XWDFileHeader        from AlienImage

raises
        OutOfRange      from Standard,
        TypeMismatch    from Standard

is
        Create returns mutable X11XWDAlienData from AlienImage ;

        Clear( me : in out mutable ) ;
        ---Level: Public
        ---Purpose: Frees memory allocated by X11XWDAlienData
        ---C++: alias ~

        Read ( me : in out mutable ; afile : in out File from OSD )
          returns Boolean from Standard ;
        ---Level: Public
          ---Purpose: Read content of a  X11XWDAlienData object from a file
          --          Returns True if file is a XWD file .

        Write( me : in immutable; afile : in out File from OSD )
          returns Boolean from Standard ;
        ---Level: Public
          ---Purpose: Write content of a  X11XWDAlienData object to a file

        SetName( me : in out mutable ;
                 aName : in AsciiString from TCollection)
        is redefined;
        ---Level: Public
          ---Purpose: Set Image name .

        Name( me : in immutable ) returns AsciiString from TCollection
        is redefined;
          ---C++: return const &
        ---Level: Public
          ---Purpose: Get Image name .

        ToImage( me : in  immutable) 
          returns mutable Image from Image 
          raises TypeMismatch from Standard ;
        ---Level: Public
          ---Purpose : convert a X11XWDAlienData object to a Image object.

        FromImage( me : in out mutable ; anImage : in Image from Image )
          raises TypeMismatch from Standard ;
        ---Level: Public
          ---Purpose : convert a Image object to a X11XWDAlienData object.

        --
        --                      Private Method
        --

        Pixel ( me : in immutable ;     X,Y : in Integer from Standard ) 
                        returns Integer from Standard
                        raises OutOfRange from Standard is private ;
        ---Level: Internal

        SetPixel( me : in out mutable; X,Y   : in Integer from Standard ;
                        Value : in Integer from Standard )
                        raises OutOfRange from Standard is private ;
        ---Level: Internal

        DataSize( me : in immutable)
                returns Integer from Standard is private ;
        ---Level: Internal
           ---Purpose: Compute the imaga data size in byte
           --          from header information

        RedShift( me : in immutable) returns Integer from Standard 
                            raises TypeMismatch from Standard is private ;
           ---Purpose: Compute the red shift for TrueColor X11XWDImage

        GreenShift( me : in immutable) returns Integer from Standard
                            raises TypeMismatch from Standard is private ;
        ---Level: Internal
           ---Purpose: Compute the red shift for TrueColor X11XWDImage

        BlueShift( me : in immutable) returns Integer from Standard
                            raises TypeMismatch from Standard is private ;
        ---Level: Internal
           ---Purpose: Compute the red shift for TrueColor X11XWDImage

        ToPseudoColorImage( me : in immutable) 
          returns PseudoColorImage from Image is private ;
        ---Level: Internal
          ---Purpose : convert a Image object to a AlienImage object.

        ToColorImage( me : in immutable) 
          returns ColorImage from Image is private ;
        ---Level: Internal
          ---Purpose : convert a Image object to a AlienImage object.

        FromPseudoColorImage( me      : in out mutable; 
                              anImage : in PseudoColorImage from Image )
                is private ;
        ---Level: Internal
          ---Purpose : convert a Image object to a X11XWDAlienData object.

        FromColorImage( me : in out mutable;
                        anImage : in ColorImage from Image)
                is private ;
        ---Level: Internal
          ---Purpose : convert a Image object to a X11XWDAlienData object.

fields

        myHeader : X11XWDFileHeader from AlienImage is protected ;

        myColors : Address from Standard  is protected ;
                        -- XColors definition

        myData   : Address from Standard is protected ;
                -- my is a ( unsigned char * ) for 8 bit image , 
                --         ( unsigned int *  ) for 24 bit image .

end ;
 
