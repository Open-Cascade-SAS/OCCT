-- Created on: 1993-07-06
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class CurveOn2Surfaces from PBRep inherits CurveRepresentation from PBRep

	---Purpose: Defines a continuity between two surfaces.

uses
    Surface  from PGeom,
    Location from PTopLoc,
    Shape    from GeomAbs
    
raises
    NullObject from Standard
    
is

    Create(S1 , S2  : Surface  from PGeom;
	   L1 , L2  : Location from PTopLoc;
	   C        : Shape    from GeomAbs)
    returns mutable CurveOn2Surfaces from PBRep;

    Surface(me) returns any Surface from PGeom
    is static;

    Surface2(me) returns any Surface from PGeom
    is static;

    Location2(me) returns Location from PTopLoc
    is static;

    Continuity(me) returns Shape from GeomAbs
    is static;
    
    IsRegularity(me) returns Boolean
	---Purpose: Returns True.
    is redefined;
    
fields
    mySurface    : Surface  from PGeom;
    mySurface2   : Surface  from PGeom;
    myLocation2  : Location from PTopLoc;
    myContinuity : Shape    from GeomAbs;

end CurveOn2Surfaces;
