-- Created on: 1993-02-03
-- Created by: Gilles DEBARBOUILLE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class InstanceParameter from Dynamic

inherits

    Parameter from Dynamic

	---Purpose: This class describes a parameter with a dynamic 
	--          fuzzy instance as value.

uses

    CString from Standard,
    OStream from Standard,
    DynamicInstance from Dynamic


is

    Create(aparameter : CString from Standard)
    
    ---Level: Public 
    
    ---Purpose: Creates an   InstanceParameter  with  <aparameter>  as
    --          identifier.
    
    returns mutable InstanceParameter from Dynamic;
    
    Create(aparameter : CString from Standard; avalue : DynamicInstance from Dynamic) 

    ---Level: Public 
    
    ---Purpose: Creates   an  InstanceParameter  with  <aparameter>  as
    --          identifier and <avalue> as initial value.

    returns mutable InstanceParameter from Dynamic;
    
    Value(me) returns DynamicInstance from Dynamic
    
    ---Level: Public 
    
    ---Purpose: Returns <thevalue>.
    
    is static;
    
    Value(me : mutable ; avalue : DynamicInstance from Dynamic)
    
    ---Level: Public 
    
    ---Purpose: Sets <avalue> to <thevalue>.
    
    is static;

    Dump(me ; astream : in out OStream from Standard)
    
    ---Level: Public 
    
    ---Purpose: Useful for debugging.
    
    is redefined;
    
fields

    thevalue : DynamicInstance from Dynamic;

end InstanceParameter;
