-- Created on: 1993-12-09
-- Created by: Bertand Lesecq
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


private generic class GPixelField from Image (Item as any)

	---Purpose: The class GPixelField represents bi-dimensionnal arrays 
	--          The range of the index start from 0 .

raises
    RangeError from Standard,
    OutOfRange from Standard,
    OutOfMemory from Standard,
    DimensionMismatch from Standard

is
    
    Create (Width, Height:  Integer from Standard) 
    returns  GPixelField from Image
	---Level: Public
    	---Purpose: Creates an array of lower bound <0><0> and upper
    	--          bound <Width-1><Height-1>.   Range from  Standard  error  is
    	--          raised when <Width-1> is less than <0> or <Height-1> is less
    	--          than <0>.
    raises 
    	RangeError  from Standard,
    	OutOfMemory from Standard;


    Create (Width, Height: Integer from Standard; V : Item) 
    returns  GPixelField from Image
	---Level: Public
    	---Purpose: Creates an array of lower bound <0><0> and upper
    	--          bound <Width-1><Height-1>.   Range from  Standard  error  is
    	--          raised when <Width-1> is less than <0> or <Height-1> is less
    	--          than <0>. The array is initialized with <V>.
    raises
    	RangeError  from Standard,
    	OutOfMemory from Standard;

    Destroy (me : in out )
	---Level: Public
    	---Purpose: Frees   the allocated   area corresponding to  the
    	--          array.   If  the array    was  constructed from  a
    	--          DoubleArray the Destroy doesn't delete the area.
        --          
        ---C++: alias ~
    is static;

    Width (me) returns Integer from Standard
	---Level: Public
    	---Purpose: Return the number of columns of <me>.
    	--          
	---C++: inline
    is static ;

    Height (me) returns Integer from Standard
	---Level: Public
    	---Purpose: Returns the number of rows of <me>.
    	--          
        ---C++: inline
    is static;

    UpperX (me) returns Integer from Standard
	---Level: Public
    	---Purpose:  Returns the upper column number of the array.
    	--          
	---C++: inline
    is static ;

    UpperY (me) returns Integer from Standard
	---Level: Public
    	---Purpose:  Returns the upper row number of the array.
    	--          
	---C++: inline
    is static ;

    SetValue (me : in out; X, Y: Integer from Standard; Value: Item) 
	---Level: Public
    	---Purpose: Sets the element of index <X><Y>
    	--          to <Value>.
	---C++: inline
    raises OutOfRange from Standard
    is static ;

    Value (me; X,Y: Integer from Standard) returns any Item
	---Level: Public
    	---Purpose: Returns the value of the element of index 
        --          <X><Y>
    	--
	---C++: inline
    	---C++: alias operator()
    	---C++: return const &
    raises OutOfRange from Standard
    is static;

    ChangeValue (me: in out; X,Y: Integer from Standard) returns any Item
	---Level: Public
    	---Purpose: Returns the value of the element of index 
        --          <X><Y>
    	--
	---C++: inline
    	---C++: alias operator()
    	---C++: return &
    raises OutOfRange from Standard
    is static;

fields

	myWidth       : Integer from Standard ;
        myHeight      : Integer from Standard ;
	myDeletable   : Boolean;
    	myData        : Address;
	
end GPixelField ;
