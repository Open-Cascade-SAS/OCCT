-- Created on: 1993-06-23
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class DSFiller from HLRTopoBRep

	---Purpose: Provides methods  to  fill a HLRTopoBRep_Data.

uses
    Real              from Standard,
    Integer           from Standard,
    Boolean           from Standard,
    Shape             from TopoDS,
    Face              from TopoDS,
    Edge              from TopoDS,
    Vertex            from TopoDS,
    ThePointOfContour from Contap,
    Contour           from Contap,
    Data              from HLRTopoBRep,
    MapOfShapeTool    from BRepTopAdaptor

is
    Insert(myclass;
    	   S     :        Shape          from TopoDS;
	   FO    : in out Contour        from Contap;
    	   DS    : in out Data           from HLRTopoBRep;
	   MST   : in out MapOfShapeTool from BRepTopAdaptor;
           nbIso :        Integer        from Standard);
    ---Purpose: Stores in <DS> the outlines of  <S> using the current
    --          outliner and stores the isolines in <DS> using a Hatcher.
    
    InsertFace(myclass;
               FI         :        Integer      from Standard;
    	       F          :        Face         from TopoDS;
	       FO         : in out Contour      from Contap;
    	       DS         : in out Data         from HLRTopoBRep;
               withPCurve :        Boolean      from Standard)
    ---Purpose: Stores in <DS> the outlines of  <F> using the current
    --          outliner.
    is private;
    
    MakeVertex(myclass;
    	       P   :        ThePointOfContour from Contap;
	       tol :        Real              from Standard;
	       DS  : in out Data              from HLRTopoBRep)
    returns Vertex from TopoDS
	---Purpose: Make a  vertex  from an intersection  point <P>and
	--          store it in the data structure <DS>.
    is private;
    
    InsertVertex(myclass;
    	         P   :        ThePointOfContour from Contap;
                 tol :        Real              from Standard;
		 E   :        Edge              from TopoDS;
	         DS  : in out Data              from HLRTopoBRep)
	---Purpose: Insert a vertex    from an internal   intersection
	--          point <P> on restriction <E>  and store it in  the
	--          data structure <DS>.
    is private;
    
    ProcessEdges(myclass; DS : in out Data from HLRTopoBRep)
	---Purpose: Split all  the edges  with  vertices in   the data
	--          structure.
    is private;
    	
end DSFiller;
