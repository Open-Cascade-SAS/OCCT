-- Created on: 1993-02-03
-- Created by: Christian CAILLET
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Protocol  from StepData  inherits Protocol from Interface

    ---Purpose : Description of Basic Protocol for Step
    --           The class Protocol from StepData itself describes a default
    --           Protocol, which recognizes only UnknownEntities.
    --           Sub-classes will redefine CaseNumber and, if necessary,
    --           NbResources and Resources.

uses CString, Type,
     SequenceOfAsciiString from TColStd, DictionaryOfTransient from Dico,
     DataMapOfTransientInteger from Interface,
     InterfaceModel from Interface,
     EDescr from StepData, ESDescr from StepData, ECDescr from StepData,
     PDescr from StepData

is

    Create returns mutable Protocol from StepData;

    NbResources (me) returns Integer;
    ---Purpose : Gives the count of Protocols used as Resource (can be zero)
    --           Here, No resource

    Resource (me; num : Integer) returns Protocol from Interface;
    ---Purpose : Returns a Resource, given a rank. Here, none

    CaseNumber (me; obj : any Transient) returns Integer  is redefined;
    ---Purpose : Returns a unique positive number for any recognized entity
    --           Redefined to work by calling both TypeNumber and, for a
    --           Described Entity (late binding) DescrNumber

    TypeNumber (me; atype : any Type) returns Integer;
    ---Purpose : Returns a Case Number, specific of each recognized Type
    --           Here, only Unknown Entity is recognized

    	-- --    Specific for StepData    -- --

    SchemaName (me) returns CString  is virtual;
    ---Purpose : Returns the Schema Name attached to each class of Protocol
    --           To be redefined by each sub-class
    --           Here, SchemaName returns "(DEFAULT)"
    -- was C++ : return const

    	-- --    General Services (defined at Norm level)    -- --

    NewModel (me) returns mutable InterfaceModel;
    ---Purpose : Creates an empty Model for Step Norm

    IsSuitableModel (me; model : InterfaceModel)  returns Boolean;
    ---Purpose : Returns True if <model> is a Model of Step Norm

    UnknownEntity (me) returns mutable Transient;
    ---Purpose : Creates a new Unknown Entity for Step (UndefinedEntity)

    IsUnknownEntity (me; ent : Transient) returns Boolean;
    ---Purpose : Returns True if <ent> is an Unknown Entity for the Norm, i.e.
    --           Type UndefinedEntity, status Unknown

    	-- --    About Descriptions (late binding)

    DescrNumber (me; adescr : any EDescr) returns Integer  is virtual;
    ---Purpose : Returns a unique positive CaseNumber for types described by
    --           an EDescr (late binding)
    --  Warning : TypeNumber and DescrNumber must give together a unique
    --           positive case number for each distinct case, type or descr

    AddDescr   (me : mutable; adescr : EDescr; CN : Integer);
    ---Purpose : Records an EDescr with its case number
    --           Also records its name for an ESDescr (simple type): an ESDescr
    --           is then used, for case number, or for type name

    HasDescr   (me) returns Boolean;
    ---Purpose : Tells if a Protocol brings at least one ESDescr, i.e. if it
    --           defines at least one entity description by ESDescr mechanism

    Descr      (me; num : Integer)  returns EDescr;
    ---Purpose : Returns the description attached to a case number, or null

    Descr      (me; name : CString; anylevel : Boolean = Standard_True)
    	returns EDescr;
    ---Purpose : Returns a description according to its name
    --           <anylevel> True (D) : for <me> and its resources
    --           <anylevel> False : for <me> only

    ESDescr    (me; name : CString; anylevel : Boolean = Standard_True)
    	returns ESDescr;
    ---Purpose : Idem as Descr but cast to simple description

    ECDescr    (me; names : SequenceOfAsciiString from TColStd;
    	    	anylevel : Boolean = Standard_True)  returns ECDescr;
    ---Purpose : Returns a complex description according to list of names
    --           <anylevel> True (D) : for <me> and its resources
    --           <anylevel> False : for <me> only


    AddPDescr  (me : mutable; pdescr : PDescr);
    ---Purpose : Records an PDescr

    PDescr     (me; name : CString; anylevel : Boolean = Standard_True)
    	returns PDescr;
    ---Purpose : Returns a parameter description according to its name
    --           <anylevel> True (D) : for <me> and its resources
    --           <anylevel> False : for <me> only

    AddBasicDescr (me : mutable; esdescr : ESDescr);
    ---Purpose : Records an ESDescr, intended to build complex descriptions

    BasicDescr    (me; name : CString; anylevel : Boolean = Standard_True)
    	returns EDescr;
    ---Purpose : Returns a basic description according to its name
    --           <anylevel> True (D) : for <me> and its resources
    --           <anylevel> False : for <me> only

fields

    thedscnum : DataMapOfTransientInteger from Interface;
    thedscnam : DictionaryOfTransient from Dico;
    thepdescr : DictionaryOfTransient from Dico;
    thedscbas : DictionaryOfTransient from Dico;

end Protocol;
