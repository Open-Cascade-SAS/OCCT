-- Created on: 1995-06-12
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class ListOfShapeOn1State from TopOpeBRepDS

---Purpose: represent a list of shape

uses
    
    ListOfShape from TopTools,
    Shape from TopoDS
    
is

    Create returns ListOfShapeOn1State from TopOpeBRepDS;

    ListOnState(me)
    returns ListOfShape from TopTools is static;
    ---C++: return const &

    ChangeListOnState(me : in out)
    returns ListOfShape from TopTools is static;
    ---C++: return &

    IsSplit(me)
    returns Boolean from Standard is static;

    Split(me : in out; B : Boolean = Standard_True) is static;
    Clear(me : in out) is static;	    

fields

    myList : ListOfShape from TopTools;
    mySplits : Integer from Standard;

end ListOfShapeOn1State from TopOpeBRepDS;
