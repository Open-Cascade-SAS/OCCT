-- Created on: 1992-04-30
-- Created by: Remi LEQUETTE
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Circle3D from Draw inherits Drawable3D from Draw

	---Purpose: 

uses
    Circ from gp,
    Color from Draw,
    Display from Draw

is

    Create(C : Circ from gp; A1,A2 : Real; col : Color)
    returns mutable Circle3D;
    
    DrawOn(me; dis : in out Display);

fields

    myCirc  : Circ from gp;
    myA1    : Real;
    myA2    : Real;
    myColor : Color;
    
end Circle3D;

