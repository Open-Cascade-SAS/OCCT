-- Created on: 1998-07-22
-- Created by: data exchange team
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ShapeTolerance from ShapeFix 

	---Purpose: Modifies tolerances of sub-shapes (vertices, edges, faces)

uses

    Shape     from TopoDS,
    ShapeEnum from TopAbs

is
    
    Create returns ShapeTolerance from ShapeFix;

    LimitTolerance (me; shape: Shape from TopoDS;
    	    	        tmin  : Real;
    	    	        tmax  : Real = 0.0;
    	    	        styp : ShapeEnum from TopAbs = TopAbs_SHAPE)
    returns Boolean;
    	---Purpose: Limits tolerances in a shape as follows :
    	--          tmin = tmax -> as SetTolerance (forces)
    	--          tmin = 0   -> maximum tolerance will be <tmax>
    	--          tmax = 0 or not given (more generally, tmax < tmin) ->
    	--             <tmax> ignored, minimum will be <tmin>
    	--          else, maximum will be <max> and minimum will be <min>
    	--          styp = VERTEX : only vertices are set
    	--          styp = EDGE   : only edges are set
    	--          styp = FACE   : only faces are set
    	--          styp = WIRE   : to have edges and their vertices set
    	--          styp = other value : all (vertices,edges,faces) are set
    	--          Returns True if at least one tolerance of the sub-shape has
    	--          been modified

    SetTolerance (me; shape: Shape from TopoDS;
    	    	      preci: Real;
    	    	      styp : ShapeEnum from TopAbs = TopAbs_SHAPE);
    	---Purpose: Sets (enforces) tolerances in a shape to the given value
    	--          styp = VERTEX : only vertices are set
    	--          styp = EDGE   : only edges are set
    	--          styp = FACE   : only faces are set
    	--          styp = WIRE   : to have edges and their vertices set
    	--          styp = other value : all (vertices,edges,faces) are set

end ShapeTolerance;
