-- Created on: 1999-10-14
-- Created by: VKH
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Updated:	GG IMP100701 Add the "depth" field and method
--              to the pixmap object.


deferred class PixMap from Aspect
inherits
    TShared from MMgt
    ---Purpose: This class allows the definition of a pixmap(bitmap)

uses
    Handle                from Aspect,
    Color                 from Quantity

raises
    PixmapDefinitionError	from Aspect,
    PixmapError           from Aspect
is
    Initialize ( aWidth, anHeight : Integer from Standard;
                 aDepth           : Integer from Standard );
    ---Level: Public
    ---Purpose: Initializes the datas of a pixmap with a pixel size
    -- <aWidth>,<anHeight> and depth.

    Destroy ( me : mutable )
    raises PixmapError from Aspect is deferred;
    ---Level: Advanced
    ---Purpose: Destroy the pixmap
    ---Category: Methods to modify the class definition

    Dump ( me ; aFilename : CString from Standard;
           aGammaValue: Real from Standard = 1.0 )
    returns Boolean
    raises PixmapError from Aspect is deferred;
    ---Level: Advanced
    ---Purpose:
    -- Dumps the Bitmap to an image file with
    -- an optional gamma correction value
    -- and returns TRUE if the dump occurs normaly.
    ---Trigger: Raises if pixmap is not defined properly

    PixelColor ( me         : in;
                 theX, theY : in Integer from Standard )
    returns Color from Quantity is deferred;
    ---Purpose:
    -- Returns the pixel color.

	  ----------------------------
    -- Category: Inquire methods
    ----------------------------

    PixmapID ( me ) returns Handle from Aspect
    is deferred;
    ---Level: Advanced
    ---Purpose: Returns the ID of the just created pixmap
    ---Category: Inquire methods

    Size ( me ; aWidth, anHeight : out Integer from Standard )
    is static;
    ---Level: Public
    ---Purpose: Returns the allocated pixmap's size in PIXEL
    ---Category: Inquire methods

    Depth ( me ) returns Integer from Standard
    is static;
    ---Level: Public
    ---Purpose: Returns the allocated pixmap's depth (planes number)
    ---Category: Inquire methods
fields
    myWidth  : Integer from Standard is protected;
    myHeight : Integer from Standard is protected;
    myDepth	 : Integer from Standard is protected;
end PixMap;
