-- File:        VertexPoint.cdl
-- Created:     Mon Dec  4 12:02:33 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWVertexPoint from RWStepShape

	---Purpose : Read & Write Module for VertexPoint

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     VertexPoint from StepShape,
     EntityIterator from Interface

is

	Create returns RWVertexPoint;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable VertexPoint from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : VertexPoint from StepShape);

	Share(me; ent : VertexPoint from StepShape; iter : in out EntityIterator);

end RWVertexPoint;
