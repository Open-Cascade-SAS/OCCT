-- Created on: 1993-04-08
-- Created by: Christian CAILLET
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class CopyControl  from Interface  inherits TShared

    ---Purpose : This deferred class describes the services required by
    --           CopyTool to work. They are very simple and correspond
    --           basically to the management of an indexed map.
    --           But they can be provided by various classes which can
    --           control a Transfer. Each Starting Entity have at most
    --           one Result (Mapping one-one)

uses Transient

raises InterfaceError

is

    Clear  (me : mutable) is deferred;
    ---Purpose : Clears List of Copy Results. Gets Ready to begin another Copy
    --           Process.

    Bind (me : mutable; ent : Transient; res : mutable Transient)
    ---Purpose : Bind a Result to a Starting Entity identified by its Number
    	raises InterfaceError  is deferred;
    --           Error if <num> is already bound or is out of range

    Search (me; ent : Transient; res : out mutable Transient)
    	returns Boolean  is deferred;
    ---Purpose : Searches for the Result bound to a Startingf Entity identified
    --           by its Number.
    --           If Found, returns True and fills <res>
    --           Else, returns False and nullifies <res>

end CopyControl;
