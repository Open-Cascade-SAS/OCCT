-- File:	Geom2d_OffsetCurve.cdl
-- Created:	Wed Mar 24 18:20:16 1993
-- Author:	Philippe DAUTRY
--		<fid@sdsun2>
-- Copyright:	 Matra Datavision 1993

---Copyright:   Matra Datavision 1991


class OffsetCurve from Geom2d inherits Curve from Geom2d

 
        --- Purpose :  
        --  This class implements the basis services for the creation,
        --  edition, modification and evaluation of planar offset curve.
        --  The offset curve is obtained by offsetting by distance along 
        --  the normal to a basis curve defined in 2D space.
        --  The offset curve in this package can be a self intersecting
        --  curve even if the basis curve does not self-intersect.
        --  The self intersecting portions are not deleted at the
        --  construction time.
        --  An offset curve is a curve at constant distance (Offset) from a
        --  basis curve and the offset curve takes its parametrization from
        --  the basis curve. The Offset curve is in the direction of the
        --  normal to the basis curve N.
        --  The distance offset may be positive or negative to indicate the
        --  preferred side of the curve :
        --  . distance offset >0 => the curve is in the direction of N
        --  . distance offset >0 => the curve is in the direction of - N
        --  On the Offset curve :
        --  Value(u) = BasisCurve.Value(U) + (Offset * (T ^ Z)) / ||T ^ Z||
        --  where T is the tangent vector to the basis curve and Z the 
        --  direction of the normal vector to the plane of the curve,
        --  N = T ^ Z defines the offset direction and should not have 
        --  null length. 
        --  
        --  Warnings :
        --  In this package we suppose that the continuity of the offset
        --  curve is one degree less than the continuity of the
        --  basis curve and we don't check that at any point ||T^Z|| != 0.0
        --  
        --  So to evaluate the curve it is better to check that the offset
        --  curve is well defined at any point because an exception could 
        --  be raised. The check is not done in this package at the creation
        --  of the offset curve because the control needs the use of an
        --  algorithm which cannot be implemented in this package.
        --  The OffsetCurve is closed if the first point and the last point
        --  are the same (The distance between these two points is lower or
        --  equal to the Resolution sea package gp) . The OffsetCurve can be
        --  closed even if the basis curve is not closed. 

uses Dir2d    from gp,
     Pnt2d    from gp,
     Trsf2d   from gp,
     Vec2d    from gp,
     Curve    from Geom2d,
     Geometry from Geom2d,
     Shape    from GeomAbs


raises ConstructionError   from Standard,
       RangeError          from Standard,
       NoSuchObject        from Standard,
       UndefinedDerivative from Geom2d,
       UndefinedValue      from Geom2d,
       NotImplemented      from Standard



is


  Create (C : Curve from Geom2d; Offset : Real)   returns mutable OffsetCurve
        --- Purpose : Constructs a curve offset from the basis curve C,
    	-- where Offset is the distance between the offset
    	-- curve and the basis curve at any point.
    	-- A point on the offset curve is built by measuring the
    	-- offset value along a normal vector at a point on C.
    	-- This normal vector is obtained by rotating the
    	-- vector tangential to C at 90 degrees in the
    	-- anti-trigonometric sense. The side of C on which
    	-- the offset value is measured is indicated by this
    	-- normal vector if Offset is positive, or in the inverse
    	-- sense if Offset is negative.
        --   Warnings :
        --  In this package the entities are not shared. The OffsetCurve is
        --  built with a copy of the curve C. So when C is modified the
        --  OffsetCurve is not modified 
	--  Warning!  ConstructionError  raised if the basis curve C is not at least C1.
        --  No check is done to know if ||V^Z|| != 0.0 at any point.
     raises ConstructionError;

        

  Reverse (me : mutable);
        --- Purpose : Changes the direction of parametrization of <me>.
    	--     As a result:
    	-- - the basis curve is reversed,
    	-- - the start point of the initial curve becomes the end
    	--   point of the reversed curve,
    	-- - the end point of the initial curve becomes the start
    	--   point of the reversed curve, and
    	-- - the first and last parameters are recomputed.


  ReversedParameter(me; U : Real) returns Real;
    	---Purpose: Computes the parameter on the reversed curve for
    	-- the point of parameter U on this offset curve.


  SetBasisCurve (me : mutable; C : Curve from Geom2d)
     raises ConstructionError;
        --- Purpose : Changes this offset curve by assigning C as the
    	-- basis curve from which it is built.
    	-- Exceptions
    	-- Standard_ConstructionError if the curve C is not at least "C1" continuous.

  SetOffsetValue (me : mutable; D : Real);
        --- Purpose :  Changes this offset curve by assigning D as the offset value.
        
  BasisCurve (me) returns Curve from Geom2d;
        --- Purpose : Returns the basis curve of this offset curve. The basis curve can be an offset curve.
    	


  Continuity (me)  returns Shape from GeomAbs;
        --- Purpose :
        --  Continuity of the Offset curve :
        --  C0 : only geometric continuity,
        --  C1 : continuity of the first derivative all along the Curve,
        --  C2 : continuity of the second derivative all along the Curve,
        --  C3 : continuity of the third derivative all along the Curve,
        --  G1 : tangency continuity all along the Curve,
        --  G2 : curvature continuity all along the Curve,
        --  CN : the order of continuity is infinite.
        --   Warnings :
        --  Returns the continuity of the basis curve - 1. 
        --  The offset curve must have a unique normal direction defined
        --  at any point.





        --- Purpose  : Value and derivatives
        --  
        --  Warnings :
        --  The exception UndefinedValue or UndefinedDerivative is 
        --  raised if it is not possible to compute a unique offset
        --  direction.
        --  If T is the first derivative with not null length and
        --  Z the direction normal to the plane of the curve, the
        --  relation ||T(U) ^ Z|| != 0  must be satisfied to evaluate
        --  the offset curve.
        --  No check is done at the creation time and we suppose
        --  in this package that the offset curve is well defined.


  D0 (me; U : Real; P : out Pnt2d)
     raises UndefinedValue;
 	---Purpose:  Warning! this should not be called 
        --          if the basis curve is not at least C1. Nevertheless
        --          if used on portion where the curve is C1, it is OK
 


  D1 (me; U : Real; P : out Pnt2d; V1 : out Vec2d)
     raises UndefinedDerivative;
        ---Purpose:  Warning! this should not be called 
        --           if the continuity of the basis curve is not C2.
        --           Nevertheless, it's OK to use it  on portion 
        --           where the curve is C2



  D2 (me; U : Real; P : out Pnt2d; V1, V2 : out Vec2d)
     raises UndefinedDerivative;
        ---Purpose:  Warning!  This  should  not  be called 
        --           if the continuity of the basis curve is not C3.
        --           Nevertheless, it's OK to use it  on portion 
        --           where the curve is C3  

  D3 (me; U : Real; P : out Pnt2d; V1, V2, V3 : out Vec2d)
     raises UndefinedDerivative;

     	---Purpose:  Warning! This should not be called 
        --           if the continuity of the basis curve is not C4.
        --           Nevertheless, it's OK to use it  on portion 
        --           where the curve is C4          

  DN (me; U : Real; N : Integer)   returns Vec2d
        --- Purpose : The returned vector gives the value of the derivative
        --  for the order of derivation N.      
    	--  Warning! this should not be called 
    	--        raises  UndefunedDerivative   if the continuity of the basis curve is not CN+1.
        --           Nevertheless, it's OK to use it  on portion 
        --           where the curve is CN+1  
    	-- raises  RangeError if N < 1. 
   	-- raises  NotImplemented if N > 3. 
    
     raises UndefinedDerivative,

            RangeError,
            NotImplemented; 



        --- Purpose : The following functions compute the value and derivatives
        --  on the offset curve and returns the derivatives on the
        --  basis curve too.  
        --  The computation of the value and derivatives on the basis
        --  curve are used to evaluate the offset curve
        --  Warnings :
        --  The exception UndefinedValue or UndefinedDerivative is 
        --  raised if it is not possible to compute a unique offset direction.


  Value (me; U : Real; P, Pbasis : out Pnt2d; V1basis : out Vec2d)
     raises UndefinedValue;

    	---Purpose:  Warning! this should not be called 
        --          if the basis curve is not at least C1. Nevertheless
        --          if used on portion where the curve is C1, it is OK 
  

  D1 (me; U : Real; P, Pbasis : out Pnt2d;
      V1, V1basis, V2basis : out Vec2d)
     raises UndefinedDerivative;

        ---Purpose:  Warning! this should not be called 
        --           if the continuity of the basis curve is not C1.
        --           Nevertheless, it's OK to use it  on portion 
        --           where the curve is C1

  D2 (me; U : Real; P, Pbasis : out Pnt2d;  V1, V2, V1basis, V2basis, 
      V3basis : out Vec2d)
     raises UndefinedDerivative;

    	---Purpose:  Warning! this should not be called 
        --           if the continuity of the basis curve is not C3.
        --           Nevertheless, it's OK to use it  on portion 
        --           where the curve is C3 

  FirstParameter (me)  returns Real;

  LastParameter (me)   returns Real;
    	---Purpose: Returns the value of the first or last parameter of this
    	-- offset curve. The first parameter corresponds to the
    	-- start point of the curve. The last parameter
    	-- corresponds to the end point.
    	-- Note: the first and last parameters of this offset curve
    	-- are also the ones of its basis curve.
        
  Offset (me)          returns Real;
    	---Purpose: Returns the offset value of this offset curve.

  IsClosed (me)   returns Boolean;
        --- Purpose :
        --  Returns True if the distance between the start point 
        --  and the end point of the curve is lower or equal to 
        --  Resolution from package gp.


  IsCN (me; N : Integer)  returns Boolean
        --- Purpose : Is the order of continuity of the curve N ?
        --   Warnings :
        --  This method answer True if the continuity of the basis curve 
        --  is N + 1.  We suppose in this class that a normal direction
        --  to the basis curve (used to compute the offset curve) is 
        --  defined at any point on the basis curve.
     raises RangeError;
        --- Purpose : Raised if N < 0.


  IsPeriodic (me)  returns Boolean;
        --- Purpose : Is the parametrization of a curve is periodic ?
        --  If the basis curve is a circle or an ellipse the corresponding
        --  OffsetCurve is periodic. If the basis curve can't be periodic 
        --  (for example BezierCurve) the OffsetCurve can't be periodic.


  Period (me) returns Real from Standard
    	---Purpose: Returns the period of this offset curve, i.e. the period
    	-- of the basis curve of this offset curve.
    	-- Exceptions
    	-- Standard_NoSuchObject if the basis curve is not periodic.
  raises  NoSuchObject from Standard
  is redefined;


  Transform (me : mutable; T : Trsf2d);
        ---Purpose : Applies the transformation T to this offset curve.
    	-- Note: the basis curve is also modified.

  TransformedParameter(me; U : Real; T : Trsf2d from gp) returns Real
	---Purpose: Returns the  parameter on the  transformed  curve for
	--          the transform of the point of parameter U on <me>.
	--          
	--          me->Transformed(T)->Value(me->TransformedParameter(U,T))
	--          
	--          is the same point as
	--          
	--          me->Value(U).Transformed(T)
	--          
	--          This methods calls the basis curve method.
     is redefined;  

  ParametricTransformation(me; T : Trsf2d from gp) returns Real
	---Purpose: Returns a  coefficient to compute the parameter on
	--          the transformed  curve  for  the transform  of the
	--          point on <me>.
	--          
	--          Transformed(T)->Value(U * ParametricTransformation(T))
	--          
	--          is the same point as
	--          
	--          Value(U).Transformed(T)
	--          
	--          This methods calls the basis curve method.
     is redefined;  



  Copy (me)  returns mutable like me;
    	---Purpose: Creates a new object, which is a copy of this offset curve.     
fields

  basisCurve  : Curve from Geom2d;
  offsetValue : Real;

end;
