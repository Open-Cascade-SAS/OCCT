-- Created on: 1993-02-22
-- Created by: Philippe DAUTRY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class CartesianPoint from PGeom inherits Point from PGeom

        ---Purpose : Point defined  in  3D space with its 3  cartesian
        --         coordinates X, Y, Z.
        --         
    	---See Also : CartesianPoint from Geom.

uses Pnt from gp

is


  Create returns mutable CartesianPoint from PGeom;
        ---Purpose : Returns a CartesianPoint with default values..
    	---Level: Internal 


  Create (aPnt : Pnt from gp) returns mutable CartesianPoint from PGeom;
        ---Purpose : Returns a CartesianPoint built with <aPnt>.
    	---Level: Internal 


  Pnt (me : mutable; aPnt : Pnt from gp);
        ---Purpose : Set the field pnt.
    	---Level: Internal 


  Pnt (me)  returns Pnt;
        ---Purpose : Returns the value of the field pnt.
    	---Level: Internal 


fields

    pnt : Pnt from gp;

end;
