-- Created on: 2000-09-29
-- Created by: Andrey BETENEV
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Tool from STEPConstruct 

    ---Purpose: Provides basic functionalities for tools which are intended
    --          for encoding/decoding specific STEP constructs
    --
    --          It is initialized by WorkSession and allows easy access to 
    --          its fields and internal data such as Model, TP and FP
    --
    --          NOTE: Call to method Graph() with True (or for a first time,
    --          if you have updated the model since last computation of model) 
    --          can take a time, so it is recommended to avoid creation of 
    --          this (and derived) tool multiple times

uses
    WorkSession      from XSControl,
    InterfaceModel   from Interface,
    Graph            from Interface,
    HGraph           from Interface,
    FinderProcess    from Transfer,
    TransientProcess from Transfer

is

    Create returns Tool;
    	---Purpose: Creates an empty tool

    Create (WS: WorkSession from XSControl) returns Tool;
    	---Purpose: Creates a tool and loads it with worksession
	
    SetWS (me: in out; WS: WorkSession from XSControl) 
    returns Boolean is protected;
    	---Purpose: Load worksession; returns True if succeeded
	--          Returns False if either FinderProcess of TransientProcess
	--          cannot be obtained or are Null
	
    WS (me) returns WorkSession from XSControl;
    	---Purpose: Returns currently loaded WorkSession
	---C++: return const &
	---C++: inline
    
    Model (me) returns InterfaceModel from Interface;
    	---Purpose: Returns current model (Null if not loaded)
	---C++: inline
    
    Graph (me; recompute: Boolean = Standard_False) returns Graph from Interface;
    	---Purpose: Returns current graph (recomputing if necessary)
	---C++: return const &
	---C++: inline
    
    TransientProcess (me) returns TransientProcess from Transfer;
    	---Purpose: Returns TransientProcess (reading; Null if not loaded)
	---C++: return const &
	---C++: inline
 
    FinderProcess (me) returns FinderProcess from Transfer;
    	---Purpose: Returns FinderProcess (writing; Null if not loaded)
	---C++: return const &
	---C++: inline
 	
fields

    myWS           : WorkSession from XSControl;
    myFinderProcess: FinderProcess from Transfer;
    myTransientProcess: TransientProcess from Transfer;
    myHGraph       : HGraph from Interface; -- for optimization (no recomutings)

end Tool;
