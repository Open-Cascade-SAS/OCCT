-- Created on: 2000-05-11
-- Created by: data exchange team
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1

class DocumentFile from StepBasic
inherits Document from StepBasic

    ---Purpose: Representation of STEP entity DocumentFile

uses
    HAsciiString from TCollection,
    DocumentType from StepBasic,
    CharacterizedObject from StepBasic

is
    Create returns DocumentFile from StepBasic;
	---Purpose: Empty constructor

    Init (me: mutable; aDocument_Id: HAsciiString from TCollection;
                       aDocument_Name: HAsciiString from TCollection;
                       hasDocument_Description: Boolean;
                       aDocument_Description: HAsciiString from TCollection;
                       aDocument_Kind: DocumentType from StepBasic;
                       aCharacterizedObject_Name: HAsciiString from TCollection;
                       hasCharacterizedObject_Description: Boolean;
                       aCharacterizedObject_Description: HAsciiString from TCollection);
	---Purpose: Initialize all fields (own and inherited)

    CharacterizedObject (me) returns CharacterizedObject from StepBasic;
	---Purpose: Returns data for supertype CharacterizedObject
    SetCharacterizedObject (me: mutable; CharacterizedObject: CharacterizedObject from StepBasic);
	---Purpose: Set data for supertype CharacterizedObject

fields
    theCharacterizedObject: CharacterizedObject from StepBasic; -- supertype

end DocumentFile;
