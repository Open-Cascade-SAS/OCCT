-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ApplicationProtocolDefinition from StepBasic 

inherits TShared from MMgt

uses

	HAsciiString from TCollection, 
	Integer from Standard, 
	ApplicationContext from StepBasic
is

	Create returns mutable ApplicationProtocolDefinition;
	---Purpose: Returns a ApplicationProtocolDefinition

	Init (me : mutable;
	      aStatus : mutable HAsciiString from TCollection;
	      aApplicationInterpretedModelSchemaName : mutable HAsciiString from TCollection;
	      aApplicationProtocolYear : Integer from Standard;
	      aApplication : mutable ApplicationContext from StepBasic) is virtual;

	-- Specific Methods for Field Data Access --

	SetStatus(me : mutable; aStatus : mutable HAsciiString);
	Status (me) returns mutable HAsciiString;
	SetApplicationInterpretedModelSchemaName(me : mutable; aApplicationInterpretedModelSchemaName : mutable HAsciiString);
	ApplicationInterpretedModelSchemaName (me) returns mutable HAsciiString;
	SetApplicationProtocolYear(me : mutable; aApplicationProtocolYear : Integer);
	ApplicationProtocolYear (me) returns Integer;
	SetApplication(me : mutable; aApplication : mutable ApplicationContext);
	Application (me) returns mutable ApplicationContext;

fields

	status : HAsciiString from TCollection;
	applicationInterpretedModelSchemaName : HAsciiString from TCollection;
	applicationProtocolYear : Integer from Standard;
	application : ApplicationContext from StepBasic;

end ApplicationProtocolDefinition;
