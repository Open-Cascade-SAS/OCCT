-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class SurfaceCurve from StepGeom 

inherits Curve from StepGeom 

uses

	HArray1OfPcurveOrSurface from StepGeom, 
	PreferredSurfaceCurveRepresentation from StepGeom, 
	PcurveOrSurface from StepGeom, 
	HAsciiString from TCollection
is

	Create returns mutable SurfaceCurve;
	---Purpose: Returns a SurfaceCurve


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aCurve3d : mutable Curve from StepGeom;
	      aAssociatedGeometry : mutable HArray1OfPcurveOrSurface from StepGeom;
	      aMasterRepresentation : PreferredSurfaceCurveRepresentation from StepGeom) is virtual;

	-- Specific Methods for Field Data Access --

	SetCurve3d(me : mutable; aCurve3d : mutable Curve);
	Curve3d (me) returns mutable Curve;
	SetAssociatedGeometry(me : mutable; aAssociatedGeometry : mutable HArray1OfPcurveOrSurface);
	AssociatedGeometry (me) returns mutable HArray1OfPcurveOrSurface;
	AssociatedGeometryValue (me; num : Integer) returns PcurveOrSurface;
	NbAssociatedGeometry (me) returns Integer;
	SetMasterRepresentation(me : mutable; aMasterRepresentation : PreferredSurfaceCurveRepresentation);
	MasterRepresentation (me) returns PreferredSurfaceCurveRepresentation;

fields

	curve3d : Curve from StepGeom;
	associatedGeometry : HArray1OfPcurveOrSurface from StepGeom; -- a SelectType
	masterRepresentation : PreferredSurfaceCurveRepresentation from StepGeom; -- an Enumeration

end SurfaceCurve;
