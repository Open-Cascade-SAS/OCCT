-- Created on: 1991-07-17
-- Created by: Isabelle GRIGNON
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class FunctionAllRoots from math 

	---Purpose: This algorithm uses a sample of the function to find
	--          all intervals on which the function is null, and afterwards
	--          uses the FunctionRoots algorithm to find the points
	--          where the function is null outside the "null intervals".
    	-- Knowledge of the derivative is required.


uses FunctionSample         from math,
     FunctionRoots          from math,
     FunctionWithDerivative from math,
     SequenceOfReal         from TColStd,
     SequenceOfInteger      from TColStd,
     OStream                from Standard

raises OutOfRange   from Standard,
       NotDone      from StdFail,
       NumericError from Standard

is

    Create(F: in out FunctionWithDerivative from math; 
           S: FunctionSample from math;
           EpsX, EpsF, EpsNul: Real)

	---Purpose: The algorithm uses the sample to find intervals on which
	--          the function is null. An interval is found if, for at least
	--          two consecutive points of the sample, Ui and Ui+1, we get
	--          |F(Ui)|<=EpsNul and |F(Ui+1)|<=EpsNul. The real bounds of
	--          an interval are computed with the FunctionRoots.
	--          algorithm.
	--          Between two intervals, the roots of the function F are
	--          calculated using the FunctionRoots algorithm.
	
	returns FunctionAllRoots
	    
	raises NumericError from Standard;


    IsDone(me)
    
	---Purpose: Returns True if the computation has been done successfully.
    	---C++: inline

    returns Boolean
    is static;


    NbIntervals(me)
	---Purpose: Returns the number of intervals on which the function
	--          is Null.
	--          An exception is raised if IsDone returns False.
        ---C++: inline

   returns Integer
   raises NotDone from StdFail
   is static;


    GetInterval(me; Index: Integer; A,B: out Real)
	---Purpose: Returns the interval of parameter of range Index.
	--          An exception is raised if IsDone returns False;
	--          An exception is raised if Index<=0 or Index >Nbintervals.
    	---C++: inline
    
    raises NotDone from StdFail, OutOfRange from Standard
    is static;


    GetIntervalState(me; Index: Integer; IFirst, ILast: out Integer)
    	---Purpose: returns the State Number associated to the interval Index.
	--          An exception is raised if IsDone returns False;
	--          An exception is raised if Index<=0 or Index >Nbintervals.
    	---C++: inline

    raises NotDone from StdFail, OutOfRange from Standard
    is static;


    NbPoints(me)
	---Purpose: returns the number of points where the function is Null.
	--          An exception is raised if IsDone returns False.
    	---C++: inline
    
    returns Integer
    raises NotDone from StdFail
    is static;


    GetPoint(me; Index: Integer)
	---Purpose: Returns the parameter of the point of range Index.
	--          An exception is raised if IsDone returns False;
	--          An exception is raised if Index<=0 or Index >NbPoints.
    	---C++: inline
    
    returns Real
    raises NotDone from StdFail, OutOfRange from Standard
    is static;


    GetPointState(me; Index: Integer)
    	---Purpose: returns the State Number associated to the point Index.
	--          An exception is raised if IsDone returns False;
	--          An exception is raised if Index<=0 or Index >Nbintervals.
    	---C++: inline

    returns Integer
    raises NotDone from StdFail, OutOfRange from Standard
    is static;


    Dump(me; o: in out OStream)
	---Purpose: Prints on the stream o information on the current state 
    	--          of the object.

    is static;

fields

    done: Boolean;
    pdeb: SequenceOfReal    from TColStd;
    pfin: SequenceOfReal    from TColStd;
    piso: SequenceOfReal    from TColStd;
    ideb: SequenceOfInteger from TColStd;
    ifin: SequenceOfInteger from TColStd;
    iiso: SequenceOfInteger from TColStd;

end FunctionAllRoots;
