-- File:        OverRidingStyledItem.cdl
-- Created:     Fri Dec  1 11:11:23 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class OverRidingStyledItem from StepVisual 

inherits StyledItem from StepVisual 

uses

	HAsciiString from TCollection, 
	HArray1OfPresentationStyleAssignment from StepVisual, 
	RepresentationItem from StepRepr
is

	Create returns mutable OverRidingStyledItem;
	---Purpose: Returns a OverRidingStyledItem


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aStyles : mutable HArray1OfPresentationStyleAssignment from StepVisual;
	      aItem : mutable RepresentationItem from StepRepr) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aStyles : mutable HArray1OfPresentationStyleAssignment from StepVisual;
	      aItem : mutable RepresentationItem from StepRepr;
	      aOverRiddenStyle : mutable StyledItem from StepVisual) is virtual;

	-- Specific Methods for Field Data Access --

	SetOverRiddenStyle(me : mutable; aOverRiddenStyle : mutable StyledItem);
	OverRiddenStyle (me) returns mutable StyledItem;

fields

	overRiddenStyle : StyledItem from StepVisual;

end OverRidingStyledItem;
