-- Created on: 1995-01-23
-- Created by: Mister rmi
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



package SelectBasics 

	---Purpose:  kernel of dynamic selection:
	--           - contains the algorithm to sort the sensitive areas
	--           before the selection action;->quick selection of
	--           an item in a set of items...
	--           - contains the entities able to give the algorithm
	--             sensitive areas .

uses
    Bnd,
    TCollection,
    TColStd,
    Standard,
    MMgt,
    gp,
    TColgp,
    TopLoc
    

is


    deferred class EntityOwner;
    ---Purpose: entity able to set multiple owners for a SensitiveEntity;

    class SortAlgo; 
    ---Purpose: sort algorithm for 2D rectangles.

    class BasicTool;
    ---Purpose: give Tools for sorting Selection results
    --          (example : sensitive entities matching)

    class ListOfBox2d instantiates List from TCollection 
    (Box2d from Bnd);
    

    class SequenceOfOwner instantiates Sequence from TCollection 
    (EntityOwner);
    


    deferred class SensitiveEntity;
    ---Purpose: general entity able to give sensitive areas 


    class ListOfSensitive instantiates List from TCollection 
    (SensitiveEntity);

    imported PickArgs;
    ---Purpose: Structure to provide all-in-one information on picking arguments
    -- for "Matches" method of SelectBasics_SensitiveEntity.

    MaxOwnerPriority returns Integer;
    
    MinOwnerPriority returns Integer;


end SelectBasics;
