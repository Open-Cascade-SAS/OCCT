-- Created on: 1995-12-06
-- Created by: Frederic MAUPAS
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class DirectionCountSelect from StepVisual

    -- a Select Type (hand generated)

uses

    Integer from Standard
    
is

    Create returns DirectionCountSelect;
    
    SetTypeOfContent(me : in out; aTypeOfContent : Integer);

    TypeOfContent(me) returns Integer;
	--        1 -> UDirectionCount
	--        2 -> VDirectionCount

    UDirectionCount(me) returns Integer from Standard;
    
    SetUDirectionCount(me : in out; aUDirectionCount : Integer from Standard);
    
    VDirectionCount(me) returns Integer from Standard;
    
    SetVDirectionCount(me : in out; aUDirectionCount : Integer from Standard);


fields

    theUDirectionCount : Integer from Standard;
    theVDirectionCount : Integer from Standard;
    theTypeOfContent   : Integer from Standard;

end DirectionCountSelect;
