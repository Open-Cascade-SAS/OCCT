-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Ellipse from StepGeom 

inherits Conic from StepGeom 

uses

	Real from Standard, 
	HAsciiString from TCollection, 
	Axis2Placement from StepGeom
is

	Create returns Ellipse;
	---Purpose: Returns a Ellipse


	Init (me : mutable;
	      aName : HAsciiString from TCollection;
	      aPosition : Axis2Placement from StepGeom) is redefined;

	Init (me : mutable;
	      aName : HAsciiString from TCollection;
	      aPosition : Axis2Placement from StepGeom;
	      aSemiAxis1 : Real from Standard;
	      aSemiAxis2 : Real from Standard) is virtual;

	-- Specific Methods for Field Data Access --

	SetSemiAxis1(me : mutable; aSemiAxis1 : Real);
	SemiAxis1 (me) returns Real;
	SetSemiAxis2(me : mutable; aSemiAxis2 : Real);
	SemiAxis2 (me) returns Real;

fields

	semiAxis1 : Real from Standard;
	semiAxis2 : Real from Standard;

end Ellipse;
