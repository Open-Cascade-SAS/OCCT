-- Created on: 1999-11-26
-- Created by: Andrey BETENEV
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0

class ClassifiedItem from StepAP203
inherits SelectType from StepData

    ---Purpose: Representation of STEP SELECT type ClassifiedItem

uses
    ProductDefinitionFormation from StepBasic,
    AssemblyComponentUsage from StepRepr

is
    Create returns ClassifiedItem from StepAP203;
	---Purpose: Empty constructor

    CaseNum (me; ent: Transient) returns Integer;
	---Purpose: Recognizes a kind of ClassifiedItem select type
	--          1 -> ProductDefinitionFormation from StepBasic
	--          2 -> AssemblyComponentUsage from StepRepr
	--          0 else

    ProductDefinitionFormation (me) returns ProductDefinitionFormation from StepBasic;
	---Purpose: Returns Value as ProductDefinitionFormation (or Null if another type)

    AssemblyComponentUsage (me) returns AssemblyComponentUsage from StepRepr;
	---Purpose: Returns Value as AssemblyComponentUsage (or Null if another type)

end ClassifiedItem;
