-- Created on: 1992-05-18
-- Created by: Stephan GARNAUD (ARM)
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Updated:       J.P. TIRAULT August 1993
--                All classes are static class.


class Directory from OSD 

 ---Purpose: Management of directories 
 
inherits FileNode 

uses Protection, Path 

is
 Create returns Directory;
    ---Purpose: Creates Directory object.
    --          It is initiliazed to an empty name.
    ---Level: Public

 Create (Name : Path) returns Directory;
    ---Purpose: Creates Directory object initialized with Name.
    ---Level: Public

 Build (me : in out ; Protect : Protection) is static;
    ---Purpose: Creates (physically) a directory.
    --          When a directory of the same name already exists, no error is
    --          returned, and only <Protect> is applied to the existing directory.
    --
    --          If Build is used and <me> is instantiated without a name,
    --          OSDError is raised.
    ---Level: Public

 BuildTemporary (myclass ) returns Directory;
    ---Purpose: Creates a temporary Directory in current directory.
    --          This directory is automatically removed when object dies.
    ---Level: Public
                                                    
end Directory from OSD;


