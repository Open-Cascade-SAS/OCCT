-- Created by: Peter KURNEV
-- Copyright (c) 2010-2012 OPEN CASCADE SAS
-- Copyright (c) 2007-2010 CEA/DEN, EDF R&D, OPEN CASCADE
-- Copyright (c) 2003-2007 OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN, CEDRAT,
--                         EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class PassKeyBoolean from BOPDS 
    inherits  PassKey from BOPDS 
	---Purpose: 

uses 
    BaseAllocator from BOPCol 
     
--raises

is 
    Create  
    	returns PassKeyBoolean from BOPDS;  
    ---C++: inline 
    ---C++: alias "virtual ~BOPDS_PassKeyBoolean();"  
      
    Create  (theAllocator: BaseAllocator from BOPCol) 
    	returns PassKeyBoolean from BOPDS;   
    ---C++: inline 
     
    Create(Other:PassKeyBoolean from BOPDS) 
    	returns PassKeyBoolean from BOPDS; 
    ---C++: inline 

    SetFlag(me:out; 
    	    theFlag: Boolean from Standard);  
    ---C++: inline 
    ---C++: alias "BOPDS_PassKeyBoolean& operator =(const BOPDS_PassKeyBoolean& );"  
     
    Flag(me)  
    	returns Boolean from Standard;   
    ---C++: inline  

fields
    myFlag: Boolean from Standard is protected; 

end PassKeyBoolean;
