-- Created on: 1996-04-12
-- Created by: Philippe MANGIN
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MinimalVariation from DrawFairCurve inherits Batten from DrawFairCurve

	---Purpose: Interactive Draw object of type "MVC"

uses MinimalVariation from FairCurve

is
   Create(TheMVC : Address)
   returns mutable MinimalVariation from DrawFairCurve;
   
   SetCurvature(me: mutable; Side : Integer; Rho : Real);
   SetPhysicalRatio(me: mutable; Ratio : Real);
   GetCurvature(me; Side : Integer) returns Real;
   GetPhysicalRatio(me) returns Real;
   FreeCurvature(me: mutable; Side : Integer);

end MinimalVariation;


