-- Created on: 1997-04-28
-- Created by: Christian CAILLET
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MakeTransformed  from StepToTopoDS    inherits Root

    ---Purpose : Produces instances by Transformation of a basic item

uses Trsf from gp, Shape from TopoDS,
     TransientProcess from Transfer,
     Axis2Placement3d from StepGeom,
     CartesianTransformationOperator3d from StepGeom,
     MappedItem       from StepRepr

is

    Create returns MakeTransformed;

    Compute (me : in out; Origin, Target : Axis2Placement3d from StepGeom)
    	returns Boolean;
    ---Purpose : Computes a transformation to pass from an Origin placement to
    --           a Target placement. Returns True when done
    --           If not done, the transformation will by Identity

    Compute (me : in out; Operator : CartesianTransformationOperator3d from StepGeom)  returns Boolean;
    ---Purpose : Computes a transformation defined by an operator 3D

    Transformation (me) returns Trsf from gp;
    ---Purpose : Returns the computed transformation (Identity if not yet or
    --           if failed)
    ---C++ : return const &

    Transform      (me; shape : in out Shape from TopoDS) returns Boolean;
    ---Purpose : Applies the computed transformation to a shape
    --           Returns False if the transformation is Identity


    TranslateMappedItem (me : in out; mapit : MappedItem from StepRepr;
    	    	    	 TP : TransientProcess from Transfer)
    	returns Shape;
    ---Purpose : Translates a MappedItem. More precisely
    --           A MappedItem has a MappingSource and a MappingTarget
    --           MappingSource has a MappedRepresentation and a MappingOrigin
    --           MappedRepresentation is the basic item to be instanced
    --           MappingOrigin is the starting placement
    --           MappingTarget is the final placement
    --           
    --           Hence, the transformation from MappingOrigin and MappingTarget
    --           is computed, the MappedRepr. is converted to a Shape, then
    --           transformed as an instance of this Shape

fields

    theTrsf : Trsf from gp;

end MakeTransformed;
