-- Created on: 2000-05-10
-- Created by: Andrey BETENEV
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1

class GroupRelationship from StepBasic
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity GroupRelationship

uses
    HAsciiString from TCollection,
    Group from StepBasic

is
    Create returns GroupRelationship from StepBasic;
	---Purpose: Empty constructor

    Init (me: mutable; aName: HAsciiString from TCollection;
                       hasDescription: Boolean;
                       aDescription: HAsciiString from TCollection;
                       aRelatingGroup: Group from StepBasic;
                       aRelatedGroup: Group from StepBasic);
	---Purpose: Initialize all fields (own and inherited)

    Name (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Name
    SetName (me: mutable; Name: HAsciiString from TCollection);
	---Purpose: Set field Name

    Description (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Description
    SetDescription (me: mutable; Description: HAsciiString from TCollection);
	---Purpose: Set field Description
    HasDescription (me) returns Boolean;
	---Purpose: Returns True if optional field Description is defined

    RelatingGroup (me) returns Group from StepBasic;
	---Purpose: Returns field RelatingGroup
    SetRelatingGroup (me: mutable; RelatingGroup: Group from StepBasic);
	---Purpose: Set field RelatingGroup

    RelatedGroup (me) returns Group from StepBasic;
	---Purpose: Returns field RelatedGroup
    SetRelatedGroup (me: mutable; RelatedGroup: Group from StepBasic);
	---Purpose: Set field RelatedGroup

fields
    theName: HAsciiString from TCollection;
    theDescription: HAsciiString from TCollection; -- optional
    theRelatingGroup: Group from StepBasic;
    theRelatedGroup: Group from StepBasic;
    defDescription: Boolean; -- flag "is Description defined"

end GroupRelationship;
