-- Created on: 1995-03-22
-- Created by: Laurent BUCHARD
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class FClass2d from BRepTopAdaptor

uses  
    Pnt2d             from gp,
    Face              from TopoDS,
    State             from TopAbs,
    SequenceOfInteger from TColStd,
    SeqOfPtr          from BRepTopAdaptor    

is 

    Create(F: Face from TopoDS; Tol: Real from Standard)
    returns FClass2d from BRepTopAdaptor;

    
    PerformInfinitePoint(me) 
    returns State from TopAbs;
    
    Perform(me; Puv: Pnt2d from gp; RecadreOnPeriodic: Boolean from Standard  =  Standard_True) 
    returns State from TopAbs;
    
    Destroy(me: in out);
    	---C++: alias ~
    

    Copy(me; Other: FClass2d from BRepTopAdaptor)
    returns FClass2d from BRepTopAdaptor;
    	---C++: return const &
      	---C++: alias operator=
     --Purpose *** Raise if called ***


    TestOnRestriction(me; Puv: Pnt2d from gp; 
                          Tol: Real from Standard;
                          RecadreOnPeriodic: Boolean from Standard  =  Standard_True) 
    returns State from TopAbs;
    ---Purpose: Test a point with +- an offset (Tol) and returns
    --          On if some points are OUT an some are IN
    --          (Caution: Internal use . see the code for more details)




fields 

    TabClass    : SeqOfPtr          from BRepTopAdaptor;
    TabOrien    : SequenceOfInteger from TColStd;
    Toluv       : Real              from Standard;
    Face        : Face              from TopoDS;
    U1          : Real              from Standard;
    V1          : Real              from Standard;    
    U2          : Real              from Standard;
    V2          : Real              from Standard;
    
    Umin        : Real              from Standard;  
    Umax        : Real              from Standard;
    Vmin        : Real              from Standard;  
    Vmax        : Real              from Standard;


end FClass2d from BRepTopAdaptor;
