-- File:        SurfaceStyleParameterLine.cdl
-- Created:     Mon Dec  4 12:02:31 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWSurfaceStyleParameterLine from RWStepVisual

	---Purpose : Read & Write Module for SurfaceStyleParameterLine

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     SurfaceStyleParameterLine from StepVisual,
     EntityIterator from Interface

is

	Create returns RWSurfaceStyleParameterLine;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable SurfaceStyleParameterLine from StepVisual);

	WriteStep (me; SW : in out StepWriter; ent : SurfaceStyleParameterLine from StepVisual);

	Share(me; ent : SurfaceStyleParameterLine from StepVisual; iter : in out EntityIterator);

end RWSurfaceStyleParameterLine;
