-- Created on: 1995-03-15
-- Created by: Laurent PAINNOT
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PolygonOnClosedSurface from BRep

    inherits PolygonOnSurface from BRep
    
    	---Purpose: Representation by two 2d polygons in the parametric
	--          space of a surface.

uses Polygon2D           from Poly,
     Surface             from Geom,
     CurveRepresentation from BRep,
     Location            from TopLoc



is
    Create(P1: Polygon2D from Poly;
    	   P2: Polygon2D from Poly;
    	   S:  Surface   from Geom;
	   L:  Location  from TopLoc)
    returns mutable PolygonOnClosedSurface from BRep;
    
    
    IsPolygonOnClosedSurface(me) returns Boolean
    	---Purpose: returns True.
    is redefined;

    Polygon2(me) returns any Polygon2D from Poly
    	---C++: return const&
    is redefined;

    Polygon2(me: mutable; P: Polygon2D from Poly)
    is redefined;
    
    
    Copy(me) returns mutable CurveRepresentation from BRep
	---Purpose: Return a copy of this representation.
    is redefined;
    
fields

myPolygon2: Polygon2D from Poly;

end PolygonOnClosedSurface;
