-- Created on: 1998-04-17
-- Created by: Andre LIEUTIER
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class  HPG0Constraint  from  NLPlate  inherits  HGPPConstraint from  NLPlate 
---Purpose: define a PinPoint G0  Constraint  used to load a Non Linear
--          Plate
uses
     XY from gp,
     XYZ from gp
     
is
    Create(UV : XY; Value : XYZ) returns mutable HPG0Constraint;
    -- create a G0 Constraint
    -- 

    SetUVFreeSliding(me: mutable; UVFree : Boolean) 
    is  redefined;
    -- If True, allow the UV value to  be modified during optimization
    --  this  is meaningless (has  no  effect) on   non G0 Constraints
    -- default is False
    -- 
    -- 

    SetIncrementalLoadAllowed(me: mutable; ILA : Boolean) 
    is  redefined;
    -- If True, allow the Constraint to be loaded incrementally during optimization
    -- default is False
    -- 


    UVFreeSliding(me)  returns  Boolean 
    is  redefined;
    -- If True, allow the UV value to be modified during optimization
    -- default is False
    -- 

    IncrementalLoadAllowed(me)  returns  Boolean 
    is redefined;
    -- If True, allow the Constraint to be loaded incrementally during optimization
    -- default is False
    -- 

    ActiveOrder(me)  returns  Integer 
    is   redefined; 
    --  returns the constraint active  order, i.e. the maximum between
    --  -- the initial constraint i.e 0 (for G0 Constraints)
    --  
    -- 

    IsG0(me) returns Boolean 
    is  redefined;

    G0Target(me) returns XYZ 
    ---C++: return const &
    is   redefined; 

fields
    myXYZTarget : XYZ from gp;
    UVIsFree : Boolean;
    IncrementalLoadingAllowed : Boolean;
end;
