-- Created on: 1993-05-19
-- Created by: Laurent PAINNOT
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

generic class SurfLeastSquare from AppCont(Surface   as any;
    	    	    	    	           SurfTool  as any)
				           ---as TheSurfTool(Surface)

    ---Purpose:


uses  Matrix          from math,
      Vector          from math,
      Constraint      from AppParCurves,
      MultiCurve      from AppParCurves,
      BezierSurface   from Geom


raises NotDone        from StdFail, 
       OutOfRange     from Standard,
       DimensionError from Standard



is

    Create(Surf: Surface; U0, U1, V0, V1: Real; 
    	   FirstCons, LastUCons, LastVCons, LastCons: Constraint; 
    	   DegU, DegV: Integer; NbPoints: Integer = 12)
    	---Purpose: given a MultiLine, this algorithm computes the
    	--          approximation of a continous Surface into a bezier
    	--          Surface.
    	--          The algorithm minimizes the volume between the 
    	--          Surface Surf and the Bezier Surface doing the 
    	--          aproximation.
    	--          NbPoints * NbPoints are taken on the Surface Surf.
    	--          The Constraints are affected to the following points:
    	--          
    	--              U0, V0 |--|---|---|---|---|---|-----| U1, V0 
    	--              FirstCons |   |   |   |   |   |     | LastUCons
    	--                     |--|---|---|---|---|---|-----|
    	--                     |--|---|---|---|---|---|-----|
    	--                     |  |   |   |   |   |   |     |
    	--              U0, V1 |--|---|---|---|---|---|-----| U1, V1
    	--              LastVCons                             LastCons


    returns SurfLeastSquare from AppCont
    raises DimensionError from Standard;    


    
    IsDone(me)
    	---Purpose: returns True if all has been correctly done.

    returns Boolean
    is static;
    
    
    Value(me: in out)
    	---Purpose: returns the result of the approximation.
    	--          An exception is raised if NotDone.
    	---C++: return const &

    returns BezierSurface from Geom
    raises NotDone from StdFail
    is static;



    Error(me; F: in out Real; MaxE3d: in out Real)
    	---Purpose: F is the sum of the square errors at each of the 
    	--          NbPoints*NbPoints and MaxE3d is the maximum value 
    	--          of these errors.
    	--          An exception is raised if NotDone.

    raises NotDone from StdFail
    is static;



fields

Done:      Boolean;
SCU:       BezierSurface from Geom;
DegreU:    Integer;
DegreV:    Integer;
Nbdiscret: Integer;
nbP:       Integer;
PointsX:   Matrix;
PointsY:   Matrix;
PointsZ:   Matrix;
PolesX:    Vector;
PolesY:    Vector;
PolesZ:    Vector;
myUParam:  Vector;
myVParam:  Vector;
VBU:       Matrix;
VBV:       Matrix;

end SurfLeastSquare from AppCont;

