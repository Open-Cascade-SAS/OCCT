-- Created on: 2002-12-12
-- Created by: data exchange team
-- Copyright (c) 2002-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class ElementMaterial from StepElement
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity ElementMaterial

uses
    HAsciiString from TCollection,
    HArray1OfMaterialPropertyRepresentation from StepRepr

is
    Create returns ElementMaterial from StepElement;
	---Purpose: Empty constructor

    Init (me: mutable; aMaterialId: HAsciiString from TCollection;
                       aDescription: HAsciiString from TCollection;
                       aProperties: HArray1OfMaterialPropertyRepresentation from StepRepr);
	---Purpose: Initialize all fields (own and inherited)

    MaterialId (me) returns HAsciiString from TCollection;
	---Purpose: Returns field MaterialId
    SetMaterialId (me: mutable; MaterialId: HAsciiString from TCollection);
	---Purpose: Set field MaterialId

    Description (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Description
    SetDescription (me: mutable; Description: HAsciiString from TCollection);
	---Purpose: Set field Description

    Properties (me) returns HArray1OfMaterialPropertyRepresentation from StepRepr;
	---Purpose: Returns field Properties
    SetProperties (me: mutable; Properties: HArray1OfMaterialPropertyRepresentation from StepRepr);
	---Purpose: Set field Properties

fields
    theMaterialId: HAsciiString from TCollection;
    theDescription: HAsciiString from TCollection;
    theProperties: HArray1OfMaterialPropertyRepresentation from StepRepr;

end ElementMaterial;
