-- Created on: 1994-09-06
-- Created by: Yves FRICAUD
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class CurAndInf2d from Geom2dLProp inherits CurAndInf from LProp

	---Purpose: An algorithm for computing local properties of a curve.
    	-- These properties include:
    	-- - the maximum and minimum curvatures
    	-- - the inflection points.
    	--   A CurAndInf2d object provides the framework for:
    	-- - defining the curve to be analyzed
    	-- - implementing the computation algorithms
    	-- - consulting the results.
    
uses
    Curve       from Geom2d
is
    Create;
 
    	--- Purpose: Initializes the framework.
    	-- Note: The curve on which the local properties are
    	-- computed is defined using one of the following
    	-- functions: Perform, PerformCurExt or PerformInf.   
        
    Perform (me : in out; C : Curve)
    	---Purpose: For the curve C, Computes both the
    	--  inflection points and the maximum and minimum curvatures.
    is static;
    
    PerformCurExt (me : in out; C : Curve)
    	---Purpose: For the curve C, Computes the locals extremas of curvature.
    is static;
    
    PerformInf    (me : in out; C : Curve)
       	---Purpose: For the curve C, Computes the inflections.
        -- After computation, the following functions can be used:
    	-- - IsDone to check if the computation was successful
    	-- - NbPoints to obtain the number of computed particular points
    	-- - Parameter to obtain the parameter on the curve for
    	--   each particular point
    	-- - Type to check if the point is an inflection point or an
    	--   extremum of curvature of the curve C.
    	--   Warning
    	-- These functions can be used to analyze a series of
    	-- curves, however it is necessary to clear the table of
    	-- results between each computation.
    is static;
    
    IsDone (me) returns Boolean
    	---Purpose: True if the solutions are found. 
    is static;
     
fields
    isDone     : Boolean   from Standard;

end CurAndInf2d;
