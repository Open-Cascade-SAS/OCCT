-- File:	StepToTopoDS_TranslateEdgeLoop.cdl
-- Created:	Wed Mar 29 08:20:18 1995
-- Author:	Frederic MAUPAS
--		<fma@pronox>
---Copyright:	 Matra Datavision 1995


class TranslateEdgeLoop from StepToTopoDS
    inherits Root from StepToTopoDS
    
    ---Purpose:
    --         

uses

    FaceBound              from StepShape,
    Surface                from StepGeom,
    Tool                   from StepToTopoDS,
    TranslateEdgeLoopError from StepToTopoDS,
    Shape                  from TopoDS,
    Surface                from Geom,
    Face                   from TopoDS,
    NMTool                 from StepToTopoDS
    
raises NotDone from StdFail

is

    Create returns TranslateEdgeLoop;
    
    Create (FB     : FaceBound     from StepShape;
            F      : Face          from TopoDS;
            S      : Surface       from Geom;
            SS     : Surface       from StepGeom;
            ss     : Boolean       from Standard;
            T      : in out Tool   from StepToTopoDS;
            NMTool : in out NMTool from StepToTopoDS)
    	returns TranslateEdgeLoop;
	    
    Init (me     : in out;
          FB     : FaceBound     from StepShape;
          F      : Face          from TopoDS;
          S      : Surface       from Geom;
          SS     : Surface       from StepGeom;
          ss     : Boolean       from Standard;
          T      : in out Tool   from StepToTopoDS;
          NMTool : in out NMTool from StepToTopoDS);

    Value (me) returns Shape from TopoDS
    	raises NotDone
	is static;
	---C++: return const &

    Error (me) returns TranslateEdgeLoopError from StepToTopoDS;
    
fields

    myError  : TranslateEdgeLoopError  from StepToTopoDS;
    
    myResult : Shape               from TopoDS;
    
end TranslateEdgeLoop;
