-- Created on: 2003-03-18
-- Created by: Oleg FEDYAEV
-- Copyright (c) 2003-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Tool from GeomLib

---Purpose:   The methods of this class compute the parameter(s) of a given point on a
-- curve or a surface. The point must be located either
-- on the curve (surface) itself or relatively to the latter at
-- a distance less than the tolerance value.
-- Return FALSE if the point is beyond the tolerance
-- limit or if computation fails.
-- Max Tolerance value is currently limited to 1.e-4 for
-- geometrical curves and 1.e-3 for BSpline, Bezier and
-- other parametrical curves.
        
uses Surface from Geom,
     Curve   from Geom,
     Curve   from Geom2d,
     Pnt     from gp,
     Pnt2d   from gp,
     Real    from Standard,
     Boolean from Standard
is

    Parameter(myclass; Curve     : in Curve from Geom;
    	    	       Point     : in Pnt   from gp;
		       Tolerance : in Real  from Standard;
		       U         : out Real from Standard)
     returns Boolean from Standard;
     ---Purpose: 
-- Extracts the parameter of a 3D point lying on a 3D curve
-- or at a distance less than the tolerance value.
     
    Parameters(myclass; Surface   : in Surface from Geom;
    	    	        Point     : in Pnt     from gp;
    	    	        Tolerance : in Real    from Standard;
     	    	        U         : out Real   from Standard;
    	    	    	V         : out Real   from Standard)
     returns Boolean from Standard;
     ---Purpose: Extracts the parameter of a 3D point lying on a surface
-- or at a distance less than the tolerance value. 
     
    Parameter(myclass; Curve     : in Curve from Geom2d;
    	    	       Point     : in Pnt2d from gp;
    	    	       Tolerance : in Real  from Standard;
     	    	       U         : out Real from Standard)
     returns Boolean from Standard;
     ---Purpose: Extracts the parameter of a 2D point lying on a 2D curve
-- or at a distance less than the tolerance value. 

end Tool;
