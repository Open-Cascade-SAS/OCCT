-- Created on: 1993-07-15
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Edge from DBRep inherits TShared from MMgt
	---Purpose: Display of an edge. Edge + color.
uses
    Edge    from TopoDS,
    Color   from Draw

is
    Create (E : Edge from TopoDS; C : Color from Draw)
    returns Edge from DBRep;
    
    Edge(me) returns Edge from TopoDS
	---C++: return const &
	---C++: inline
    is static;

    Edge(me : mutable; E : Edge from TopoDS)
	---C++: inline
    is static;

    Color(me) returns Color from Draw
	---C++: return const &
	---C++: inline
    is static;

    Color(me : mutable; C : Color from Draw)
	---C++: inline
    is static;

fields
    myEdge  : Edge  from TopoDS;
    myColor : Color from Draw;

end Edge;
