-- Created on: 1993-01-08
-- Created by: Philippe DAUTRY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package Sweep

    ---Purpose: This package contains generic classes usefull to create
    --          swept 3D primitives.

uses

    Standard, 
    TCollection, 
    TColStd,
    TopAbs

is
    
    --
    --     The following classes provides a directing topology for the
    --     LinearRegularSweep. This  is  the  topology of an  open  or
    --     closed loop of edges.
    --     

    class NumShape;

    class NumShapeTool;

    class NumShapeIterator;

end Sweep;


