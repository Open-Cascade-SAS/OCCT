-- Created on: 1994-07-19
-- Created by: Guest Kernel
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Convert from Quantity

    	---Purpose: Services to manage units conversion between Front-ends and Engines.
    	-- This conversion is managed by a table of correspondance between the quantities
    	-- and their "conversion coefficient".
    	-- This table is implemented like an external array (TCollection_Array1) regarding 
    	-- to the quantities enumeration.
     
uses 
    AsciiString from TCollection,
    PhysicalQuantity from Quantity,
    Coefficient from Quantity
	     
is

    Create returns Convert from Quantity;
    	---Purpose: Creates an object;

    SetQuantity(myclass ; 
                aQuantity : PhysicalQuantity from Quantity ;
	        aCoef: Coefficient from Quantity);	    
    	---Purpose: Updates the conversion table (correspondances between 
    	-- Quantities and conversion coefficients).
    	---C++: inline

    ConvertUserToSI(myclass ; 
                    aQuantity : PhysicalQuantity from Quantity ;
          	    aVal : Real from Standard)
    returns Real from Standard;
        ---Purpose: Converts, from the conversion table, the value <aVal>
    	-- from the user system to the SI system. 
    	---C++: inline

    ConvertSIToUser(myclass ; 
                    aQuantity : PhysicalQuantity from Quantity ;
          	    aVal : Real from Standard)
    returns Real from Standard;
    	---Purpose: Converts, from the conversion table, the value <aVal>
   	-- from the SI system to the user system. 
    	---C++: inline

    IsPhysicalQuantity(myclass; 
                       aTypeName : AsciiString from TCollection ; 
                       anEnum : in out AsciiString from TCollection)
    returns Boolean from Standard;
    	---Purpose:
    	-- if (aType is a physical quantity)
    	--    returns True and the name of the associated PhysicalQuantity .
    	-- else 
    	--    returns False.

end Convert from Quantity;
	        	







































































































