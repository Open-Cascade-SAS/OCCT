-- Created on: 1993-03-10
-- Created by: JCV
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



deferred class BoundedCurve from Geom inherits Curve from Geom


    	---Purpose : The abstract class BoundedCurve describes the
    	-- common behavior of bounded curves in 3D space. A
    	-- bounded curve is limited by two finite values of the
    	-- parameter, termed respectively "first parameter" and
    	-- "last parameter". The "first parameter" gives the "start
    	-- point" of the bounded curve, and the "last parameter"
    	-- gives the "end point" of the bounded curve.
    	-- The length of a bounded curve is finite.
    	-- The Geom package provides three concrete classes of bounded curves:
    	-- - two frequently used mathematical formulations of complex curves:
    	--   - Geom_BezierCurve,
    	--   - Geom_BSplineCurve, and
    	-- - Geom_TrimmedCurve to trim a curve, i.e. to only
    	--   take part of the curve limited by two values of the
    	--   parameter of the basis curve.


uses Pnt from gp

is

  EndPoint (me)   returns Pnt
        ---Purpose : Returns the end point of the curve.
     is deferred;


  StartPoint (me)  returns Pnt
        ---Purpose : Returns the start point of the curve.
     is deferred;


end;
