-- Created on: 1995-01-30
-- Created by: Mister rmi
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ModedPresentation from PrsMgr

uses
    Presentation from PrsMgr

is
    Create 
    returns  ModedPresentation from PrsMgr;
    
    Create(aPresentation:Presentation from PrsMgr;
           aMode: Integer from Standard) 
    returns  ModedPresentation from PrsMgr;
    
    Presentation(me) returns Presentation from PrsMgr
    is static;

    Mode(me) returns Integer from Standard;

    
fields

    myPresentation: Presentation from PrsMgr;
    myMode: Integer from Standard;
    
end ModedPresentation from PrsMgr;
    
