-- Created on: 1992-09-28
-- Created by: Remi GILET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class MakeRotation

from GC

    ---Purpose: This class implements elementary construction algorithms for a
    -- rotation in 3D space. The result is a
    -- Geom_Transformation transformation.
    -- A MakeRotation object provides a framework for:
    -- -   defining the construction of the transformation,
    -- -   implementing the construction algorithm, and
    -- -   consulting the result.

uses Pnt            from gp,
     Lin            from gp,
     Ax1            from gp,
     Dir            from gp,
     Transformation from Geom,
     Real           from Standard

is

Create(Line  : Lin from gp      ;
       Angle : Real  from Standard) returns MakeRotation;
    --- Purpose: Constructs a rotation through angle Angle about the axis defined by the line Line.
Create(Axis  : Ax1  from gp      ;
       Angle : Real from Standard) returns MakeRotation;
    ---Purpose: Constructs a rotation through angle Angle about the axis defined by the axis Axis.
Create(Point : Pnt  from gp      ;
       Direc : Dir  from gp      ; 
       Angle : Real from Standard) returns MakeRotation;
    ---Purpose: Constructs a rotation through angle Angle about the axis
    -- defined by the point Point and the unit vector Direc.
    
Value(me) returns Transformation from Geom
    is static;
    ---Purpose: Returns the constructed transformation.
    ---C++: return const&
  
Operator(me) returns Transformation from Geom
    is static;
    ---C++: return const&
    ---C++: alias "Standard_EXPORT operator Handle_Geom_Transformation() const;"

fields

    TheRotation : Transformation from Geom;

end MakeRotation;
