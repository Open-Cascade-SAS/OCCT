-- Created on: 1992-10-22
-- Created by: Gilles DEBARBOUILLE
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package Materials 

    ---Purpose: This package is useful  for creating Material objects,
    --          which contain a sequence of  physical properties.  All
    --          applications  which  request physical properties  on a
    --          given material, should reference this package.
    --          
    --          A predefined sequence  of materials  is given  by  the
    --          dictionary of  materials, and  the sequence   of known
    --          properties is given by the material definition.
    --          
    --          Only the  package  methods   are public,   except  the
    --          DictionaryOfMaterials class which   is called  by  the
    --          method Material.

uses

    TCollection,
    Quantity,
    Dynamic

is

    class Color; 
    class MaterialDefinition;    
    
    class MaterialsDictionary;    
    
    class FuzzyInstance instantiates FuzzyInstance from Dynamic(MaterialDefinition from Materials);
    
    class Material;
    
    class MtsSequence instantiates
          Sequence from TCollection (Material from Materials);
    class MaterialsSequence instantiates 
          HSequence from TCollection (Material from Materials, MtsSequence);
    
    MaterialFile(afile : CString from Standard); 
    ---Level: Public 
    ---Purpose: Sets the  location and the name  of the  file defining
    --          the definition of a material, in term of properties.
    
    MaterialsFile(afile : CString from Standard);
    ---Level: Public 
    ---Purpose: Sets  the location and  the name of  the file defining
    --          the dictionary of materials.
    
    MaterialsFile returns CString from Standard;   
    ---Level: Internal   
    ---Purpose: Returns  the location and the   name of the dictionary
    --          file of materials.
    
    DictionaryOfMaterials returns MaterialsDictionary from Materials; 
    ---Level: Internal 
    ---Purpose: Returns  the dictionary of materials.The dictionary is
    --          created at  the first call to this  method, or  if the
    --          dictionary is not up to date  with respect to the file
    --          date.
    
    ExistMaterial(aName : CString from Standard) returns Boolean from Standard;
    ---Purpose: True if the materialofname aName exists ...

    Material(amaterial : CString from Standard) returns Material from Materials;   
    ---Level: Public    
    ---Purpose: Retrieves from the dictionary the object material with
    --          <amaterial> as name.
    
    NumberOfMaterials returns Integer from Standard;   
    ---Level: Public   
    ---Purpose: Returns  the number of  materials previously stored in
    --          the dictionary.
    
    Material(anindex : Integer from Standard) returns Material from Materials;
    ---Level: Public 
    ---Purpose: This method used  with  the previous  one, allows  the
    --          exploration of    all the  dictionary.  It   returns a
    --          Material instance.
    
end Materials;








