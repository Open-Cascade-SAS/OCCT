-- Created on: 1995-12-07
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class Result from BRepCheck inherits TShared from MMgt

	---Purpose: 

uses Shape                                       from TopoDS,
     ListOfStatus                                from BRepCheck,
     DataMapOfShapeListOfStatus                  from BRepCheck,
     DataMapIteratorOfDataMapOfShapeListOfStatus from BRepCheck

raises NoSuchObject from Standard

is

    Initialize;

    Init(me: mutable; S: Shape from TopoDS);


    InContext(me: mutable; ContextShape: Shape from TopoDS)
    
    	is deferred;


    Minimum(me: mutable)
    
    	is deferred;

    
    Blind(me: mutable)
    
    	is deferred;

    SetFailStatus(me: mutable; S: Shape from TopoDS);


    Status(me)
    
    	returns ListOfStatus from BRepCheck
	---C++: return const&
	---C++: inline
	is static;

    IsMinimum(me)
    
    	returns Boolean from Standard
	---C++: inline
	is static;


    IsBlind(me)
    
    	returns Boolean from Standard
	---C++: inline
	is static;


    StatusOnShape(me: mutable; S: Shape from TopoDS)
	---Purpose: If  not  already   done,  performs the   InContext
	--          control and returns the list of status.
    	returns ListOfStatus from BRepCheck
	---C++: return const&
	raises
	    NoSuchObject from Standard
	is static;


    InitContextIterator(me: mutable)
    
    	is static;


    MoreShapeInContext(me)
    
    	returns Boolean from Standard
	---C++: inline
	is static;


    ContextualShape(me)
    
    	returns Shape from TopoDS
	---C++: return const&
	---C++: inline
	raises
	    NoSuchObject from Standard
	is static;


    StatusOnShape(me)
    
    	returns ListOfStatus from BRepCheck
	---C++: return const&
	---C++: inline
	raises
	    NoSuchObject from Standard
	is static;


    NextShapeInContext(me: mutable)
    
    	is static;


fields

    myShape : Shape                      from TopoDS    is protected;
    myMin   : Boolean                    from Standard  is protected;
    myBlind : Boolean                    from Standard  is protected;
    myMap   : DataMapOfShapeListOfStatus from BRepCheck is protected;
    myIter  : DataMapIteratorOfDataMapOfShapeListOfStatus from BRepCheck;

end Result;
