-- File:	StepShape_AngularLocation.cdl
-- Created:	Tue Apr 18 16:42:57 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0
-- Copyright:	Matra Datavision 1999

class AngularLocation from StepShape
inherits DimensionalLocation from StepShape

    ---Purpose: Representation of STEP entity AngularLocation

uses
    HAsciiString from TCollection,
    ShapeAspect from StepRepr,
    AngleRelator from StepShape

is
    Create returns AngularLocation from StepShape;
	---Purpose: Empty constructor

    Init (me: mutable; aShapeAspectRelationship_Name: HAsciiString from TCollection;
                       hasShapeAspectRelationship_Description: Boolean;
                       aShapeAspectRelationship_Description: HAsciiString from TCollection;
                       aShapeAspectRelationship_RelatingShapeAspect: ShapeAspect from StepRepr;
                       aShapeAspectRelationship_RelatedShapeAspect: ShapeAspect from StepRepr;
                       aAngleSelection: AngleRelator from StepShape);
	---Purpose: Initialize all fields (own and inherited)

    AngleSelection (me) returns AngleRelator from StepShape;
	---Purpose: Returns field AngleSelection
    SetAngleSelection (me: mutable; AngleSelection: AngleRelator from StepShape);
	---Purpose: Set field AngleSelection

fields
    theAngleSelection: AngleRelator from StepShape;

end AngularLocation;
