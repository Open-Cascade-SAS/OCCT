-- Created on: 1993-07-22
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



deferred class MakeOneAxis from BRepPrimAPI inherits MakeShape from BRepBuilderAPI

	---Purpose: The abstract class MakeOneAxis is the root class of
    	-- algorithms used to construct rotational primitives.

uses
    Address from Standard,
    Face    from TopoDS,
    Shell   from TopoDS,
    Solid   from TopoDS

raises
    NotDone     from StdFail

is
    OneAxis(me : in out) returns Address from Standard
	---Purpose: The inherited commands should provide the algorithm.
	--          Returned as a pointer.
	---Level: Public
    is deferred;
    
    Build(me : in out)
	---Purpose: Stores the solid in myShape.
	---Level: Public
    is redefined;

    Face(me : in out) 
	---Purpose: Returns the lateral face of the rotational primitive.
	--          
	---C++: return const &
	---C++: alias "Standard_EXPORT operator TopoDS_Face();" 
	---Level: Public
    returns Face from TopoDS
    is static;

    Shell(me : in out) 
	---Purpose: Returns the constructed rotational primitive as a shell.
    	---C++: return const &
	---C++: alias "Standard_EXPORT operator TopoDS_Shell();" 
    returns Shell from TopoDS
    is static;

    Solid(me : in out) 
	---Purpose: Returns the constructed rotational primitive as a solid.
	---C++: return const &
	---C++: alias "Standard_EXPORT operator TopoDS_Solid();" 
    returns Solid from TopoDS 
    is static;


end MakeOneAxis;
