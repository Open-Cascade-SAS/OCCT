-- Created on: 2005-04-18
-- Created by: Eugeny NAPALKOV <eugeny.napalkov@opencascade.com>
-- Copyright (c) 2005-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package BinMXCAFDoc

uses
    BinMDF,
    BinObjMgt,
    TopLoc,
    CDM,
    TDF,
    BinTools
is

    class AreaDriver;
    
    class CentroidDriver;
    
    class ColorDriver;
    
    class GraphNodeDriver;
    
    class LocationDriver;
    
    class VolumeDriver;
    
    class DatumDriver;
    class DimTolDriver;
    class MaterialDriver;
    
    class ColorToolDriver;
    class DocumentToolDriver;
    class LayerToolDriver;
    class ShapeToolDriver;
    class DimTolToolDriver;
    class MaterialToolDriver;

    AddDrivers (theDriverTable : ADriverTable  from BinMDF;
                theMsgDrv        : MessageDriver from CDM);
        ---Purpose: Adds the attribute drivers to <theDriverTable>.
end;
