-- Created on: 1996-04-05
-- Created by: Joelle CHAUVET
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


---Purpose : 
-- inherits class Cutting; contains a list of preferential points (di)i
-- if Cutting is necessary in [a,b], we cut at the di nearest from (a+b)/2.

class PrefCutting from AdvApprox inherits Cutting from AdvApprox

uses Array1OfReal from TColStd
    
is
    Create(CutPnts : Array1OfReal) returns PrefCutting;
    
    Value(me; a,b : Real;
              cuttingvalue : out Real)
    returns Boolean 
    is redefined;


fields

    myPntOfCutting : Array1OfReal from TColStd;


end PrefCutting;






























