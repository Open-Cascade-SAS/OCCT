-- Created on: 2018-03-15
-- Created by: Stephan GARNAUD (ARM)
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Printer from OSD 

 ---Purpose: Selects a printer (used by File).

uses Error, AsciiString from TCollection
raises ConstructionError, NullObject, OSDError

is
  Create (Name : AsciiString) returns Printer
   ---Purpose: Initializes printer to use with its name.
   --          The string must contain only ASCII characters
   --          between ' ' and '~'; this means no control character 
   --          and no extended ASCII code. If it is not the case the
   --          exception ConstructionError is raised.
   ---Level: Advanced
  raises ConstructionError;

  SetName (me : in out; Name : AsciiString)
  ---Purpose: Changes name of printer to use.
  ---Level: Advanced
  raises ConstructionError, NullObject is static;

  Name (me ;Name : out AsciiString) is static;
  ---Purpose: Returns name of current printer
  ---Level: Advanced

 Failed (me) returns Boolean is static;
  ---Purpose: Returns TRUE if an error occurs
  ---Level: Advanced

 Reset (me : in out) is static;
  ---Purpose: Resets error counter to zero
  ---Level: Advanced
      
 Perror (me : in out) 
  ---Level: Advanced
  ---Purpose: Raises OSD_Error
   raises OSDError is static;

 Error (me) returns Integer is static;
  ---Purpose: Returns error number if 'Failed' is TRUE.
  ---Level: Advanced

fields

  myName  : AsciiString;
  myError : Error;
end Printer from OSD;


