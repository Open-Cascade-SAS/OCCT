-- Created on: 1990-12-11
-- Created by: Remi Lequette
-- Copyright (c) 1990-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Update:      Frederic Maupas


class HShape from PTopoDS inherits ExternShareable from ObjMgt

    ---Purpose: The PTopoDS_HShape is the Persistent view of a TopoDS_Shape.
  -- This can be a vertex, an edge, a wire, a face, a shell, a solid and so on.
 -- It can be shared by other objects.
    --  a  HShape contains :
    --          
    --          - a reference to a TShape.
    --          
    --          - a Location  to put the TShape in  a local coordinate
    --          system.
    --          
    --          - an Orientation.
    --          
    --          It inherits from ExternShareable, so that it can be shared
    --          by other objects located outside the container.
    
uses

    Orientation   from TopAbs,
    TShape        from PTopoDS,
    Location      from PTopLoc
    
is
    Create returns mutable HShape from PTopoDS;
    ---Level: Internal 

    TShape(me) returns any TShape from PTopoDS
    ---Level: Internal 
    is static;

    TShape(me : mutable; T : TShape from PTopoDS)
    ---Level: Internal 
    is static;

    Location(me) returns Location from PTopLoc
    ---Level: Internal 
    is static;
	
    Location(me : mutable; L : Location from PTopLoc)
    ---Level: Internal 
    is static;
	
    Orientation(me) returns Orientation from TopAbs
    ---Level: Internal 
    is static;

    Orientation(me: mutable; O : Orientation from TopAbs)
    ---Level: Internal 
    is static;
    
fields
    myTShape   : TShape      from PTopoDS;
    myLocation : Location    from PTopLoc;
    myOrient   : Orientation from TopAbs;

end HShape;
