-- File:        MeasureQualification.cdl
-- Created:     Mon Dec  4 12:02:23 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWMeasureQualification from RWStepShape

	---Purpose : Read & Write Module for MeasureQualification

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     MeasureQualification from StepShape,
     EntityIterator from Interface

is

	Create returns RWMeasureQualification;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable MeasureQualification from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : MeasureQualification from StepShape);

	Share(me; ent : MeasureQualification from StepShape; iter : in out EntityIterator);

end RWMeasureQualification;
