-- Created on: 1993-01-09
-- Created by: CKY / Contract Toubro-Larsen ( Kiran )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Point from IGESGeom  inherits IGESEntity

        ---Purpose: defines IGESPoint, Type <116> Form <0>
        --          in package IGESGeom

uses

        SubfigureDef from IGESBasic,
        Pnt          from gp,
        XYZ          from gp
is

        Create returns Point;

        -- Specific Methods pertaining to the class

        Init (me : mutable; aPoint : XYZ; aSymbol : SubfigureDef);
        ---Purpose : This method is used to set the fields of the class Point
        --       - aPoint  : Coordinates of point
        --       - aSymbol : SubfigureDefinition entity specifying the
        --                   display symbol if there exists one, or zero

        Value (me) returns Pnt;
        ---Purpose : returns co-ordinates of the point

        TransformedValue (me) returns Pnt;
        ---Purpose : returns co-ordinates of the point after applying Transf. Matrix

        HasDisplaySymbol (me) returns Boolean;
        ---Purpose : returns True if symbol exists

        DisplaySymbol (me) returns SubfigureDef;
        ---Purpose : returns display symbol entity if it exists

fields

--
-- Class    : IGESGeom_Point
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class Point.
--
-- Reminder : A Point instance is defined by :
--            The coordinates of the point and display symbol if any

        thePoint  : XYZ;
        theSymbol : SubfigureDef;

end Point;
