-- Created on: 2004-05-11
-- Created by: Sergey ZARITCHNY <szy@opencascade.com>
-- Copyright (c) 2004-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package BinTools 

	---Purpose: Tool to keep shapes in binary format

uses 
    Geom2d, 
    Geom,
    TColStd,
    TopoDS, 
    TopAbs, 
    TopLoc,
    BRep,
    BRepTools, 
    TopTools
is
    
    class  ShapeSet; 

    class  Curve2dSet; 

    class  CurveSet;  

    class  SurfaceSet; 
     
    class  LocationSet;
    
    pointer LocationSetPtr to LocationSet from BinTools;


    PutReal (OS : out OStream from Standard; theValue : Real from Standard) returns OStream; 
    ---C++: return & 
    
    PutInteger (OS : out OStream from Standard; theValue : Integer from Standard) returns OStream;
    ---C++: return &  

    PutBool (OS : out OStream from Standard; theValue : Boolean from Standard) returns OStream;
    ---C++: return &  

    PutExtChar (OS : out OStream from Standard; theValue : ExtCharacter from Standard) returns OStream;
    ---C++: return &

    GetReal (IS : out IStream from Standard; theValue : out Real from Standard) returns IStream; 
    ---C++: return & 

    GetInteger (IS : out IStream from Standard; theValue : out Integer from Standard) returns IStream; 
    ---C++: return &  
     
    GetBool (IS : out IStream from Standard; theValue : out Boolean from Standard) returns IStream; 
    ---C++: return & 
     
    GetExtChar (IS : out IStream from Standard; theValue : out ExtCharacter from Standard) returns IStream; 
    ---C++: return &

end BinTools;

