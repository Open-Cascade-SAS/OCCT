-- Created by: Peter KURNEV
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class WireSplitter from BOPAlgo 
    	inherits Algo from BOPAlgo 
	 
	---Purpose: 

uses   
    Wire from TopoDS, 
    BaseAllocator from BOPCol, 
    ListOfShape from BOPCol, 
    WireEdgeSet from BOPAlgo,
    PWireEdgeSet from BOPAlgo, 
    ConnexityBlock from BOPTools, 
    ListOfConnexityBlock from BOPTools 
    
    
--raises

is 
    Create 
    	returns WireSplitter from BOPAlgo; 
    ---C++: alias "Standard_EXPORT virtual ~BOPAlgo_WireSplitter();" 
     
    Create(theAllocator: BaseAllocator from BOPCol)  
    	returns WireSplitter from BOPAlgo; 
     
    SetWES(me:out; 
    	    theWES: WireEdgeSet from BOPAlgo);  
    
    
    WES(me:out) 
    	returns WireEdgeSet from BOPAlgo; 
    ---C++:  return &  

    Perform(me:out) 
	is redefined; 
	 
    MakeWire(myclass; 
    	    theLE:out ListOfShape from BOPCol; 
    	    theW :out Wire from TopoDS);  
    ---C++: inline 
     
    CheckData(me:out) 
	is redefined protected;    
	
    MakeConnexityBlocks(me:out)  
    	is protected;  
     
    MakeWires(me:out)  
    	is protected;  
	 
    SplitBlock(me:out; 
    	    theCB:out ConnexityBlock from BOPTools)  
    	is protected; 
    
fields 
    myWES   : PWireEdgeSet from BOPAlgo is protected;
    myLCB   : ListOfConnexityBlock from BOPTools is protected; 
    
end WireSplitter;
