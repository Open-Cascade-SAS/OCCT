-- File:        SurfaceOfLinearExtrusion.cdl
-- Created:     Mon Dec  4 12:02:31 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWSurfaceOfLinearExtrusion from RWStepGeom

	---Purpose : Read & Write Module for SurfaceOfLinearExtrusion

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     SurfaceOfLinearExtrusion from StepGeom,
     EntityIterator from Interface

is

	Create returns RWSurfaceOfLinearExtrusion;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable SurfaceOfLinearExtrusion from StepGeom);

	WriteStep (me; SW : in out StepWriter; ent : SurfaceOfLinearExtrusion from StepGeom);

	Share(me; ent : SurfaceOfLinearExtrusion from StepGeom; iter : in out EntityIterator);

end RWSurfaceOfLinearExtrusion;
