-- Created on: 2002-10-29
-- Created by: Michael SAZONOV
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DocumentStorageDriver from BinDrivers inherits DocumentStorageDriver from BinLDrivers

    ---Purpose: persistent implemention of storage a document in a binary file

uses   
    OStream          from Standard,
    MessageDriver    from CDM, 
    DocumentSection  from BinLDrivers,
    ADriverTable     from BinMDF
is
    -- ===== Public methods =====

    Create returns DocumentStorageDriver from BinDrivers;
	---Purpose: Constructor


    AttributeDrivers  (me : mutable; theMsgDriver: MessageDriver from CDM)
	returns ADriverTable from BinMDF
	is redefined virtual; 
	 
    WriteShapeSection    (me: mutable; theDocSection : in out DocumentSection from BinLDrivers;
                                       theOS         : in out OStream from Standard)
        is redefined  virtual; 
        ---Purpose: implements the procedure of writing a shape section to file 	

end DocumentStorageDriver;
