-- Created on: 1997-01-24
-- Created by: Robert COUBLANC
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

private class GlobalStatus from AIS inherits TShared from MMgt

	---Purpose: Stores  information  about objects in graphic context:
	--          - Status Of Display : in the main viewer 
	--                                hidden in the main viewer
	--          - Displayed Modes 
	--          - Active Selection Modes
	--          - is the Interactive Object Current ?
	--          - Layer Index

uses 
    ListOfInteger from TColStd,
    DisplayStatus from AIS,
    NameOfColor from Quantity

is

    Create returns GlobalStatus from AIS;

    Create (aStat             : DisplayStatus from AIS;
    	    aDispMode,aSelMode: Integer from Standard;
	    ishilighted       : Boolean from Standard=Standard_False;
	    TheHiCol          : NameOfColor from Quantity = Quantity_NOC_WHITE;
	    aLayerIndex       : Integer from Standard = 0)
	    returns GlobalStatus from AIS;

		    ---Category: Modifications.

    SetGraphicStatus(me:mutable; aStat :  DisplayStatus from AIS);
    ---C++: inline
    AddDisplayMode(me:mutable; aMode: Integer from Standard);
    ---C++: inline    
    AddSelectionMode(me:mutable; aMode : Integer from Standard);
    ---C++: inline    
    SetLayerIndex (me: mutable ; AnIndex : Integer from Standard);
    ---C++: inline  
    SetHilightStatus (me: mutable; aStat:Boolean from Standard);
    ---C++: inline    
    SetHilightColor(me:mutable;aHiCol : NameOfColor from Quantity);
    ---C++: inline    



    IsSubIntensityOn(me) returns Boolean from Standard;
    ---C++: inline
    SubIntensityOn (me: mutable);
    ---C++: inline    
    SubIntensityOff (me: mutable);
    ---C++: inline    

    

    RemoveDisplayMode(me:mutable; aMode : Integer from Standard);

    RemoveSelectionMode(me:mutable; aMode : Integer from Standard);
    ClearSelectionModes(me:mutable);


 		    ---Category: Information.

   
    GraphicStatus(me) returns DisplayStatus from AIS;
    ---C++: inline
	    
    DisplayedModes(me) returns ListOfInteger from TColStd;
    ---C++: return const &
    ---C++: inline
    ---Purpose: keeps the information of displayed modes in the 
    --          main viewer.

    SelectionModes(me) returns ListOfInteger from TColStd;
    ---C++: return const &
    ---C++: inline
    ---Purpose: keeps the active selection modes of the object
    --          in the main viewer.

    IsHilighted(me) returns Boolean from Standard;
    ---C++: inline

    HilightColor(me) returns NameOfColor from Quantity;
    ---C++: inline

    IsDModeIn(me; aMode : Integer from Standard) returns Boolean from Standard;

    IsSModeIn(me; aMode : Integer from Standard) returns Boolean from Standard;
    
    
fields

    myStatus     : DisplayStatus from AIS;
    myDispModes  : ListOfInteger from TColStd;
    mySelModes   : ListOfInteger from TColStd;
    myLayerIndex : Integer       from Standard;
    myIsHilit    : Boolean       from Standard;
    myHiCol      : NameOfColor   from Quantity;
    mySubInt     : Boolean;
end GlobalStatus;
