-- Created on: 1994-09-02
-- Created by: Frederic MAUPAS
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MakeEllipse from GeomToStep inherits Root from GeomToStep

    ---Purpose: This class implements the mapping between classes 
    --          Ellipse from Geom, and Circ from gp, and the class
    --          Ellipse from StepGeom which describes a Ellipse from
    --          Prostep. 
  
uses Elips from gp,
     Elips2d from gp,
     Ellipse from Geom,
     Ellipse from Geom2d,
     Ellipse from StepGeom
     
raises NotDone from StdFail
     
is 

Create ( C : Elips from gp ) returns MakeEllipse;

Create ( C : Ellipse from Geom ) returns MakeEllipse;

Create ( C : Ellipse from Geom2d ) returns MakeEllipse;

Value (me) returns Ellipse from StepGeom
    raises NotDone
    is static;
    ---C++: return const&
  
fields

    theEllipse : Ellipse from StepGeom;
    	-- The solution from StepGeom
    	
end MakeEllipse;


