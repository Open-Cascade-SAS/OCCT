-- Created on: 1995-03-09
-- Created by: Laurent PAINNOT
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class Polygon2D from Poly inherits TShared from MMgt

    	---Purpose: Provides a polygon in 2D space (for example, in the
    	-- parametric space of a surface). It is generally an
    	-- approximate representation of a curve.
    	-- A Polygon2D is defined by a table of nodes. Each node is
    	-- a 2D point. If the polygon is closed, the point of closure is
    	-- repeated at the end of the table of nodes.


uses Array1OfPnt2d  from TColgp

raises NullObject from Standard

is

    Create(Nodes: Array1OfPnt2d from TColgp) 
    returns mutable Polygon2D from Poly;
    	---Purpose: Constructs a 2D polygon defined by the table of points, <Nodes>.
    
    Deflection(me) returns Real;
    	---Purpose: Returns the deflection of this polygon.
    	--  Deflection is used in cases where the polygon is an
    	-- approximate representation of a curve. Deflection
    	-- represents the maximum distance permitted between any
    	-- point on the curve and the corresponding point on the polygon.
    	-- By default the deflection value is equal to 0. An algorithm
    	-- using this 2D polygon with a deflection value equal to 0
    	-- considers that it is working with a true polygon and not with
    	-- an approximate representation of a curve. The Deflection
    	-- function is used to modify the deflection value of this polygon.
    	-- The deflection value can be used by any algorithm working  with 2D polygons.
    	-- For example:
    	-- -   An algorithm may use a unique deflection value for all
    	--   its polygons. In this case it is not necessary to use the
    	--   Deflection function.
    	-- -   Or an algorithm may want to attach a different
    	--   deflection to each polygon. In this case, the Deflection
    	--   function is used to set a value on each polygon, and
    	--   later to fetch the value.
    
    Deflection(me : mutable; D : Real);
    	---Purpose: Sets the deflection of this polygon to D    

    NbNodes(me) returns Integer;
	---Purpose: Returns the number of nodes in this polygon.
    	-- Note: If the polygon is closed, the point of closure is
    	-- repeated at the end of its table of nodes. Thus, on a closed
    	-- triangle, the function NbNodes returns 4.
    	---C++: inline

    Nodes(me) returns Array1OfPnt2d from TColgp
	---Purpose: Returns the table of nodes for this polygon.
	---C++: return const &
    raises NullObject from Standard;
    	
    
fields

    myDeflection: Real;
    myNbNodes:    Integer;
    myNodes:      Array1OfPnt2d from TColgp;

end Polygon2D;
