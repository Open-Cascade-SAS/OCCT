-- Created on: 2002-12-12
-- Created by: data exchange team
-- Copyright (c) 2002-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class UniformSurfaceSection from StepElement
inherits SurfaceSection from StepElement

    ---Purpose: Representation of STEP entity UniformSurfaceSection

uses
    MeasureOrUnspecifiedValue from StepElement

is
    Create returns UniformSurfaceSection from StepElement;
	---Purpose: Empty constructor

    Init (me: mutable; aSurfaceSection_Offset: MeasureOrUnspecifiedValue from StepElement;
                       aSurfaceSection_NonStructuralMass: MeasureOrUnspecifiedValue from StepElement;
                       aSurfaceSection_NonStructuralMassOffset: MeasureOrUnspecifiedValue from StepElement;
                       aThickness: Real;
                       aBendingThickness: MeasureOrUnspecifiedValue from StepElement;
                       aShearThickness: MeasureOrUnspecifiedValue from StepElement);
	---Purpose: Initialize all fields (own and inherited)

    Thickness (me) returns Real;
	---Purpose: Returns field Thickness
    SetThickness (me: mutable; Thickness: Real);
	---Purpose: Set field Thickness

    BendingThickness (me) returns MeasureOrUnspecifiedValue from StepElement;
	---Purpose: Returns field BendingThickness
    SetBendingThickness (me: mutable; BendingThickness: MeasureOrUnspecifiedValue from StepElement);
	---Purpose: Set field BendingThickness

    ShearThickness (me) returns MeasureOrUnspecifiedValue from StepElement;
	---Purpose: Returns field ShearThickness
    SetShearThickness (me: mutable; ShearThickness: MeasureOrUnspecifiedValue from StepElement);
	---Purpose: Set field ShearThickness

fields
    theThickness: Real;
    theBendingThickness: MeasureOrUnspecifiedValue from StepElement;
    theShearThickness: MeasureOrUnspecifiedValue from StepElement;

end UniformSurfaceSection;
