-- Created on: 1996-04-09
-- Created by: Yves FRICAUD
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Collect from BRepBuilderAPI 

	---Purpose: 

uses
    Shape                     from TopoDS,
    DataMapOfShapeListOfShape from TopTools,
    MapOfShape                from TopTools,
    MakeShape                 from BRepBuilderAPI
    
is

    Create returns Collect from BRepBuilderAPI;
    
    Add  (me : in out; SI  : Shape            from TopoDS  ;
		       MKS : in out MakeShape from BRepBuilderAPI );
    	---Purpose: 
   
    AddGenerated  (me : in out; S   : Shape from TopoDS  ;  
		                 Gen : Shape from TopoDS  );
       ---Purpose:

    AddModif  (me : in out; S      : Shape from TopoDS  ;  
		             Mod    : Shape from TopoDS  ); 
       ---Purpose: 
		   
    Filter     (me : in out; SF : Shape from TopoDS  );
	---Purpose: 

    Modification (me) returns DataMapOfShapeListOfShape from TopTools;
    ---C++: return const &

    Generated    (me) returns DataMapOfShapeListOfShape from TopTools;
    ---C++: return const &
    
    
fields
    myInitialShape : Shape from TopoDS;
    myDeleted      : MapOfShape from TopTools;
    myMod          : DataMapOfShapeListOfShape from TopTools;
    myGen          : DataMapOfShapeListOfShape from TopTools;
end Collect;
