-- Created by: DAUTRY Philippe
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

--      	--------------

---Version:	0.0
--Version	Date		Purpose
--		0.0	Sep 17 1997	Creation


class XLink from PDocStd inherits Attribute from PDF

	---Purpose: This attribute define a persistant external link.

uses

    HAsciiString from PCollection

-- raises

is

    Create
    returns XLink from PDocStd;
    ---Purpose: Returns an empty persistent external reference.


    DocumentEntry(me : mutable; aDocEntry : HAsciiString from PCollection);
    ---Purpose: Sets the field <myDocEntry> with <aDocEntry>.
    
    DocumentEntry(me)
    returns HAsciiString from PCollection;
    ---Purpose: Returns the contents of the field <myDocEntry>.

    LabelEntry(me : mutable; aLabEntry : HAsciiString from PCollection);
    ---Purpose: Sets the field <myLabEntry> with <aLabEntry>.

    LabelEntry(me)
    returns HAsciiString from PCollection;
    ---Purpose: Returns the contents of the field <myLabEntry>.


fields

    myDocEntry       : HAsciiString from PCollection;
    myLabEntry       : HAsciiString from PCollection;

end XLink from PDocStd;
