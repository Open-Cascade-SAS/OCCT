-- Created on: 1994-08-26
-- Created by: Frederic MAUPAS
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MakeAxisPlacement from StepToGeom

    ---Purpose: This class implements the mapping between classes 
    --          Axis2Placement2d from Step and AxisPlacement from Geom2d

uses AxisPlacement from Geom2d,
     Axis2Placement2d from StepGeom
     
is 

    Convert ( myclass; SA : Axis2Placement2d from StepGeom;
                       CA : out AxisPlacement from Geom2d )
    returns Boolean from Standard;

end MakeAxisPlacement;
