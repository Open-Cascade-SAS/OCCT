-- Created on: 2009-04-06
-- Created by: Sergey ZARITCHNY
-- Copyright (c) 2009-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Shape from TDataXtd inherits Attribute from TDF

	---Purpose: A Shape is associated in the framework with :
	--          a NamedShape attribute 


uses Attribute       from TDF,
     Label           from TDF,
     NamedShape      from TNaming,
     GUID            from Standard,
     DataSet         from TDF,
     RelocationTable from TDF,
     Shape           from TopoDS
is    


    ---Purpose: class methods
    --          =============
    
    Find (myclass; current : Label from TDF; S : in out Shape from TDataXtd)
    ---Purpose: try to retrieve a Shape attribute at <current> label
    --           or in  fathers  label of  <current>. Returns True  if
    --          found and set <S>.
    returns Boolean from Standard;
    
    New (myclass; label : Label from TDF)
    ---Purpose: Find, or create, a Shape attribute.  the Shape attribute
    --          is returned. Raises if <label> has attribute.
    returns Shape from TDataXtd;

    Set (myclass; label : Label from TDF; shape : Shape from TopoDS)
    ---Purpose: Create or update associated NamedShape attribute.  the
    --          Shape attribute is returned.
    returns Shape from TDataXtd;    

    Get (myclass; label : Label from TDF)
    ---Purpose:   the Shape from  associated NamedShape attribute
    --            is returned.
    returns Shape from TopoDS;
    
    GetID (myclass)   
    ---C++: return const &  
    returns GUID from Standard;

    ---Purpose: Shape methods
    --          ============

    Create
    returns mutable Shape from TDataXtd;

    
    ---Category: methodes de TDF_Attribute
    --           =========================
 
	
    ID (me)
    ---C++: return const & 
    returns GUID from Standard;

    Restore (me: mutable; with : Attribute from TDF);

    NewEmpty (me)
    returns mutable Attribute from TDF;

    Paste (me; into : mutable Attribute from TDF;
	       RT   : mutable RelocationTable from TDF);       

    References (me; DS : DataSet from TDF) is redefined;   

    Dump(me; anOS : in out OStream from Standard)
    returns OStream from Standard
     is redefined;
	---C++: return &

end Shape;

