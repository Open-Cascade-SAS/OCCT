-- Created on: 2001-12-13
-- Created by: Peter KURNEV
-- Copyright (c) 2001-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PntOn2Faces from IntTools 

	---Purpose: Contains two points PntOnFace from IntTools and a flag

uses
    PntOnFace from IntTools
---raises

is 
    Create 
    	returns PntOn2Faces from IntTools; 
	---Purpose:
	--- Empty constructor
	---
	 
    Create(aP1:	PntOnFace from IntTools;
           aP2:	PntOnFace from IntTools);
    	---Purpose:
	--- Initializes me by two points aP1 and aP2
	---
	    
    SetP1 (me:out; 
    	aP1: PntOnFace from IntTools);
	---Purpose:
	--- Modifier
	---
	 
    SetP2 (me:out; 
    	aP2: PntOnFace from IntTools);
	---Purpose:
	--- Modifier
	---

    SetValid(me:out; 
	bF : Boolean from Standard); 
	---Purpose:
	--- Modifier
	---
     
    P1(me) 
    	returns PntOnFace from IntTools; 
    	---C++:  return const &  
	---Purpose:
	--- Selector
	---
     
    P2(me) 
    	returns PntOnFace from IntTools; 
    	---C++:  return const & 
	---Purpose:
	--- Selector
	---

    IsValid(me) 
	returns Boolean from Standard; 
	---Purpose:
	--- Selector
	---

fields
  
    myIsValid : Boolean from Standard;    
    myPnt1    : PntOnFace from IntTools;
    myPnt2    : PntOnFace from IntTools;
    
     
end PntOn2Faces;
