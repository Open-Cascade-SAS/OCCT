-- Created on: 1993-01-11
-- Created by: CKY / Contract Toubro-Larsen ( Arun MENON )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ReferenceDesignator from IGESAppli  inherits IGESEntity

        ---Purpose: defines ReferenceDesignator, Type <406> Form <7>
        --          in package IGESAppli
        --          Used to attach a text string containing the value of
        --          a component reference designator to an entity being
        --          used to represent a component.

uses

        HAsciiString from TCollection

is

        Create returns mutable ReferenceDesignator;

        -- Specific Methods pertaining to the class

        Init (me        : mutable; 
              nbPropVal : Integer; 
              aText     : HAsciiString);
        ---Purpose : This method is used to set the fields of the class
        --           ReferenceDesignator
        --       - nbPropVal : Number of property values = 1
        --       - aText     : Reference designator text

        NbPropertyValues (me) returns Integer;
        ---Purpose : returns the number of property values
        -- is always 1

        RefDesignatorText (me) returns HAsciiString from TCollection;
        ---Purpose : returns the Reference designator text

fields

--
-- Class    : IGESAppli_ReferenceDesignator
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class ReferenceDesignator.
--
-- Reminder : A ReferenceDesignator instance is defined by :
--            - Number of property values (always = 1)
--            - Reference designator text

        theNbPropertyValues : Integer;
        theRefDesigText     : HAsciiString;

end ReferenceDesignator;
