-- File:	QANewBRepNaming_Fillet.cdl
-- Created:	Fri Oct  8 09:09:14 1999
-- Author:	Vladislav ROMASHKO
--		<v-romashko@opencascade.com>
---Copyright:	 Open CASCADE 2003

class Fillet from QANewBRepNaming inherits TopNaming from QANewBRepNaming

	---Purpose: For topological naming of a fillet

uses

     MakeFillet from BRepFilletAPI,
     Shape      from TopoDS,
     Label      from TDF

is

    Create returns Fillet from QANewBRepNaming;

    Create(ResultLabel : Label from TDF)
    returns Fillet from QANewBRepNaming;

    Init(me : in out; ResultLabel : Label from TDF);


    Load (me; part     :        Shape      from TopoDS;
    	      mkFillet : in out MakeFillet from BRepFilletAPI);
      ---Purpose: Loads a fillet in a data framework

    DeletedFaces(me)
    ---Purpose: Returns a label for deleted faces of the part.
    returns Label from TDF;

    ModifiedFaces(me)
    ---Purpose: Returns a label for modified faces of the part.
    returns Label from TDF;

    FacesFromEdges(me)
    ---Purpose: Returns a label for faces generated from edges of the part.
    returns Label from TDF;

    FacesFromVertices(me)
    ---Purpose: Returns a label for faces generated from vertices of the part.
    returns Label from TDF;

    WRFace1(me)
    ---Purpose: Returns a label for WorkAround Face number 1
    returns Label from TDF;

    WRFace2(me)
    ---Purpose: Returns a label for WorkAround Face number 2
    returns Label from TDF;

    WREdge1(me)
    ---Purpose: Returns a label for WorkAround Edge number 1
    returns Label from TDF;

    WREdge2(me)
    ---Purpose: Returns a label for WorkAround Edge number 2
    returns Label from TDF;


end Fillet;
