-- Created on: 1993-09-21
-- Created by: Christian CAILLET
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class ToolLocation  from IGESData  inherits TShared

    ---Purpose : This Tool determines and gives access to effective Locations
    --           of IGES Entities as defined by the IGES Norm. These Locations
    --           can be for each Entity :
    --           - on one part, explicitly defined by a Transf in Directory
    --             Part (this Transf can be itself compound); if not defined,
    --             no proper Transformation is defined
    --           - on the other part, implicitly defined by a reference from
    --             another Entity : its Parent
    --           Both implicit and explicit locations are combinable.
    --           
    --           Implicit definition can be itself defined, either through the
    --           definition of an Entity (i.e. a Composite Curve references
    --           a list of Curves), or by a specific Associativity, of type
    --           SingleParentEntity, by which the Location of the Parent is
    --           applied to the Childs defined by this Associativity.
    --           Remark that a Transf itself has no Location, but it can be
    --           compound
    --           
    --           This is a TShared object, then it is easier to use in an
    --           interactive session


uses GTrsf from gp, Trsf from gp, Array1OfInteger from TColStd,
     GeneralLib, IGESEntity, IGESModel, Protocol from IGESData

raises DomainError

is

    Create (amodel : IGESModel; protocol : Protocol from IGESData)
    	returns mutable ToolLocation;
    ---Purpose : Creates a ToolLocation on a given Model, filled with the help
    --           of a Protocol (which allows to known Entities referenced by
    --           other ones)

    Load (me : mutable);
    ---Purpose : Does the effective work of determining Locations of Entities

    SetPrecision (me : mutable; prec : Real) is static;
    ---Purpose : Sets a precision for the Analysis of Locations
    --           (default by constructor is 1.E-05)

    	-- --    Internal Actions to Compute and Edit the Result    -- --

    SetReference      (me : mutable; parent, child : IGESEntity)  is static;
    ---Purpose : Sets the "Reference" information for <child> as being <parent>
    --           Sets an Error Status if already set (see method IsAmbiguous)

    SetParentAssoc    (me : mutable; parent, child : IGESEntity)  is static;
    ---Purpose : Sets the "Associativity" information for <child> as being
    --           <parent> (it must be the Parent itself, not the Associativity)

    ResetDependences  (me : mutable; child : IGESEntity)  is static;
    ---Purpose : Resets all informations about dependences for <child>

    SetOwnAsDependent (me : mutable; ent : IGESEntity);
    ---Purpose : Unitary action which defines Entities referenced by <ent>
    --           (except those in Directory Part and Associativities List)
    --           as Dependent (their Locations are related to that of <ent>)

    	-- --    Queries  -- --

    IsTransf         (me; ent : IGESEntity) returns Boolean  is static;
    ---Purpose : Returns True if <ent> is kind of TransfEntity. Then, it has
    --           no location, while it can be used to define a Location)

    IsAssociativity  (me; ent : IGESEntity) returns Boolean  is static;
    ---Purpose : Returns True if <ent> is an Associativity (IGES Type 402).
    --           Then, Location does not apply.

    HasTransf        (me; ent : IGESEntity) returns Boolean  is static;
    ---Purpose : Returns True if <ent> has a Transformation Matrix in proper
    --           (referenced from its Directory Part)

    ExplicitLocation (me; ent : IGESEntity) returns GTrsf from gp  is static;
    ---Purpose : Returns the Explicit Location defined by the Transformation
    --           Matrix of <ent>. Identity if there is none


    IsAmbiguous      (me; ent : IGESEntity) returns Boolean  is static;
    ---Purpose : Returns True if more than one Parent has been determined for
    --           <ent>, by adding direct References and Associativities

    HasParent        (me; ent : IGESEntity) returns Boolean
    ---Purpose : Returns True if <ent> is dependent from one and only one other
    --           Entity, either by Reference or by Associativity
    	raises DomainError  is static;
    --           Error if more than one Parent has been noted

    Parent           (me; ent : IGESEntity) returns IGESEntity
    ---Purpose : Returns the unique Parent recorded for <ent>.
    --           Returns a Null Handle if there is none
    	raises DomainError  is static;
    --           Error if more than one Parent has been noted

    HasParentByAssociativity (me; ent : IGESEntity) returns Boolean
    ---Purpose : Returns True if the Parent, if there is one, is defined by
    --           a SingleParentEntity Associativity
    --           Else, if HasParent is True, it is by Reference
    	raises DomainError  is static;
    --           Error if more than one Parent has been noted

    ParentLocation    (me; ent : IGESEntity) returns GTrsf from gp
    ---Purpose : Returns the effective Location of the Parent of <ent>, if
    --           there is one : this Location is itself given as compound
    --           according dependences on the Parent, if there are some.
    --           Returns an Identity Transformation if no Parent is recorded.
    	raises DomainError  is static;
    --           Error if more than one Parent has been noted

    EffectiveLocation (me; ent : IGESEntity) returns GTrsf from gp
    ---Purpose : Returns the effective Location of an Entity, i.e. the
    --           composition of its proper Transformation Matrix (returned by
    --           Transf) and its Parent's Location (returned by ParentLocation)
    	raises DomainError  is static;
    --           Error if more than one Parent has been noted

    AnalyseLocation (me; loc : GTrsf from gp; result : out Trsf from gp)
    	returns Boolean  is static;
    ---Purpose : Analysis a Location given as a GTrsf, by trying to convert it
    --           to a Trsf (i.e. to a True Location of which effect is
    --           described by an Isometry or a Similarity)
    --           Works with the Precision given by default or by SetPrecision
    --           Calls ConvertLocation (see below)

    ConvertLocation (myclass; prec : Real;
    	     loc : GTrsf from gp; result : out Trsf from gp; uni : Real = 1)
     returns Boolean;
    ---Purpose : Convertion of a Location, from GTrsf form to Trsf form
    --           Works with a precision given as argument.
    --           Returns True if the Conversion is possible, (hence, <result>
    --           contains the converted location), False else
    --           <unit>, if given, indicates the unit in which <loc> is defined
    --           in meters. It concerns the translation part (to be converted.
    --           
    --           As a class method, it can be called separately


fields

    theprec   : Real;
    themodel  : IGESModel;
    thelib    : GeneralLib;
    therefs   : Array1OfInteger from TColStd;
    theassocs : Array1OfInteger from TColStd;

end ToolLocation;
