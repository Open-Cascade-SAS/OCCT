-- Created on: 1991-04-03
-- Created by: Remi GILET
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Lin2d2Tan

from GccAna

	---Purpose: This class implements the algorithms used to 
	--          create 2d lines tangent to 2 other elements which
	--          can be circles or points.
    	--          Describes functions for building a 2D line:
    	--          -   tangential to 2 circles, or
    	--          -   tangential to a circle and passing through a point, or
    	--          -   passing through 2 points.
    	--          A Lin2d2Tan object provides a framework for:
    	--          -   defining the construction of 2D line(s),
    	--          -   implementing the construction algorithm, and 
        --          consulting the result(s).
    	--          Some constructors may check the type of the qualified argument 
    	--          and raise BadQualifier Error in case of incorrect couple (qualifier,
    	--          curv).
    	--          For example: "EnclosedCirc".

uses Pnt2d         from gp, 
     Lin2d         from gp,
     QualifiedCirc from GccEnt,
     Array1OfLin2d from TColgp,
     Array1OfPnt2d from TColgp,
     Array1OfReal  from TColStd,
     Position         from GccEnt,
     Array1OfPosition from GccEnt
     

raises OutOfRange   from Standard,
       BadQualifier from GccEnt,
       NotDone      from StdFail

is



Create (ThePoint1  : Pnt2d         from gp      ;
        ThePoint2  : Pnt2d         from gp      ;
        Tolerance  : Real          from Standard) returns Lin2d2Tan;
	---Purpose: This methods implements the algorithms used to 
	--          create 2d lines passing thrue 2 points.
	--          Tolerance is used because we can't create a line 
	--          when the distance between the two points is too small.

Create (Qualified1 : QualifiedCirc from GccEnt  ;
        ThePoint   : Pnt2d         from gp      ;
        Tolerance  : Real          from Standard) returns Lin2d2Tan
raises BadQualifier;
	---Purpose: This methods implements the algorithms used to 
	--          create 2d lines tangent to one circle and passing
	--          thrue a point.
	--          Exception BadQualifier is raised in the case of 
	--          EnclosedCirc
      	--          Tolerance is used because there is no solution 
      	--          when the point is inside the solution according to 
      	--          the tolerance.

Create (Qualified1 : QualifiedCirc from GccEnt  ;
        Qualified2 : QualifiedCirc from GccEnt  ;
        Tolerance  : Real          from Standard) returns Lin2d2Tan
raises BadQualifier;
	---Purpose: This methods implements the algorithms used to 
	--          create 2d lines tangent to 2 circles.
	--          Exception BadQualifier is raised in the case of 
	--          EnclosedCirc

--------------------------------------------------------------------------

IsDone (me) returns Boolean from Standard
is static;
    	---Purpose: This method returns true when there is a solution 
    	--          and false in the other cases.

NbSolutions(me) returns Integer from Standard
    	---Purpose: This method returns the number of solutions.
    	--          Raises NotDone if the construction algorithm didn't succeed. 
raises NotDone
is static;
  

ThisSolution(me                           ; 
    	     Index : Integer from Standard) returns Lin2d 
    	---Purpose : Returns the solution number Index and raises OutOfRange 
    	--           exception if Index is greater than the number of solutions.
    	--           Be carefull: the Index is only a way to get all the 
    	--           solutions, but is not associated to theses outside the 
    	--           context of the algorithm-object. Raises OutOfRange is raised if Index is greater than 
    	--           the number of solutions.
    	--           It raises NotDone if the algorithm failed.
raises OutOfRange, NotDone
is static;
  

WhichQualifier(me                                  ;
    	       Index   :     Integer  from Standard;
	       Qualif1 : out Position from GccEnt  ;
	       Qualif2 : out Position from GccEnt  )
raises OutOfRange, NotDone
is static;
    	---Purpose: Returns the qualifiers Qualif1 and Qualif2 of the
    	-- tangency arguments for the solution of index Index
    	-- computed by this algorithm.
    	-- The returned qualifiers are:
    	-- -   those specified at the start of construction when the
    	--   solutions are defined as enclosing or outside with
    	--   respect to the arguments, or
    	-- -   those computed during construction (i.e. enclosing or
    	--   outside) when the solutions are defined as unqualified
    	--   with respect to the arguments, or
    	-- -   GccEnt_noqualifier if the tangency argument is a point.
    	--  Exceptions
    	-- Standard_OutOfRange if Index is less than zero or
    	-- greater than the number of solutions computed by this algorithm.
    	-- StdFail_NotDone if the construction fails.


Tangency1(me                                     ;
          Index         : Integer   from Standard;
          ParSol,ParArg : out Real  from Standard;
          PntSol        : out Pnt2d from gp      )
    	---Purpose : Returns informations about the tangency point between the 
    	--           result number Index and the first argument.
    	--           ParSol is the intrinsic parameter of the point PntSol on
    	--           the solution curv.
    	--           ParArg is the intrinsic parameter of the point PntSol on 
    	--           the argument curv. Raises OutOfRange is raised if Index is greater than 
    	--           the number of solutions.
    	--           It raises NotDone if the algorithm failed.
raises OutOfRange, NotDone
is static;
  
Tangency2(me                                     ;
          Index         : Integer   from Standard;
          ParSol,ParArg : out Real  from Standard;
          PntSol        : out Pnt2d from gp      )
    	---Purpose : Returns informations about the tangency point between the 
   	--           result number Index and the second argument.
    	--           ParSol is the intrinsic parameter of the point ParSol on
    	--           the solution curv.
    	--           ParArg is the intrinsic parameter of the point PntSol on 
    	--           the argument curv. Raises OutOfRange is raised if Index is greater than 
    	--          the number of solutions.
    	--          It raises NotDone if the algorithm failed.
raises OutOfRange, NotDone
is static;
  

fields

    WellDone : Boolean from Standard;
    	---Purpose : True if the algorithm succeeded.

    NbrSol   : Integer from Standard;
    	---Purpose : The number of possible solutions. We have to decide about the
    	--           status of the multiple solutions...

    linsol   : Array1OfLin2d from TColgp;
    	---Purpose : Thesolutions.

    qualifier1 : Array1OfPosition from GccEnt;
    	---Purpose: The qualifiers of the first argument.

    qualifier2 : Array1OfPosition from GccEnt;
   	---Purpose: The qualifiers of the second argument.

    pnttg1sol   : Array1OfPnt2d from TColgp;
    	---Purpose: The tangency point between the solution and the first 
    	--          argument on the solution.

    pnttg2sol   : Array1OfPnt2d from TColgp;
    	---Purpose: The tangency point between the solution and the second 
    	--          argument on the solution.

    par1sol   : Array1OfReal from TColStd;
    	---Purpose: The parameter of the tangency point between the solution 
    	--          and the first argument on the solution.

    par2sol   : Array1OfReal from TColStd;
    	---Purpose: The parameter of the tangency point between the solution 
    	--          and the second argument on the solution.

    pararg1   : Array1OfReal from TColStd;
    	---Purpose: The parameter of the tangency point between the solution 
    	--          and the first argument on the first argument.

    pararg2   : Array1OfReal from TColStd;
    	---Purpose: The parameter of the tangency point between the solution 
    	--          and the second argument on the second argument.

end Lin2d2Tan;
