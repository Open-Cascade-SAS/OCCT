-- Created on: 1993-03-09
-- Created by: Jean-Louis Frenkel
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class HLRToolShape from StdPrs

uses 
    Shape          from TopoDS,
    Curve          from BRepAdaptor,
    Data           from HLRBRep,
    EdgeIterator   from HLRAlgo,
    Projector      from HLRAlgo

is
    Create (TheShape    : Shape     from TopoDS;
            TheProjector: Projector from HLRAlgo) 
    	    returns HLRToolShape from StdPrs;
    NbEdges(me) returns Integer from Standard;
    InitVisible(me: in out; EdgeNumber: Integer from Standard);
    MoreVisible(me) returns Boolean from Standard;
    NextVisible(me: in out);
    Visible(me: in out ; TheEdge : out Curve from BRepAdaptor;
                U1,U2   : out Real from Standard);
    InitHidden(me:in out; EdgeNumber: Integer from Standard);
    MoreHidden(me) returns Boolean from Standard;
    NextHidden(me: in out);
    Hidden(me: in out; TheEdge : out Curve from BRepAdaptor; 
                U1,U2  : out Real from Standard);

fields
    MyData              : Data         from HLRBRep;
    myEdgeIterator      : EdgeIterator from HLRAlgo;
    MyCurrentEdgeNumber : Integer      from Standard;

end HLRToolShape from StdPrs;
