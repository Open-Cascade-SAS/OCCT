-- Created on: 1997-09-11
-- Created by: Roman BORISOV
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class ApproxCurve from Geom2dConvert 
    	---Purpose: A framework to convert a 2D curve to a BSpline.
    	--  This is done by approximation within a given tolerance.
	
uses 
    Curve          from  Geom2d, 
    BSplineCurve   from  Geom2d, 
    Shape          from  GeomAbs,
    OutOfRange     from  Standard          
    
raises  OutOfRange   from Standard

is
 
    Create  (Curve:  Curve  from  Geom2d; 
    	    Tol2d:  Real; 
    	    Order:  Shape  from  GeomAbs; 
    	    MaxSegments:  Integer; 
    	    MaxDegree:  Integer)  returns  ApproxCurve  from  Geom2dConvert; 
        ---Purpose: Constructs an approximation framework defined by
    	-- -   the 2D conic Curve
    	-- -   the tolerance value Tol2d
    	-- -   the degree of continuity Order
    	-- -   the maximum number of segments allowed MaxSegments
    	-- -   the highest degree MaxDegree which the
    	--   polynomial defining the BSpline is allowed to have.
     
    Curve(me)  returns  BSplineCurve  from  Geom2d; 
    	---Purpose: Returns the 2D BSpline curve resulting from the
    	--  approximation algorithm.
        
    IsDone(me)  returns  Boolean  from  Standard; 
    	---Purpose:  returns  Standard_True  if  the  approximation  has   
    	-- been  done  with  within  requiered tolerance  
     
    HasResult(me) returns Boolean; 
    	---Purpose: returns  Standard_True if the approximation did come out 
    	-- with a result that  is not NECESSARELY within the required tolerance 
    
    MaxError(me)  returns  Real  from  Standard; 
    	---Purpose: Returns the greatest distance between a point on the
    	-- source conic and the BSpline curve resulting from the
    	-- approximation. (>0 when an approximation 
    	--  has  been  done, 0  if  no  approximation) 
     
    Dump(me;  o:  in  out  OStream); 
    	---Purpose:  Print on the stream  o  information about the object

fields
    myCurve     : Curve           from  Geom2d;
    myIsDone    : Boolean         from  Standard; 
    myHasResult : Boolean         from  Standard; 
    myBSplCurve : BSplineCurve    from  Geom2d; 
    myMaxError  : Real            from  Standard; 
    
end ApproxCurve;
