-- Created on: 2001-05-25
-- Created by: Peter KURNEV
-- Copyright (c) 2001-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class SolidSolid from BOP inherits ShellSolid from BOP

	---Purpose:  
    	---        Performs Boolean Operations  (BO)  
    	---        Common,Cut,Fuse for solids as      
	---        arguments 
	---
uses 
    DSFiller     from BOPTools, 
     
    WireEdgeSet  from BOP,   
    ShellFaceSet from BOP, 

    HistoryCollector from BOP,
    IndexedDataMapOfIntegerIndexedMapOfInteger from BOPTColStd,
    DataMapOfShapeInteger from TopTools,
    Shape        from TopoDS,
    Solid        from TopoDS,
    State        from TopAbs,
    
    ListOfShape  from TopTools
    
    
is 
    Create   
    	returns SolidSolid from BOP; 
    	---Purpose:  
    	--- Empty constructor;
    	---
    DoWithFiller      (me:out; 
    	     aDSF: DSFiller from BOPTools) 
    	is  redefined; 
    	---Purpose:  
    	--- See base classes, please 
    	---
    Destroy (me: in out) 
    	is redefined; 
    	---C++: alias "Standard_EXPORT virtual ~BOP_SolidSolid(){Destroy();}"  
    	---Purpose:   
    	--- Destructor 
    	---
    DoNewFaces(me: out)    
    	is redefined;  
    	---Purpose:  
    	--- See base classes, please 
    	---
    BuildResult (me: out)
    	is  redefined; 
     	---Purpose:  
    	--- See base classes, please 
    	---

    SetHistoryCollector(me: in out; theHistory: HistoryCollector from BOP)
    	is redefined virtual;

    --- 
    ---              P  r  i  v  a  t  e    b  l  o  c  k   
    ---	     
    PrepareSFS  (me:out; 
    	    aFaces: ListOfShape from TopTools; 
	    aSFS  : out ShellFaceSet from BOP) 
	is  private;	     

    PrepareFaceSplits(me: out)
    	is private;

    PropagateFaceStateByEdges(me: in out; theFace:           Shape from TopoDS;
    	    	    	    	    	  theMapOfEdgeIndex: DataMapOfShapeInteger from TopTools;
    	    	    	    	    	  theState:          out State from TopAbs)
    	returns Boolean from Standard
    	is private;
	
    ComputeStateByInsidePoints(me: in out; theFaceIndex: Integer from Standard;
    	    	    	    	    	   theBaseFaceIndex: Integer from Standard;
    	    	    	    	    	   theFaceRank:  Integer from Standard;
					   theFFMap:     IndexedDataMapOfIntegerIndexedMapOfInteger from BOPTColStd;
    	    	    	    	    	   theState:     out State from TopAbs)
    	returns Boolean from Standard
    	is private;

    TakeOnSplit(me; theFaceIndex: Integer from Standard;
    	    	    theBaseFaceIndex: Integer from Standard)
    	returns Boolean from Standard
    	is private;
     
    PrepareReferences(me:out) 
    	is protected; 
    
fields  
    myRefObject: Solid from TopoDS is protected;   
    myRefTool  : Solid from TopoDS is protected;     
    
end SolidSolid;
