-- Created on: 1996-12-25
-- Created by: Alexander BRIVIN
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Cube from Vrml 

	---Purpose: defines a Cube node of VRML specifying geometry shapes.
    	-- This  node  represents  a  cuboid aligned with  the coordinate  axes. 
        -- By  default ,  the  cube  is  centred  at  (0,0,0) and  measures  2  units
	-- in  each  dimension, from -1  to  +1. 
    	-- A cube's width is its extent along its object-space X axis, its height is  
    	-- its extent along the object-space Y axis, and its depth is its extent along its
	-- object-space Z axis. 
is

    Create ( aWidth  : Real from Standard = 2;
    	     aHeight : Real from Standard = 2;
	     aDepth  : Real from Standard = 2 )
        returns Cube from Vrml;
    
    SetWidth ( me : in out; aWidth : Real from Standard );
    Width ( me  )  returns Real  from  Standard;
    
    SetHeight ( me : in out; aHeight : Real from Standard );
    Height ( me  )  returns Real  from  Standard;
    
    SetDepth ( me : in out; aDepth : Real from Standard );
    Depth ( me )  returns Real  from  Standard;

    Print  ( me;  anOStream: in out OStream from Standard) returns OStream from Standard;
    ---C++:  return  & 

fields

    myWidth  : Real from Standard;  -- Size in x dimension
    myHeight : Real from Standard;  -- Size in y dimension
    myDepth  : Real from Standard;  -- Size in z dimension

end Cube;

