-- Created on: 1994-07-19
-- Created by: Guest Kernel
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Convert from Quantity

    	---Purpose: Services to manage units conversion between Front-ends and Engines.
    	-- This conversion is managed by a table of correspondance between the quantities
    	-- and their "conversion coefficient".
    	-- This table is implemented like an external array (TCollection_Array1) regarding 
    	-- to the quantities enumeration.
     
uses 
    AsciiString from TCollection,
    PhysicalQuantity from Quantity,
    Coefficient from Quantity
	     
is

    Create returns Convert from Quantity;
    	---Purpose: Creates an object;

    SetQuantity(myclass ; 
                aQuantity : PhysicalQuantity from Quantity ;
	        aCoef: Coefficient from Quantity);	    
    	---Purpose: Updates the conversion table (correspondances between 
    	-- Quantities and conversion coefficients).
    	---C++: inline

    ConvertUserToSI(myclass ; 
                    aQuantity : PhysicalQuantity from Quantity ;
          	    aVal : Real from Standard)
    returns Real from Standard;
        ---Purpose: Converts, from the conversion table, the value <aVal>
    	-- from the user system to the SI system. 
    	---C++: inline

    ConvertSIToUser(myclass ; 
                    aQuantity : PhysicalQuantity from Quantity ;
          	    aVal : Real from Standard)
    returns Real from Standard;
    	---Purpose: Converts, from the conversion table, the value <aVal>
   	-- from the SI system to the user system. 
    	---C++: inline

    IsPhysicalQuantity(myclass; 
                       aTypeName : AsciiString from TCollection ; 
                       anEnum : in out AsciiString from TCollection)
    returns Boolean from Standard;
    	---Purpose:
    	-- if (aType is a physical quantity)
    	--    returns True and the name of the associated PhysicalQuantity .
    	-- else 
    	--    returns False.

end Convert from Quantity;
	        	







































































































