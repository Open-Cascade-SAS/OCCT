-- Created on: 1999-09-24
-- Created by: Sergey ZARITCHNY
-- Copyright (c) 1999-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package QANewBRepNaming 

	---Purpose: Implements  methods   to   load  the  Make   Shape
	--          operations in  the  naming data-structure (package
	--          TNaming),  which    provides  topological   naming
	--          facilities.  Shape  generation, modifications  and
	--          deletions   are  recorded in   the  data-framework
	--          (package  TDF)   using the builder  from   package
	--          TNaming.

uses 
 
    TDF,
    TNaming,
    TopAbs,
    TopLoc,
    TopTools,
    TopoDS, 
--    FeatAlgo, 
    BRepAlgo,
    BRepAlgoAPI,
    BRepPrimAPI, 
    BRepBuilderAPI, 
    BRepOffsetAPI, 
    BRepFilletAPI,
    QANewModTopOpe
    
is

    ---Level: Public

    enumeration TypeOfPrimitive3D is
	SHELL,
	SOLID
    end TypeOfPrimitive3D;

    class LoaderParent;

    class Loader;

    deferred class TopNaming;

    	---Level: Primitives

    	class Box;
    
    	class Prism; 
     
    	class Revol; 

    	--class Cone;

    	class Cylinder;

    	class Sphere; 
	 
	--class Torus; 
	 
	--class Pipe;

	--class PipeShell;

	--class CircularPipe;


    	---Level: Boolean operation (Cut, Fuse, Common)

    	class BooleanOperation;      -- creation of a new part (primitive)

    	deferred class BooleanOperationFeat;  -- modification one of the shapes (feature)
	
    	    class Common;

    	    class Cut;

    	    class Fuse;

    	    --class Section;


    	---Level: Fillet & Chamfer

    	class Fillet;

    	class Chamfer;

    
    	---Level: Importation

    	class ImportShape;

    	class Gluing;
	
	class Intersection;
	
	class Limitation;


    	---Level: Offset

        --class Draft;		  
 
    	--class ThickSolid; 
	 
	--class ThruSections; 
	 
	--class Vary;


    	---Level: Features

	--class DPrism; 
	 
    	--class Hole;

    	--class LinearForm; 
	 
	--class Mirror; 
	 
	--class PipeFeat;

    	--class Scale;

    	--class PrismFeat; 
	 
	--class RevolFeat;

    	CleanStructure (theLabel : Label from TDF);

    	LoadNamedShape (theBuilder : in out Builder from TNaming;
			theEvol : Evolution from TNaming;
			theOS : Shape from TopoDS;
			theNS : Shape from TopoDS);

    	Displace (theLabel : Label from TDF;
                  theLoc : Location from TopLoc;
                  theWithOld : Boolean from Standard);

end QANewBRepNaming;
