-- Created on: 1999-03-05
-- Created by: Fabrice SERVANT
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Edge from IntPolyh

uses
    
    Pnt from gp


is


    Create;
    
    Create(i1,i2,i3,i4: Integer from Standard) ; 
    
    FirstPoint(me) 
    returns Integer from Standard
    is static;

    SecondPoint(me) 
    returns Integer from Standard
    is static;
    
    FirstTriangle(me) 
    returns Integer from Standard
    is static;

    SecondTriangle(me) 
    returns Integer from Standard
    is static;
    
    AnalysisFlag(me) 
    returns Integer from Standard
    is static;
    
--    GetTriangles(me; T1,T2: Integer from Standard)
--    is static;

    SetFirstPoint(me: in out; v: Integer from Standard) 
    is static;
	
    SetSecondPoint(me: in out; v: Integer from Standard) 
    is static;
    
    SetFirstTriangle(me: in out; v: Integer from Standard) 
    is static;
	
    SetSecondTriangle(me: in out; v: Integer from Standard) 
    is static;
    
    SetAnalysisFlag(me: in out; v: Integer from Standard) 
    is static;
    
--    SetTriangles(me: in out; T1,T2: in out Integer from Standard) 
--    is static;
    
    Dump(me; v: Integer from Standard) 
    is static;
     	
fields

    p1,p2 : Integer from Standard;
    t1,t2 : Integer from Standard;
    ia    : Integer from Standard;
    
end Edge from IntPolyh;
