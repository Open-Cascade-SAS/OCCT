-- Created on: 2002-01-25
-- Created by: doneux <doneux@samcef.com>
-- Copyright (c) 2002-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Real2String from OSD 

	---Purpose:  Convertion of CString to Real and reciprocally

is 

    Create
    	returns Real2String from OSD;
 
    RealToCString(me;
    	    	  aReal: Real;
    	    	  aString:out PCharacter) 
     returns Boolean ;
    ---Purpose:
    --  Converts aReal into aCstring in exponential format with maximum
    --  17 digits. The size of the destination string must be sufficient (at least 23 characters)
    --  The decimal separator account for locale setting, but 
    --  neither thousand separator nor grouping of digits in the output string.
    --  

    CStringToReal(me: in out;
    	          aString: CString; 
    	    	  aReal: out Real) returns Boolean ;
    ---Purpose:
    --  Converts aCstring representing a real. The first occurence of the decimal separator
    --  (comma or period) defines it values for further readings.
   --  Neither thousand separator nor grouping of digits are allowed in the CString

fields

    myReadDecimalPoint: Integer from Standard;
    myLocalDecimalPoint: Integer from Standard;

end Real2String;
