-- Created on: 2000-02-14
-- Created by: Denis PASCAL
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class CopyShape from TNaming 

	---Purpose: 

uses Shape from TopoDS,
     IndexedDataMapOfTransientTransient from TColStd,
     TranslateTool from TNaming,
     Location from TopLoc

is

    CopyTool (myclass;
              aShape    :  Shape      from TopoDS;
    	      aMap      :  in out  IndexedDataMapOfTransientTransient from TColStd; 
	      aResult   :  in  out Shape  from  TopoDS);
	---Purpose:      Makes  copy  a  set  of  shape(s),  using the  aMap 
	 
	  
    Translate (myclass;
               aShape  : Shape          from TopoDS; 
	       aMap    : in out  IndexedDataMapOfTransientTransient from TColStd; 
	       aResult : in  out Shape  from  TopoDS;
    	       TrTool  : TranslateTool  from TNaming); 
	     
	 ---Purpose: Translates  a  Transient  shape(s)  to  Transient     
	    
    Translate (myclass;
               L : Location from TopLoc; 
     	       aMap :  in out  IndexedDataMapOfTransientTransient from TColStd)   	       
    returns Location from TopLoc; 
     ---Purpose: Translates a Topological  Location  to an  other  Top.
     --          Location 

end CopyShape;
