-- Created on: 2004-06-22
-- Created by: STV
-- Copyright (c) 2004-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class ColorScale from Aspect inherits TShared from MMgt
        ---Purpose: Defines a color scale for viewer.
uses

       TypeOfColorScaleData     from Aspect,
       TypeOfColorScalePosition from Aspect,
       SequenceOfColor          from Aspect,
       Color                    from Quantity,
       AsciiString              from TCollection,
       ExtendedString           from TCollection,
       SequenceOfExtendedString from TColStd

is

	---Category: Public

       FindColor( me; theValue : Real from Standard;
                      theColor : in out Color from Quantity ) returns Boolean from Standard;
       ---Purpose: Calculate color according passed value; returns true if value is in range or false, if isn't


       FindColor( myclass; theValue : Real from Standard;
                           theMin, theMax : Real from Standard;
                           theColorsCount : Integer from Standard;
                           theColor : in out Color from Quantity ) returns Boolean from Standard;

       GetMin(me)
       returns Real from Standard;
       ---Purpose: Returns minimal value of color scale;

       GetMax(me)
       returns Real from Standard;
       ---Purpose: Returns maximal value of color scale;

       GetRange(me; theMin : in out Real from Standard;
                    theMax : in out Real from Standard);
       ---Purpose: Returns minimal and maximal values of color scale;

       GetLabelType(me)
       returns TypeOfColorScaleData from Aspect;
       ---Purpose: Returns the type of labels;
       ---         Aspect_TOCSD_AUTO - labels as boundary values for intervals
       ---         Aspect_TOCSD_USER - user specified label is used

	GetColorType(me)
       returns TypeOfColorScaleData from Aspect;
       ---Purpose: Returns the type of colors;
       ---         Aspect_TOCSD_AUTO - value between Red and Blue
       ---         Aspect_TOCSD_USER - user specified color from color map

       GetNumberOfIntervals(me)
       returns Integer from Standard;
       ---Purpose: Returns the number of color scale intervals;

       GetTitle(me)
       returns ExtendedString from TCollection;
       ---Purpose: Returns the color scale title string;

       GetFormat(me)
       returns AsciiString from TCollection;
       ---Purpose: Returns the format for numbers.
       --         The same like format for function printf().
       --         Used if GetLabelType() is TOCSD_AUTO;

	GetLabel(me; theIndex : Integer from Standard)
       returns ExtendedString from TCollection;
       ---Purpose: Returns the user specified label with index <anIndex>.
       --         Returns empty string if label not defined.

	GetColor(me; theIndex : Integer from Standard)
       returns Color from Quantity;
       ---Purpose: Returns the user specified color from color map with index <anIndex>.
       --         Returns default color if index out of range in color map.

       GetLabels(me; theLabels : in out SequenceOfExtendedString from TColStd);
       ---Purpose: Returns the user specified labels.

       GetColors(me; theColors : in out SequenceOfColor from Aspect);
       ---Purpose: Returns the user specified colors.

       GetLabelPosition(me)
       returns TypeOfColorScalePosition from Aspect;
       ---Purpose: Returns the position of labels concerning color filled rectangles.

	GetTitlePosition(me)
       returns TypeOfColorScalePosition from Aspect;
       ---Purpose: Returns the position of color scale title.

	IsReversed(me)
       returns Boolean from Standard;
	---Purpose: Returns true if the labels and colors used in reversed order.

	IsLabelAtBorder(me)
       returns Boolean from Standard;
	---Purpose: Returns true if the labels placed at border of color filled rectangles.

       SetMin(me : mutable; theMin : Real from Standard);
       ---Purpose: Sets the minimal value of color scale.

       SetMax(me : mutable; theMax : Real from Standard);
       ---Purpose: Sets the maximal value of color scale.

       SetRange(me : mutable; theMin : Real from Standard;
                              theMax : Real from Standard);
       ---Purpose: Sets the minimal and maximal value of color scale.

       SetLabelType(me : mutable; theType : TypeOfColorScaleData from Aspect);
       ---Purpose: Sets the type of labels.
       --         Aspect_TOCSD_AUTO - labels as boundary values for intervals
       --         Aspect_TOCSD_USER - user specified label is used

       SetColorType(me : mutable; theType : TypeOfColorScaleData from Aspect);
       ---Purpose: Sets the type of colors.
       --         Aspect_TOCSD_AUTO - value between Red and Blue
       --         Aspect_TOCSD_USER - user specified color from color map

       SetNumberOfIntervals(me : mutable; theNum : Integer from Standard);
       ---Purpose: Sets the number of color scale intervals.

       SetTitle(me : mutable; theTitle : ExtendedString from TCollection);
       ---Purpose: Sets the color scale title string.

       SetFormat(me : mutable; theFormat : AsciiString from TCollection);
       ---Purpose: Sets the color scale auto label format specification.

       SetLabel(me : mutable; theLabel  : ExtendedString from TCollection;
                              anIndex : Integer from Standard = -1);
       ---Purpose: Sets the color scale label at index. Index started from 1.

       SetColor(me : mutable; theColor  : Color from Quantity;
                              theIndex : Integer from Standard = -1);
       ---Purpose: Sets the color scale color at index. Index started from 1.

       SetLabels(me : mutable; theSeq : SequenceOfExtendedString from TColStd);
       ---Purpose: Sets the color scale labels.

       SetColors(me : mutable; theSeq : SequenceOfColor from Aspect);
       ---Purpose: Sets the color scale colors.

       SetLabelPosition(me : mutable; thePos : TypeOfColorScalePosition from Aspect);
       ---Purpose: Sets the color scale labels position concerning color filled rectangles.

       SetTitlePosition(me : mutable; thePos : TypeOfColorScalePosition from Aspect);
       ---Purpose: Sets the color scale title position.

	SetReversed(me : mutable; theReverse : Boolean from Standard);
	---Purpose: Sets true if the labels and colors used in reversed order.

	SetLabelAtBorder(me : mutable; theOn : Boolean from Standard);
	---Purpose: Sets true if the labels placed at border of color filled rectangles.

       --- Size and position management
       --- Size and position are values relative to view size (between 0 and 1)

       GetSize(me; theWidth  : in out Real from Standard;
                   theHeight : in out Real from Standard);
	---Purpose: Returns the size of color scale.

       GetWidth(me)
       returns Real from Standard;
	---Purpose: Returns the width of color scale.

       GetHeight(me)
       returns Real from Standard;
	---Purpose: Returns the height of color scale.

       SetSize(me : mutable; theWidth  : Real from Standard;
                             theHeight : Real from Standard);
	---Purpose: Sets the size of color scale.

       SetWidth(me : mutable; theWidth : Real from Standard);
	---Purpose: Sets the width of color scale.

       SetHeight(me : mutable; theHeight : Real from Standard);
	---Purpose: Sets the height of color scale.

       GetPosition(me; theX : in out Real from Standard;
                       theY : in out Real from Standard);
	---Purpose: Returns the position of color scale.

       GetXPosition(me)
       returns Real from Standard;
	---Purpose: Returns the X position of color scale.

       GetYPosition(me)
       returns Real from Standard;
	---Purpose: Returns the height of color scale.

       SetPosition(me : mutable; theX : Real from Standard;
                                 theY : Real from Standard);
	---Purpose: Sets the position of color scale.

       SetXPosition(me : mutable; theX : Real from Standard);
	---Purpose: Sets the X position of color scale.

       SetYPosition(me : mutable; theY : Real from Standard);
	---Purpose: Sets the Y position of color scale.

	GetTextHeight(me)
	returns Integer from Standard;
 ---Purpose: Returns the height of text of color scale.

	SetTextHeight(me: mutable; theHeight :  Integer from Standard);
 ---Purpose: Sets the height of text of color scale.

	---Category: Protected


	Initialize
       returns ColorScale from Aspect
       is protected;
	---Purpose: Default constructor.

       SizeHint(me; theWidth  : in out Integer from Standard;
                    theHeight : in out Integer from Standard)
       is protected;
	---Purpose: Returns the size of color scale.
    -- @param theWidth [out] the width of color scale.
    -- @param theHeight [out] the height of color scale.


       UpdateColorScale(me : mutable)
       is virtual protected;
	---Purpose: updates color scale parameters.

       DrawScale(me : mutable; theBgColor : Color from Quantity;
                      theX, theY, theWidth, theHeight : Integer from Standard)
       is protected;
	---Purpose: Draws color scale.
    -- @param theBgColor [in] background color
    -- @param theX [in] the X coordinate of color scale position.
    -- @param theY [in] the Y coordinate of color scale position.
    -- @param theWidth [in] the width of color scale.
    -- @param theHeight [in] the height of color scale.

	BeginPaint(me : mutable)
       returns Boolean from Standard
       is virtual protected;

	EndPaint(me : mutable)
       returns Boolean from Standard
       is virtual protected;

       PaintRect(me : mutable; theX, theY, theWidth, theHeight : Integer from Standard;
                               theColor     : Color from Quantity;
                               theFilled    : Boolean from Standard = Standard_False)
       is deferred;
    ---Purpose: Draws a rectangle.
    -- @param theX [in] the X coordinate of rectangle position.
    -- @param theY [in] the Y coordinate of rectangle position.
    -- @param theWidth [in] the width of rectangle.
    -- @param theHeight [in] the height of rectangle.
    -- @param theColor [in] the color of rectangle.
    -- @param theFilled [in] defines if rectangle must be filled.

	PaintText(me : mutable; theText : ExtendedString from TCollection;
                               theX, theY : Integer from Standard;
                               theColor : Color from Quantity)
       is deferred;
    ---Purpose: Draws a text.
    -- @param theText [in] the text to draw.
    -- @param theX [in] the X coordinate of text position.
    -- @param theY [in] the Y coordinate of text position.
    -- @param theColor [in] the color of text.

	TextWidth(me; theText : ExtendedString from TCollection)
       returns Integer from Standard
       is deferred;
    ---Purpose: Returns the width of text.
    -- @param theText [in] the text of which to calculate width.

	TextHeight(me; theText : ExtendedString from TCollection)
       returns Integer from Standard
       is deferred;
    ---Purpose: Returns the height of text.
    -- @param theText [in] the text of which to calculate height.

	---Category: Private

       Format(me)
       returns AsciiString from TCollection
       is private;
    ---Purpose: Returns the format of text.

       GetNumber(me; theIndex : Integer from Standard)
       returns Real from Standard
       is private;
    ---Purpose: Returns the value of given interval.

       HueFromValue(myclass; theValue : Integer from Standard;
                             theMin   : Integer from Standard;
                             theMax   : Integer from Standard)
       returns Integer from Standard
       is private;
    ---Purpose: Returns the color's hue for the given value in the given interval.
    -- @param theValue [in] the current value of interval.
    -- @param theMin [in] the min value of interval.
    -- @param theMax [in] the max value of interval.

fields

       myMin, myMax            : Real from Standard;
       myTitle                 : ExtendedString from TCollection;
       myFormat                : AsciiString from TCollection;
       myInterval              : Integer from Standard;
       myColorType             : TypeOfColorScaleData from Aspect;
       myLabelType             : TypeOfColorScaleData from Aspect;

       myAtBorder              : Boolean from Standard;
       myReversed              : Boolean from Standard;

       myColors                : SequenceOfColor          from Aspect;
       myLabels                : SequenceOfExtendedString from TColStd;

       myLabelPos              : TypeOfColorScalePosition from Aspect;
       myTitlePos              : TypeOfColorScalePosition from Aspect;

       myXPos,  myYPos         : Real from Standard;
       myWidth, myHeight       : Real from Standard;

       myTextHeight            : Integer from Standard;

end ColorScale;
