-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class DimensionalExponents from StepBasic 

inherits TShared from MMgt

uses

	Real from Standard
is

	Create returns mutable DimensionalExponents;
	---Purpose: Returns a DimensionalExponents

	Init (me : mutable;
	      aLengthExponent : Real from Standard;
	      aMassExponent : Real from Standard;
	      aTimeExponent : Real from Standard;
	      aElectricCurrentExponent : Real from Standard;
	      aThermodynamicTemperatureExponent : Real from Standard;
	      aAmountOfSubstanceExponent : Real from Standard;
	      aLuminousIntensityExponent : Real from Standard) is virtual;

	-- Specific Methods for Field Data Access --

	SetLengthExponent(me : mutable; aLengthExponent : Real);
	LengthExponent (me) returns Real;
	SetMassExponent(me : mutable; aMassExponent : Real);
	MassExponent (me) returns Real;
	SetTimeExponent(me : mutable; aTimeExponent : Real);
	TimeExponent (me) returns Real;
	SetElectricCurrentExponent(me : mutable; aElectricCurrentExponent : Real);
	ElectricCurrentExponent (me) returns Real;
	SetThermodynamicTemperatureExponent(me : mutable; aThermodynamicTemperatureExponent : Real);
	ThermodynamicTemperatureExponent (me) returns Real;
	SetAmountOfSubstanceExponent(me : mutable; aAmountOfSubstanceExponent : Real);
	AmountOfSubstanceExponent (me) returns Real;
	SetLuminousIntensityExponent(me : mutable; aLuminousIntensityExponent : Real);
	LuminousIntensityExponent (me) returns Real;

fields

	lengthExponent : Real from Standard;
	massExponent : Real from Standard;
	timeExponent : Real from Standard;
	electricCurrentExponent : Real from Standard;
	thermodynamicTemperatureExponent : Real from Standard;
	amountOfSubstanceExponent : Real from Standard;
	luminousIntensityExponent : Real from Standard;

end DimensionalExponents;
