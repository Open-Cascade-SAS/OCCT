-- Created on: 1993-03-23
-- Created by: BBL,JLF
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class XPR from ImageUtility

	---Version: 0.0

	---Purpose: Performs a "xpr" with a XAlienImage build
	-- 		 from any Image , any AlienImage .

	---Keywords:
	---Warning:
	---References:

uses
	AlienUserImage 	from AlienImage,
	XAlienImage  	from AlienImage,
	File  		from OSD,
	Image 		from Image

raises
	TypeMismatch 	from Standard

is
	XPR ( myclass ; aImage          : in Image from Image; 
			aName           : CString from Standard;
			xprOptions      : CString from Standard 
						= "" ) ;
	---Level: Internal
	  ---Purpose: Write content of a Image object to aTmpFile and
	  --          execute a Spawn "xpr xprOptions aTmpFile | lpr &" .

	XPR ( myclass ; aAlienUserImage : in AlienUserImage from AlienImage; 
			aName           : CString from Standard ;
			xprOptions      : CString from Standard 
						= "" ) ;
	---Level: Internal
	  ---Purpose: Write content of a  AlienImage object to aTmpFile and
	  --          execute a Spawn "xpr xprOptions aTmpFile| lpr  &" .

	XPR ( myclass ; aXAlienImage    : in XAlienImage from AlienImage ;
			xprOptions      : CString from Standard 
						= "" ) ;
	---Level: Internal
	  ---Purpose: Write content of a  XAlienImage object to aTmpFile and
	  --          execute a Spawn "xpr xprOptions aTmpFile| lpr  &" .

	XPR ( myclass ; aFile           : in File from OSD ;
			xprOptions      : CString from Standard 
						= "" ) ;
	---Level: Internal
	  ---Purpose: execute a Spawn 
	  --	"xpr xprOptions /aFile.SystemName()/ | lpr &" .

	XPR ( myclass ; aFileName       : CString from Standard ;
			xprOptions      : CString from Standard 
						= "" ) ;
	---Level: Internal
	  ---Purpose: execute a Spawn "xpr xprOptions aFileName | lpr &" .



end ;
