-- File:	StepShape_MeasureQualification.cdl
-- Created:	Tue Apr 24 13:58:11 2001
-- Author:	Christian CAILLET
--		<cky@photox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 2001

class MeasureQualification  from StepShape    inherits TShared

    ---Purpose : Added for Dimensional Tolerances

uses
    HAsciiString from TCollection,
    MeasureWithUnit from StepBasic,
    ValueQualifier from StepShape,
    HArray1OfValueQualifier from StepShape

is

    Create returns mutable MeasureQualification;

    Init (me : mutable; name : HAsciiString from TCollection;
    	    description : HAsciiString from TCollection;
	    qualified_measure : MeasureWithUnit from StepBasic;
	    qualifiers : HArray1OfValueQualifier from StepShape);

    Name (me) returns HAsciiString from TCollection;
    SetName (me : mutable; name : HAsciiString from TCollection);

    Description (me) returns HAsciiString from TCollection;
    SetDescription (me : mutable; description : HAsciiString from TCollection);

    QualifiedMeasure (me) returns MeasureWithUnit from StepBasic;
    SetQualifiedMeasure (me : mutable; qualified_measure : MeasureWithUnit from StepBasic);

    Qualifiers (me) returns HArray1OfValueQualifier from StepShape;
    NbQualifiers (me) returns Integer;
    SetQualifiers (me : mutable; qualifiers : HArray1OfValueQualifier from StepShape);
    QualifiersValue (me; num : Integer) returns ValueQualifier from StepShape;
    SetQualifiersValue (me : mutable; num : Integer; aqualifier : ValueQualifier from StepShape);

fields

    theName : HAsciiString from TCollection;
    theDescription : HAsciiString from TCollection;
    theQualifiedMeasure : MeasureWithUnit from StepBasic;
    theQualifiers : HArray1OfValueQualifier from StepShape;

end MeasureQualification;
