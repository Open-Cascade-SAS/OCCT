-- Created on: 2000-09-07
-- Created by: TURIN  Anatoliy <ati@nnov.matra-dtv.fr>
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Application from AppStd inherits Application from TDocStd

uses MessageDriver            from CDM,
     SequenceOfExtendedString from TColStd, 
     ExtendedString           from TCollection

is
   
    Create returns mutable Application from AppStd; 

    MessageDriver(me: mutable)
        returns MessageDriver from CDM
    is redefined;

    Formats(me: mutable; theFormats: out SequenceOfExtendedString from TColStd) 
    ---Purpose: returns supported format for application documents.
    is redefined;    

    ResourcesName (me: mutable)
    ---Purpose: returns   the file  name  which  contains  application
    --          resources
        returns CString from Standard;

fields
    myMessageDriver : MessageDriver from CDM;

end Application;
