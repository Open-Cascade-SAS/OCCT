-- File:	TopoDS_Face.cdl
-- Created:	Mon Dec 17 11:12:03 1990
-- Author:	Remi Lequette
---Copyright:	 Matra Datavision 1990, 1992


class Face from TopoDS inherits Shape from TopoDS

	---Purpose: Describes a face which
-- - references an underlying face with the potential to
--   be given a location and an orientation
-- - has a location for the underlying face, giving its
--   placement in the local coordinate system
-- - has an orientation for the underlying face, in terms
--   of its geometry (as opposed to orientation in relation to other shapes).

is
    Create returns Face from TopoDS;
    ---C++: inline
	---Purpose: Undefined Face.

end Face;
