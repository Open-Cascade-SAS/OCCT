-- Created on: 1995-03-10
-- Created by: Mister rmi
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Modified on july 97 by ROB : Field HArray instead Of ArrayOfPnt3D
--                      (connected entities)


class SensitiveCurve   from Select3D 
inherits SensitivePoly from Select3D

    ---Purpose: A framework to define a sensitive 3D curve.
    -- In some cases this class can raise Standard_ConstructionError and 
    -- Standard_OutOfRange exceptions. For more details see Select3D_SensitivePoly.

uses
    Pnt             from gp,
    Pnt2d           from gp,
    Projector       from Select3D,
    Lin             from gp,
    EntityOwner     from SelectBasics,
    ListOfBox2d     from SelectBasics,
    PickArgs        from SelectBasics,
    Curve           from Geom,
    Array1OfPnt     from TColgp,
    Array1OfPnt2d   from TColgp,
    HArray1OfPnt     from TColgp,
    Box2d           from Bnd,
    Location                 from TopLoc, 
    SensitiveEntity   from Select3D

raises
    ConstructionError from Standard,
    OutOfRange from Standard
is


    Create (OwnerId      : EntityOwner from SelectBasics;
            TheCurve     : Curve from Geom;
            MaxPoints    : Integer = 17)
     returns mutable SensitiveCurve;
        ---Level: Public 
        ---Purpose: Constructs a sensitive curve object defined by the
        -- owner OwnerId, the curve TheCurve, and the
        -- maximum number of points on the curve: MaxPoints.

    Create (OwnerId      : EntityOwner from SelectBasics;
            ThePoints    : HArray1OfPnt from TColgp)
     returns mutable SensitiveCurve;
        ---Level: Public 
        ---Purpose: Constructs a sensitive curve object defined by the
        -- owner OwnerId and the set of points ThePoints.
        
    Create (OwnerId      : EntityOwner from SelectBasics;
            ThePoints    : Array1OfPnt from TColgp)
     returns mutable SensitiveCurve;
        ---Level: Public 
        ---Purpose: Creation of Sensitive Curve from Points.
        --          Warning : This Method should disappear in the next version...

    Matches (me : mutable;
             thePickArgs : PickArgs from SelectBasics;
             theMatchDMin, theMatchDepth : out Real from Standard)
    returns Boolean is redefined static;
    ---Level: Public
    ---Purpose: Checks whether the sensitive entity matches the picking
    -- detection area (close to the picking line).
    -- For details please refer to base class declaration.

    Matches (me  :mutable; 
             XMin,YMin,XMax,YMax : Real from Standard;
             aTol: Real from Standard)
    returns Boolean
    is static;
     
    Matches (me  :mutable; 
             Polyline:Array1OfPnt2d from TColgp;
             aBox:Box2d from Bnd;
             aTol: Real from Standard) 
    returns Boolean
    is redefined virtual;
        ---Level: Public 
    

    ComputeDepth (me;
                  thePickLine : Lin from gp;
                  theDetectedIndex : Integer from Standard)
    returns Real from Standard;
    ---Level: Public
    ---Purpose: Compute depth of sensitive circle for the detected sub-part.
    -- @param thePickLine [in] the picking line.
    -- @param theDetectedIndex [in] index of the detected sub-part.
    -- @return depth on the picking line.
 
    GetLastDetected(me) returns Integer from Standard;
    ---Purpose: Gets index of last detected segment 
    ---C++: inline


        ---Category: Internal Methods
    Dump(me; S: in out OStream;FullDump : Boolean from Standard = Standard_True) is redefined virtual; 
     
    LoadPoints(me:mutable;aCurve:Curve from Geom;NbPoints: Integer) is static private; 

    GetConnected(me: mutable; theLocation : Location from TopLoc) 
    returns SensitiveEntity from Select3D 
    is redefined virtual; 
        ---Level: Public 
        ---Purpose: Returns the copy of this

fields
    mylastseg : Integer        from Standard;
    myCurve  : Curve from Geom;
end SensitiveCurve;

