-- Created on: 1997-05-06
-- Created by: Jean-Louis Frenkel, Remi Lequette
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package CDM


uses TCollection,TColStd,Resource

is

    enumeration CanCloseStatus is CCS_OK, CCS_NotOpen, CCS_UnstoredReferenced,CCS_ModifiedReferenced,CCS_ReferenceRejection
    end CanCloseStatus from CDM;


    class MetaData;

    deferred class MessageDriver;

    deferred class Document;

    class ReferenceIterator;
    
    class NullMessageDriver; 
    ---Purpose: a MessageDriver that writes nowhere.

    class COutMessageDriver;
    ---Purpose: aMessageDriver for output to COUT (only ASCII strings)

---Category: classes to manager automatic naming of documents.

    private alias NamesDirectory is DataMapOfStringInteger from TColStd;
    ---Purpose: this map will allows to get a directory object from a name.

    private class PresentationDirectory instantiates DataMap from TCollection 
    ---Purpose: this map will allows to get a directory object from a name.
        (ExtendedString from TCollection,
         Document from CDM,
         ExtendedString from TCollection);
         
    private pointer DocumentPointer to Document from CDM;
    private class Reference;    

    private class ListOfReferences instantiates List from TCollection(Reference from CDM);
    deferred class Application;
    
    private class MetaDataLookUpTable instantiates DataMap from TCollection(ExtendedString from TCollection, MetaData from CDM, ExtendedString from TCollection);
         
         
---Category: reusable classes

    class DocumentHasher instantiates MapHasher from TCollection(Document from CDM);
    class MapOfDocument instantiates Map from TCollection(Document from CDM, DocumentHasher from CDM);
    class ListOfDocument instantiates List from TCollection(Document from CDM);

end CDM;
