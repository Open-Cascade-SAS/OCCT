-- Created on: 1991-09-06
-- Created by: NW,JPB,CAL
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

--      27/09/97 ; PCT : add manual control of  textures
--              11/97 ; CAL : ajout polyline par 2 points
--      16/06/2000 : ATS: Study G005 - Group store presentations of it's objects in field
--                        MyListOfPArray to avoid deletion of handle-manipulating 
--                        primitives.
class Group from Graphic3d inherits TShared
    
        ---Version:

        ---Purpose: This class allows the definition of groups
        --     of primitives inside of graphic objects (presentations).
        --     A group contains the primitives and attributes
        --     for which the range is limited to this group.
        --     The primitives of a group can be globally suppressed.
        --
        --      There are two main group usage models:
        --
        --        1) Non-modifiable, or unbounded, group ('black box'). 
        --           Developers can repeat a sequence of 
        --           SetPrimitivesAspect() with AddPrimitiveArray() methods arbitrary number of times
        --           to define arbitrary number of primitive "blocks" each having individual apect values.
        --           Any modification of such a group is forbidden, as aspects and primitives are mixed 
        --           in memory without any high-level logical structure, and any modification is very likely to result
        --           in corruption of the group internal data.
        --           It is necessary to recreate such a group as a whole when some attribute should be changed.
        --           (for example, in terms of AIS it is necessary to re-Compute() the whole presentation each time).
        --        2) Bounded group. Developers should specify the necessary group aspects with help of
        --           SetGroupPrimitivesAspect() and then add primitives to the group.
        --           Such a group have simplified organization in memory (a single block of attributes
        --           followed by a block of primitives) and therefore it can be modified, if it is necessary to
        --           change parameters of some aspect that has already been set, using methods:
        --           IsGroupPrimitivesAspectSet() to detect which aspect was set for primitives;
        --           GroupPrimitivesAspect() to read current aspect values
        --           and SetGroupPrimitivesAspect() to set new values.
        -- 
        --        Developers are strongly recommended to take all the above into account when filling Graphic3d_Group
        --        with aspects and primitives and choose the group usage model beforehand out of application needs.

        ---Warning:
        ---References:
    
    uses
    
        Array1OfInteger             from TColStd,
        Array1OfReal                from TColStd,
        HArray1OfByte               from TColStd,
    
        ExtendedString              from TCollection,
    
        PlaneAngle                  from Quantity,
    
        Array1OfEdge                from Aspect,
        Edge                        from Aspect,
    
    	GroupAspect	            from Graphic3d,
        AspectLine3d                from Graphic3d,
        AspectMarker3d              from Graphic3d,
        AspectText3d                from Graphic3d,
        AspectFillArea3d            from Graphic3d,
        HorizontalTextAlignment     from Graphic3d,
        CBitFields4                 from Graphic3d,
        CGroup                      from Graphic3d,
        GraphicDriver               from Graphic3d,
        Structure                   from Graphic3d,
        TextPath                    from Graphic3d,
        Vector                      from Graphic3d,
        Array1OfVertex              from Graphic3d,
        Array2OfVertex              from Graphic3d,
        Vertex                      from Graphic3d,
        VerticalTextAlignment       from Graphic3d, 
        ArrayOfPrimitives           from Graphic3d,
        ListOfPArray                from Graphic3d,
        TransModeFlags              from Graphic3d,
        CBounds                     from Graphic3d
    
    raises
    
        GroupDefinitionError        from Graphic3d,
        PickIdDefinitionError       from Graphic3d,
    OutOfRange          from Standard
    
    is
        Create ( AStructure : Structure from Graphic3d )
            returns mutable Group from Graphic3d;
        ---Level: Public
        ---Purpose: Creates a group in the structure <AStructure>.
    
        ---------------------------------------------------
        -- Category: Methods to modify the class definition
        ---------------------------------------------------
    
        Clear ( me  : mutable;
                theUpdateStructureMgr : Boolean from Standard = Standard_True )
            is static;
        ---Level: Public
        ---Purpose: Supress all primitives and attributes of <me>.
        --          To clear group without update in Graphic3d_StructureManager
        --          pass Standard_False as <theUpdateStructureMgr>. This
        --          used on context and viewer destruction, when the pointer
        --          to structure manager in Graphic3d_Structure could be 
        --          already released (pointers are used here to avoid handle 
        --          cross-reference);
        ---Category: Methods to modify the class definition
    
        Destroy ( me    : mutable )
            is static;
        ---Level: Public
        ---Purpose: Supress the group <me> in the structure.
        ---Category: Methods to modify the class definition
        ---C++: alias ~
    
        Remove ( me : mutable )
            is static;
        ---Level: Public
        ---Purpose: Supress the group <me> in the structure.
        --  Warning: No more graphic operations in <me> after this call.
        ---Category: Methods to modify the class definition

        --SetTransformPersistence( me     : mutable;
        --                         AFlag  : TransModeFlags from Graphic3d )
        ---Level: Public
    ---Purpose: Modifies the current modelling transform persistence (pan, zoom or rotate)
        --is static;

    --TransformPersistence( me )
    --      returns TransModeFlags from Graphic3d
        ---Level: Public
    ---Purpose: Get the current modelling transform persistence (pan, zoom or rotate)
        --is static;
    
        SetGroupPrimitivesAspect ( me   : mutable )
            is static;
        ---Level: Public
        ---Purpose: Removes the context for all the line primitives
        --      of the group.
        ---Category: Methods to modify the class definition
    
        SetGroupPrimitivesAspect ( me   : mutable;
                                   CTX  : AspectLine3d from Graphic3d )
            is static;
        ---Level: Public
        ---Purpose: Modifies the context for all the line primitives
        --      of the group.
        ---Category: Methods to modify the class definition
    
        SetGroupPrimitivesAspect ( me   : mutable;
                                   CTX  : AspectFillArea3d from Graphic3d )
            is static;
        ---Level: Public
        ---Purpose: Modifies the context for all the face primitives
        --      of the group.
        ---Category: Methods to modify the class definition
    
        SetGroupPrimitivesAspect ( me   : mutable;
                                   CTX  : AspectText3d from Graphic3d )
            is static;
        ---Level: Public
        ---Purpose: Modifies the context for all the text primitives
        --      of the group.
        ---Category: Methods to modify the class definition
    
        SetGroupPrimitivesAspect ( me   : mutable;
                                   CTX  : AspectMarker3d from Graphic3d )
            is static;
        ---Level: Public
        ---Purpose: Modifies the context for all the marker primitives
        --      of the group.
        ---Category: Methods to modify the class definition
    
        SetPrimitivesAspect ( me    : mutable;
                              CTX   : AspectLine3d from Graphic3d )
            is static;
        ---Level: Public
        ---Purpose: Modifies the current context of the group to give
        --      another aspect for all the line primitives created
        --      after this call in the group.
        ---Category: Methods to modify the class definition
    
        SetPrimitivesAspect ( me    : mutable;
                              CTX   : AspectFillArea3d from Graphic3d )
            is static;
        ---Level: Public
        ---Purpose: Modifies the current context of the group to give
        --      another aspect for all the face primitives created
        --      after this call in the group.
        ---Category: Methods to modify the class definition
    
        SetPrimitivesAspect ( me    : mutable;
                              CTX   : AspectText3d from Graphic3d )
            is static;
        ---Level: Public
        ---Purpose: Modifies the current context of the group to give
        --      another aspect for all the text primitives created
        --      after this call in the group.
        ---Category: Methods to modify the class definition
    
        SetPrimitivesAspect ( me    : mutable;
                              CTX   : AspectMarker3d from Graphic3d )
            is static;
        ---Level: Public
        ---Purpose: Modifies the current context of the group to give
        --      another aspect for all the marker primitives created
        --      after this call in the group.
        ---Category: Methods to modify the class definition
    
        SetMinMaxValues ( me                : mutable;
                          XMin, YMin, ZMin  : Real from Standard;
                          XMax, YMax, ZMax  : Real from Standard )
            is static;
        ---Level: Public
        ---Purpose: Sets the coordinates of the boundary box of the
        --      group <me>.
        ---Category: Methods to modify the class definition

        -----------------------------------
        -- Category: Methods to create Text
        -----------------------------------
    
        --------------------------------------------
        -- Summary of Texts                       --
        --                                        --
        -- Text  has  geometric  and nongeometric --
        -- attributes.                            --
        --                                        --
        -- The geometric text attributes are :    --
        --                                        --
        --  Character Height.                 --
        --  Character Up Vector.              --
        --  Text Path.                        --
        --  Text Alignment Horizontal.        --
        --  Text Alignment Vertical.          --
        --                                        --
        -- The nongeometric text attributes are : --
        --                                        --
        --  Text Font.                        --
        --  Character Spacing.                --
        --  Character Expansion Factor.       --
        --  Text Color.                       --
        --------------------------------------------
    
        Text (  me  : mutable;
            AText   : CString from Standard;
            APoint  : Vertex from Graphic3d;
            AHeight : Real from Standard;
            AAngle  : PlaneAngle from Quantity;
            ATp : TextPath from Graphic3d;
            AHta    : HorizontalTextAlignment from Graphic3d;
            AVta    : VerticalTextAlignment from Graphic3d;
            EvalMinMax  : Boolean from Standard = Standard_True )
            is static;
        ---Level: Public
        ---Purpose: Creates the string <AText> at position <APoint>.
        --      The 3D point of attachment is projected. The text is
        --      written in the plane of projection.
        --      The attributes are given with respect to the plane of
        --      projection.
        --      AHeight : Height of text.
        --            (Relative to the Normalized Projection
        --              Coordinates (NPC) Space).
        --      AAngle  : Orientation of the text
        --            (with respect to the horizontal).
        ---Category: Methods to create Text
    
        Text ( me   : mutable;
               AText    : CString from Standard;
               APoint   : Vertex from Graphic3d;
               AHeight  : Real from Standard;
               EvalMinMax   : Boolean from Standard = Standard_True )
            is static;
        ---Level: Public
        ---Purpose: Creates the string <AText> at position <APoint>.
        --      The 3D point of attachment is projected. The text is
        --      written in the plane of projection.
        --      The attributes are given with respect to the plane of
        --      projection.
        --      AHeight : Height of text.
        --            (Relative to the Normalized Projection
        --              Coordinates (NPC) Space).
        --      The other attributes have the following default values:
        --      AAngle  : PI / 2.
        --      ATp     : TP_RIGHT
        --      AHta    : HTA_LEFT
        --      AVta    : VTA_BOTTOM
        ---Category: Methods to create Text
    
        Text (  me          : mutable;
                AText       : ExtendedString from TCollection;
                APoint      : Vertex from Graphic3d;
                AHeight     : Real from Standard;
                AAngle      : PlaneAngle from Quantity;
                ATp         : TextPath from Graphic3d;
                AHta        : HorizontalTextAlignment from Graphic3d;
                AVta        : VerticalTextAlignment from Graphic3d;
                EvalMinMax  : Boolean from Standard = Standard_True )
            is static;
        ---Level: Internal
        ---Purpose: Creates the string <AText> at position <APoint>.
        --      The 3D point of attachment is projected. The text is
        --      written in the plane of projection.
        --      The attributes are given with respect to the plane of
        --      projection.
        --      AHeight : Height of text.
        --            (Relative to the Normalized Projection
        --              Coordinates (NPC) Space).
        --      AAngle  : Orientation of the text
        --            (with respect to the horizontal).
        ---Category: Methods to create Text
    
        Text ( me           : mutable;
               AText        : ExtendedString from TCollection;
               APoint       : Vertex from Graphic3d;
               AHeight      : Real from Standard;
               EvalMinMax   : Boolean from Standard = Standard_True )
            is static;
        ---Level: Internal
        ---Purpose: Creates the string <AText> at position <APoint>.
        --      The 3D point of attachment is projected. The text is
        --      written in the plane of projection.
        --      The attributes are given with respect to the plane of
        --      projection.
        --      AHeight : Height of text.
        --            (Relative to the Normalized Projection
        --              Coordinates (NPC) Space).
        --      The other attributes have the following default values:
        --      AAngle  : PI / 2.
        --      ATp     : TP_RIGHT
        --      AHta    : HTA_LEFT
        --      AVta    : VTA_BOTTOM
        ---Category: Methods to create Text
    
        ---------------------------------------
        ---Category: Methods to create Triangle
        ---------------------------------------

    AddPrimitiveArray( me      : mutable;
                       elem    : ArrayOfPrimitives from Graphic3d;
          EvalMinMax: Boolean from Standard = Standard_True );
        ---Level: Public
    ---Purpose: Adds an array of primitives for display

    UserDraw ( me           : mutable;
               AnObject     : Address from Standard; 
               EvalMinMax   : Boolean from Standard = Standard_True; 
               ContainsFacet: Boolean from Standard = Standard_False
    )
    ---Level: Public
    ---Purpose: Creates an UserDraw primitive
    --  Category: Methods to create UserDraw
    --  Warning: Raises GroupDefinitionError if ...
    raises GroupDefinitionError from Graphic3d is static;

    SetStencilTestOptions (me          : mutable;
                           theIsEnabled: Boolean from Standard);
    ---Purpose: sets the stencil test to theIsEnabled state;

        ----------------------------
        -- Category: Inquire methods
        ----------------------------

        IsGroupPrimitivesAspectSet ( me;
                    theAspect : GroupAspect from Graphic3d )
            returns Boolean from Standard
            is static;
        ---Level: Public
        ---Purpose: Returns TRUE if aspect is set for the group.
        ---Category: Inquire methods

    	GroupPrimitivesAspect ( me;
    				CTXL	: AspectLine3d from Graphic3d;
    				CTXT	: AspectText3d from Graphic3d;
    				CTXM	: AspectMarker3d from Graphic3d;
    				CTXF	: AspectFillArea3d from Graphic3d )
    		is static;
    	---Level: Public
    	---Purpose: Returns the context of all the primitives of the group.
    	---Category: Inquire methods
    
    	PrimitivesAspect ( me;
    			   CTXL	: AspectLine3d from Graphic3d;
    			   CTXT	: AspectText3d from Graphic3d;
    			   CTXM	: AspectMarker3d from Graphic3d;
    			   CTXF	: AspectFillArea3d from Graphic3d )
    		is static;
    	---Level: Public
    	---Purpose: Returns the last inserted context in the group <me>
    	--	    foreach kind of primitives.
    	---Category: Inquire methods

        ContainsFacet ( me )
            returns Boolean from Standard
            is static;
        ---Level: Internal
        ---Purpose: Returns Standard_True if the group <me> contains
        --      Polygons, Triangles or Quadrangles.
        ---Category: Inquire methods
    
        IsDeleted ( me )
            returns Boolean from Standard
            is static;
        ---Level: Public
        ---Purpose: Returns Standard_True if the group <me> is deleted.
        --      <me> is deleted after the call Remove (me) or the
        --      associated structure is deleted.
        ---Category: Inquire methods
    
        IsEmpty ( me )
            returns Boolean from Standard
            is static;
        ---Level: Public
        ---Purpose: Returns Standard_True if the group <me> is empty.
        ---Warning: A group is empty if the MinMaxValues method returns :
        --      XMin = YMin = ZMin = RealFirst ().
        --      XMax = YMax = ZMax = RealLast ().
        ---Category: Inquire methods
    
        MinMaxValues ( me;
                       XMin, YMin, ZMin : out Real from Standard;
                       XMax, YMax, ZMax : out Real from Standard )
            is static;
        ---Level: Public
        ---Purpose: Returns the coordinates of the boundary box of the
        --      group <me>.
        ---Warning: If the group <me> is empty then :
        --      XMin = YMin = ZMin = RealFirst ().
        --      XMax = YMax = ZMax = RealLast ().
        ---Category: Inquire methods
    
        Structure ( me )
            returns mutable Structure from Graphic3d
            is static;
        ---Level: Public
        ---Purpose: Returns the structure containing the group <me>.
        ---Category: Inquire methods
    
        ----------------------------
        -- Category: Private methods
        ----------------------------
        
        MinMaxCoord ( me;
                      XMin, YMin, ZMin : out Real from Standard;
                      XMax, YMax, ZMax : out Real from Standard )
            is static private;
        ---Level: Internal
        ---Purpose: Returns the extreme coordinates found in the group.
        ---Warning: If the group <me> is empty then :
        --      XMin = YMin = ZMin = RealFirst ().
        --      XMax = YMax = ZMax = RealLast ().
        ---Category: Private methods
    
        Update ( me )
            is static private;
        ---Level: Internal
        ---Purpose: Calls the Update method of the StructureManager which
        --      contains the associated Structure of the Group <me>.
        ---Category: Private methods
    
    fields
    
    --
    -- Class    :   Graphic3d_Group
    --
    -- Purpose  :   Declaration of variables specific to groups
    --          of primitives.
    --
    -- Reminder :   A group is defined in a structure
    --          It acts as the smallest editable entity.
    
        -- the associated C structure 
        MyCGroup        :   CGroup from Graphic3d;
    
        -- the graphic driver used
        MyGraphicDriver     :   GraphicDriver from Graphic3d;
    
        -- the state of the different contexts for primitives
        MyCBitFields        :   CBitFields4 from Graphic3d;
    
        -- the structure contains the group
        MyPtrStructure      :   Address from Standard;
    
        -- the min-max
    MyBounds                :       CBounds from Graphic3d;

    MyListOfPArray          :   ListOfPArray from Graphic3d;

    MyMarkArray             :       HArray1OfByte from TColStd;
    MyMarkWidth             :       Integer from Standard;
    MyMarkHeight            :       Integer from Standard;

    friends
    
        Remove from class Structure from Graphic3d
            ( me : mutable; AGroup : Group from Graphic3d )
    
    end Group;
