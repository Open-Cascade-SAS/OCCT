-- File:	TDataStd_DeltaOnModificationOfRealArray.cdl
-- Created:	Tue Oct 30 16:49:40 2007
-- Author:	Sergey ZARITCHNY
--		<sergey.zaritchny@opencascade.com>
---Copyright:	Open CasCade SA 2007


class DeltaOnModificationOfRealArray from TDataStd inherits DeltaOnModification from TDF

	---Purpose: This class provides default services for an
	--          AttributeDelta on a MODIFICATION action

uses

    Attribute      from TDF,
    HArray1OfReal  from TColStd,
    HArray1OfInteger from TColStd,
    RealArray      from TDataStd

is

    Create (Arr : RealArray     from TDataStd)
    	returns mutable DeltaOnModificationOfRealArray from TDataStd;
	---Purpose: Initializes a TDF_DeltaOnModification.

    Apply (me : mutable)
    	is redefined virtual;
    	---Purpose: Applies the delta to the attribute.
fields
  
 myIndxes  :  HArray1OfInteger from TColStd; 
 myValues  :  HArray1OfReal from TColStd;
 myUp1     :  Integer       from Standard;
 myUp2     :  Integer       from Standard;

end DeltaOnModificationOfRealArray;
