-- Created on: 1992-09-23
-- Created by: Christian CAILLET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class GraphContent  from Interface  inherits EntityIterator

    	---Purpose : Defines general form for classes of graph algorithms on
    	--           Interfaces, this form is that of EntityIterator
    	--           Each sub-class fills it according to its own algorithm
    	--           This also allows to combine any graph result to others,
    	--           all being given under one unique form

uses Transient, Graph

is

    Create returns GraphContent;
    ---Purpose : Creates an empty GraphContent, ready to be filled

    Create (agraph : Graph) returns GraphContent;
    ---Purpose : Creates with all entities designated by a Graph

    Create (agraph : Graph; stat : Integer) returns GraphContent;
    ---Purpose : Creates with entities having specific Status value in a Graph

    Create (agraph : Graph; ent : Transient) returns GraphContent;
    ---Purpose : Creates an Iterator with Shared entities of an entity
    --           (equivalente to EntityIterator but with a Graph) 

    GetFromGraph (me : in out; agraph : Graph);
    ---Purpose : Gets all Entities designated by a Graph (once created), adds
    --           them to those already recorded

    GetFromGraph (me : in out; agraph : Graph; stat : Integer);
    ---Purpose : Gets entities from a graph which have a specific Status value
    --           (one created), adds them to those already recorded

    Result (me : in out) returns EntityIterator;
    ---Purpose : Returns Result under the exact form of an EntityIterator :
    --           Can be used when EntityIterator itself is required (as a
    --           returned value for instance), whitout way for a sub-class

    	-- --    Evaluation - Iteration    -- --
    	--   Made by Start-More-Next-Value  inherited from EntityIterator
    	--   Start is redefined to call Evaluate moreover
    	--   Default for Evaluate is given as doing nothing

--    Start (me : in out)  is redefined;
    Begin (me : in out);
    ---Purpose : Does the Evaluation before starting the iteration itself
    --           (in out)

    Evaluate (me : in out)  is virtual;
    ---Purpose : Evaluates list of Entities to be iterated. Called by Start
    --           Default is set to doing nothing : intended to be redefined
    --           by each sub-class

end GraphContent;
