-- File:	StepBasic_EffectivityAssignment.cdl
-- Created:	Wed May 10 15:09:06 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class EffectivityAssignment from StepBasic
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity EffectivityAssignment

uses
    Effectivity from StepBasic

is
    Create returns EffectivityAssignment from StepBasic;
	---Purpose: Empty constructor

    Init (me: mutable; aAssignedEffectivity: Effectivity from StepBasic);
	---Purpose: Initialize all fields (own and inherited)

    AssignedEffectivity (me) returns Effectivity from StepBasic;
	---Purpose: Returns field AssignedEffectivity
    SetAssignedEffectivity (me: mutable; AssignedEffectivity: Effectivity from StepBasic);
	---Purpose: Set field AssignedEffectivity

fields
    theAssignedEffectivity: Effectivity from StepBasic;

end EffectivityAssignment;
