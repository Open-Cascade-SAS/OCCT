-- Created on: 1994-06-24
-- Created by: Frederic MAUPAS
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MakeShellBasedSurfaceModel from TopoDSToStep inherits
    Root from TopoDSToStep

    ---Purpose: This class implements the mapping between classes 
    --          Face, Shell or Solid from TopoDS and ShellBasedSurfaceModel
    --          from StepShape. All the topology and geometry comprised 
    --          into the shape are taken into account and translated.
  
uses Face  from TopoDS,
     Shell from TopoDS,
     Solid from TopoDS,
     ShellBasedSurfaceModel from StepShape,
     FinderProcess from Transfer
          
raises NotDone from StdFail
     
is 

Create ( F  : Face from TopoDS;
         FP : FinderProcess from Transfer)
        returns MakeShellBasedSurfaceModel;

Create ( S           : Shell from TopoDS;
         FP          : FinderProcess from Transfer)
        returns MakeShellBasedSurfaceModel;

Create ( S  : Solid from TopoDS;
         FP : FinderProcess from Transfer)
        returns MakeShellBasedSurfaceModel;

Value (me) returns ShellBasedSurfaceModel from StepShape
    raises NotDone
    is static;
    ---C++: return const&

fields

    theShellBasedSurfaceModel : ShellBasedSurfaceModel from StepShape;

    	-- The solution from StepShape
    	
end MakeShellBasedSurfaceModel;

