-- File:	IGESDimen_ToolNewGeneralNote.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolNewGeneralNote  from IGESDimen

    ---Purpose : Tool to work on a NewGeneralNote. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses NewGeneralNote from IGESDimen,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolNewGeneralNote;
    ---Purpose : Returns a ToolNewGeneralNote, ready to work


    ReadOwnParams (me; ent : mutable NewGeneralNote;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : NewGeneralNote;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : NewGeneralNote;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a NewGeneralNote <ent>, from
    --           its specific (own) parameters

    DirChecker (me; ent : NewGeneralNote) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : NewGeneralNote;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : NewGeneralNote; entto : mutable NewGeneralNote;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : NewGeneralNote;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolNewGeneralNote;
