-- File:	PGeom_Axis1Placement.cdl
-- Created:	Mon Feb 22 16:04:21 1993
-- Author:	Philippe DAUTRY
--		<fid@phobox>
-- Copyright:	 Matra Datavision 1993


class Axis1Placement from PGeom inherits AxisPlacement from PGeom

	---Purpose : This class describes an axis  one placement built
	--         with a point and a direction.
	--          

uses Ax1 from gp

is


  Create returns mutable Axis1Placement from PGeom;
        --- Purpose : Creates an Axis1Placement with Ax1 default value.
    	---Level: Internal 

  Create (aAxis : Ax1 from gp) returns mutable Axis1Placement from PGeom;
        --- Purpose : Creates an Axis1Placement with <aAxis>.
    	---Level: Internal 


end;


