-- Created on: 1996-02-13
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class MakeRevol from BRepFeat inherits Form from BRepFeat

	---Purpose: Describes functions to build revolved shells from basis shapes.

uses Shape                     from TopoDS,
     Face                      from TopoDS,
     Edge                      from TopoDS,
     DataMapOfShapeListOfShape from TopTools,
     Ax1                       from gp,
     DataMapOfShapeShape       from TopTools,
     SequenceOfCurve           from TColGeom,
     Curve                     from Geom,
     SequenceOfCurve           from TColGeom,
     StatusError               from BRepFeat
     
    raises ConstructionError from Standard

is


    Create

    	returns MakeRevol from BRepFeat;
	---Purpose: initializes the revolved shell class.
	---C++: inline


    Create(Sbase     : Shape   from TopoDS;
           Pbase     : Shape   from TopoDS;
           Skface    : Face    from TopoDS;
	   Axis      : Ax1     from gp;
           Fuse      : Integer from Standard;
           Modify    : Boolean from Standard)
    
	---Purpose: a face Pbase is selected in the
    	--   shape Sbase to serve as the basis for the
    	--   revolved shell. The revolution will be defined
    	--   by the axis Axis and Fuse offers a choice between:
    	--   -   removing matter with a Boolean cut using the setting 0
    	--   -   adding matter with Boolean fusion using the setting 1.
    	--     The sketch face Skface serves to determine
    	-- the type of operation. If it is inside the basis
    	-- shape, a local operation such as glueing can be performed.
    	---C++: inline
    	    	returns MakeRevol from BRepFeat;


    Init(me: in out; Sbase     : Shape   from TopoDS;
                     Pbase     : Shape   from TopoDS;
                     Skface    : Face    from TopoDS;
                     Axis      : Ax1     from gp;
	             Fuse      : Integer from Standard;
                     Modify    : Boolean from Standard)
    
    	is static;


    Add(me: in out; E: Edge from TopoDS; OnFace: Face from TopoDS)

	---Purpose: Indicates that the edge <E> will slide on the face
	-- <OnFace>. Raises ConstructionError if the  face does not belong to the
	-- basis shape, or the edge to the prismed shape.
    	raises ConstructionError from Standard
	
	is static;


    Perform(me: in out; Angle: Real from Standard)
    
    	is static;


    Perform(me: in out; Until: Shape from TopoDS)
    
    	is static;


    Perform(me: in out; From : Shape from TopoDS;
                        Until: Shape from TopoDS)
    
    	is static;
    	---Purpose: Reconstructs the feature topologically.

    PerformThruAll(me: in out)
    
    	is static;
    	---Purpose: Builds an infinite shell. The infinite descendants
    	-- will not be kept in the result.

    PerformUntilAngle(me: in out; Until :  Shape from TopoDS;
                        Angle :  Real  from Standard)
    
    	is static;
    	---Purpose: Assigns both a limiting shape, Until from
    	-- TopoDS_Shape, and an angle, Angle at
    	-- which to stop generation of the revolved shell feature.
    Curves(me: in out; S : in out SequenceOfCurve from TColGeom);
    

    BarycCurve(me: in out)    
    	returns Curve from Geom;


fields

    myPbase  : Shape                     from TopoDS;
    mySlface : DataMapOfShapeListOfShape from TopTools;
    myAxis   : Ax1                       from gp;
    myCurves : SequenceOfCurve           from TColGeom;
    myBCurve : Curve                     from Geom;
    myStatusError : StatusError          from BRepFeat;

end MakeRevol;
