-- Created on: 1997-07-25
-- Created by: Jerome LEMONIER
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class AppFuncRst from BRepBlend inherits AppFuncRoot from BRepBlend
	---Purpose: Function to approximate by AppSurface for Edge/Face          
	---Level: Advanced

uses 
 Line            from BRepBlend,
 Point           from Blend,
 SurfRstFunction from Blend,
 AppFunction     from Blend,
 Vector          from math

 
raises OutOfRange from  Standard

is   
     
   Create(Line : in out Line from BRepBlend;
    	  Func  : in  out SurfRstFunction from Blend; 
          Tol3d: Real;
          Tol2d: Real)
   returns AppFuncRst from BRepBlend;

   Point(me;
    	 Func  : AppFunction from Blend; 
	 Param : Real;
	 Sol   : Vector from math;
	 Pnt   : in out Point from Blend);
	
   Vec(me;
       Sol : in out Vector from math;
       Pnt : Point from Blend);
	
end AppFuncRst;
