-- Created by: DAUTRY Philippe
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

--      	-----------------------

---Version:	0.0
--Version	Date		Purpose
--		0.0	May  7 1997	Creation



generic class RelocationTable from MDF
    (TheSourceType as any;
     TheTargetType as any;
     TheOtherSourceType as any;
     TheOtherTargetType as any;
     TheMapType    as any)
    inherits TShared from MMgt

	---Purpose: Storage Relocation Table
	--          (Transient->Persistent). It is a relocation
	--          dictionnary.

uses

    Tool from MDF

-- raises

is

    Create(theSelfRelocation : Boolean from Standard = Standard_False) 
    returns mutable RelocationTable from MDF;
	---Purpose: Creates a relocation table. 
	--          <theSelfRelocation> status says that the relocation table allows self relocation.

    SetSelfRelocation(me : mutable; theStatus : Boolean from Standard = Standard_True);
    ---Purpose: Sets self relocation status.

    IsSelfRelocation(me) 
    ---Purpose: Returns true if the self relocation status is set.
    returns Boolean from Standard;


    -- Attribute relocation methods.
    -- ---------

    SetRelocation(me : mutable;
    	    	  aSourceAttribute : TheSourceType;
    	    	  aTargetAttribute : TheTargetType);
	---Purpose: Sets the relocation value of <aSourceAttribute> to
	--          <aTargetAttribute>.

    HasRelocation(me : mutable;
    	    	  aSourceAttribute :                TheSourceType;
    	    	  aTargetAttribute : in out mutable TheTargetType)
	returns Boolean from Standard;
	---Purpose: Finds the relocation value of <aSourceAttribute>
	--          and returns it into <aTargetAttribute>.
	--          
	--          If a value is found, returns True; False otherwise.


    -- Transient other types object relocation methods.
    -- ---------------------

    SetOtherRelocation(me : mutable;
    	               aSource : TheOtherSourceType;
    	               aTarget : TheOtherTargetType);
	---Purpose: Sets the relocation value of <aSourceTransient> to
	--          <aTargetTransient>.

    HasOtherRelocation(me : mutable;
    	    	       aSource :                TheOtherSourceType;
    	    	       aTarget : in out mutable TheOtherTargetType)
	returns Boolean from Standard;
	---Purpose: Finds the relocation value of <aSource>
	--          and returns it into <aTarget>.
	--          
	--          If a value is found, returns True; False otherwise.


    -- Try not to use the following methods...

    AttributeTable(me : mutable)
    	returns TheMapType;
	---Purpose: Returns <myAttributeTable> to be read or
	--          updated. Please, for a better security, avoid to
	--          use this method.
	--          
	---C++: return &

    OtherTable(me : mutable)
    	returns TheMapType;
	---Purpose: Returns <myOtherTable> to be read or
	--          updated. Please, for a better security, avoid to
	--          use this method.
	--          
	---C++: return &


fields

    myAttributeTable : TheMapType;
    myOtherTable     : TheMapType;
    mySelfRelocation : Boolean from Standard;

end RelocationTable;
