--
-- File:	Aspect_Background.cdl
-- Created:	Mercredi 2 Octobre 1991
-- Author:	NW,JPB,CAL
--
---Copyright:	MatraDatavision 1991,1992,1993
--

class Background from Aspect


	---Purpose: This class allows the definition of
	--	    a window background.

uses

	Color	from Quantity

is

	Create
		returns Background from Aspect;
	---Level: Public
	---Purpose: Creates a window background.
	--	    Default color : NOC_MATRAGRAY.

	Create ( AColor : Color from Quantity )
		returns Background from Aspect;
	---Level: Public
	---Purpose: Creates a window background with the colour <AColor>.

	---------------------------------------------------
	-- Category: Methods to modify the class definition
	---------------------------------------------------

	SetColor ( me		: in out;
		   AColor	: Color from Quantity );
	---Level: Public
	---Purpose: Modifies the colour of the window background <me>.
	---Category: Methods to modify the class definition

	----------------------------
	-- Category: Inquire methods
	----------------------------

	Color ( me )
		returns Color from Quantity;
	---Level: Public
	---Purpose: Returns the colour of the window background <me>.
	---Category: Inquire methods

--

fields

--
-- Class	:	Aspect_Background
--
-- Purpose	:	Declaration of variables specific to the window
--			background.
--
-- Reminder	:	A background is defined by one colour
--

	-- the colour associated with the window background
	MyColor	:	Color from Quantity;

end Background;
