-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Axis2Placement2d from StepGeom 

inherits Placement from StepGeom 

uses

	Direction from StepGeom, 
	Boolean from Standard, 
	HAsciiString from TCollection, 
	CartesianPoint from StepGeom
is

	Create returns Axis2Placement2d;
	---Purpose: Returns a Axis2Placement2d


	Init (me : mutable;
	      aName : HAsciiString from TCollection;
	      aLocation : CartesianPoint from StepGeom) is redefined;

	Init (me : mutable;
	      aName : HAsciiString from TCollection;
	      aLocation : CartesianPoint from StepGeom;
	      hasArefDirection : Boolean from Standard;
	      aRefDirection : Direction from StepGeom) is virtual;

	-- Specific Methods for Field Data Access --

	SetRefDirection(me : mutable; aRefDirection : Direction);
	UnSetRefDirection (me:mutable);
	RefDirection (me) returns Direction;
	HasRefDirection (me) returns Boolean;

fields

	refDirection : Direction from StepGeom;   -- OPTIONAL can be NULL
	hasRefDirection : Boolean from Standard;

end Axis2Placement2d;
