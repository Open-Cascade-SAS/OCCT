-- Created on: 1992-12-02
-- Created by: Isabelle GRIGNON
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class CelGProps  from GProp inherits GProps from GProp

	--- Purpose  : 
	--  Computes the  global properties of bounded curves 
	--  in 3D space. 
	--  It can be an elementary curve from package gp such as 
	--  Lin, Circ, Elips, Parab .

uses  Circ  from gp,
      Lin   from gp,
      Parab from gp,
      Pnt   from gp
       
is

    Create returns CelGProps;
  
    Create (C : Circ from gp; CLocation : Pnt)   returns CelGProps;

    Create (C : Circ from gp; U1, U2 : Real; CLocation : Pnt)returns CelGProps;

    Create (C : Lin from gp; U1, U2 : Real; CLocation : Pnt) returns CelGProps;

    SetLocation(me : in out;CLocation : Pnt) ;

    Perform(me : in out; C :Circ; U1,U2 : Real);
    
    Perform(me : in out; C : Lin ; U1,U2 : Real);

end CelGProps;


