-- File:	MPrsStd_PositionRetrievalDriver.cdl
-- Created:	Tue Apr  7 14:58:29 1998
-- Author:	Jean-Pierre COMBE
--		<jpr@chariox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1998

class PositionRetrievalDriver from MPrsStd inherits ARDriver from MDF
	---Purpose: 



uses RRelocationTable from MDF,
     Attribute        from PDF,
     Attribute        from TDF, 
     MessageDriver    from CDM

is


    Create(theMessageDriver : MessageDriver from CDM)  -- Version 0
    returns mutable PositionRetrievalDriver from MPrsStd;
    

    VersionNumber(me) returns Integer from Standard;
	---Purpose: Returns the version number from which the driver
	--          is available: 0.

    SourceType(me) returns Type from Standard;
	---Purpose: Returns the type: ColorAttribute from PGraphicAttribute.

    NewEmpty (me)  returns mutable Attribute from TDF;


    Paste(me;
    	  Source     :         Attribute from PDF;
    	  Target     : mutable Attribute from TDF;
    	  RelocTable : RRelocationTable  from MDF);

end PositionRetrievalDriver;
