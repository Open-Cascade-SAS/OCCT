-- Created on: 1999-11-05
-- Created by: Vladislav ROMASHKO
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Revol from QANewBRepNaming inherits TopNaming from QANewBRepNaming 

    ---Purpose: To load the Revol results 

uses 
 
    MakeRevol from BRepPrimAPI, 
    Shape     from TopoDS,
    Label     from TDF

is 
 
    Create returns Revol from QANewBRepNaming;

    Create(ResultLabel : Label from TDF) 
    returns Revol from QANewBRepNaming;

    Init(me : in out; ResultLabel : Label from TDF);


    Load (me; mkRevol : in out MakeRevol from BRepPrimAPI;
	      basis   : in     Shape     from TopoDS);
    ---Purpose: Loads the revol in the data framework 
      
    Start(me)
    ---Purpose: Returns the insertion label of the start face of the Revol.  
    returns Label from TDF;

    End(me) 
    ---Purpose: Returns the insertion label of the end face of the Revol. 
    returns Label from TDF;
       
    Lateral(me) 
    ---Purpose: Returns the insertion label of the lateral faces of the Revol.
    returns Label from TDF; 
    
    Degenerated(me)
    ---Purpose: Returns the label of degenerated edges.
    returns Label from TDF;
    
    Content(me)
    ---Purpose: Returns the label of the content of the result.
    returns Label from TDF;    
    

end Revol;
