-- Created on: 1997-03-27
-- Created by: Denis PASCAL
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



package DDataStd 

	---Purpose: commands for Standard Attributes.
	--          =================================


uses Draw,
     TDF,
     TDataStd,     
     TDataXtd,
     TopoDS,
     MMgt,
     Standard,
     TNaming, 
     TCollection

is 

    ---Purpose: attribute display presentation
    --          ==============================

    class DrawPresentation;
    
    class DrawDriver;
    ---Purpose: root class of drivers to build draw variables from TDF_Label.

   ---Purpose: attribute tree presentation
    --         ===========================

    class TreeBrowser;
    ---Purpose: Used to browse tree nodes.

    ---Purpose: commands
    --          ========

    AllCommands (I : in out Interpretor from Draw);
    ---Purpose: command to set and get modeling attributes

    NamedShapeCommands (I : in out Interpretor from Draw);
    ---Purpose: to set and get NamedShape

    BasicCommands  (I : in out Interpretor from Draw);
    ---Purpose: to set and get Integer, Real,  Reference, Geometry

    DatumCommands (I : in out Interpretor from Draw);
    ---Purpose: to set and get Datum attributes

    ConstraintCommands (I : in out Interpretor from Draw);
    ---Purpose: to set and get Constraint and Constraint  attributes    

    ObjectCommands (I : in out Interpretor from Draw);
    ---Purpose: to set and get Objects attributes

    DrawDisplayCommands  (I : in out Interpretor from Draw);
    ---Purpose: to display standard attributes

    NameCommands (I: in out Interpretor from Draw);
    ---Purpose: to set and get Name attribute    
    
    TreeCommands (I: in out Interpretor from Draw);    
    ---Purpose: to build, edit and browse an explicit tree of labels
    
    ---Purpose: package methods
    --          ===============

    DumpConstraint (C : Constraint from TDataXtd; S : in out OStream);


end DDataStd;

