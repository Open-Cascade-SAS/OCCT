-- File:	StepRepr_StructuralResponsePropertyDefinitionRepresentation.cdl
-- Created:	Sun Dec 15 10:59:25 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class StructuralResponsePropertyDefinitionRepresentation from StepRepr
inherits PropertyDefinitionRepresentation from StepRepr

    ---Purpose: Representation of STEP entity StructuralResponsePropertyDefinitionRepresentation

uses
    PropertyDefinition from StepRepr,
    Representation from StepRepr

is
    Create returns StructuralResponsePropertyDefinitionRepresentation from StepRepr;
	---Purpose: Empty constructor

end StructuralResponsePropertyDefinitionRepresentation;
