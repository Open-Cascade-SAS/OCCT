-- Created on: 1996-12-26
-- Created by: Alexander BRIVIN and Dmitry TARASOV
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class IndexedFaceSet from Vrml inherits  TShared  from  MMgt

	---Purpose: defines a IndexedFaceSet node of VRML specifying geometry shapes. 
    	--  This node represents a 3D shape formed by constructing faces (polygons) from  
    	--  vertices located at the current coordinates. IndexedFaceSet uses the indices  
    	--  in its coordIndex to define polygonal faces. An index of -1 separates faces  
    	--  (so a -1 at the end of the list is optional). 

    	--  The vertices of the faces are transformed by the current transformation matrix. 
        --  Treatment of the current material and normal binding is as follows: The PER_PART  
    	--  and PER_FACE bindings specify a material or normal for each face. PER_VERTEX  
    	--  specifies a material or normal for each vertex. The corresponding _INDEXED bindings  
    	--  are the same, but use the materialIndex or normalIndexindices. The DEFAULT material  
    	--  binding is equal to OVERALL. The DEFAULT normal binding is equal to PER_VERTEX_INDEXED;  
    	--  if insufficient normals exist in the state, vertex normals will be generated
	--  automatically. When materialIndex or normalIndex are specified on a per vertex basis,  
    	--  an index of -1 is used in the same way as coordIndex.
uses

    HArray1OfInteger from TColStd

is

    Create ( aCoordIndex        : HArray1OfInteger from TColStd;
    	     aMaterialIndex     : HArray1OfInteger from TColStd;
	     aNormalIndex       : HArray1OfInteger from TColStd;
	     aTextureCoordIndex : HArray1OfInteger from TColStd )
        returns mutable IndexedFaceSet from Vrml;

    Create  returns mutable IndexedFaceSet from Vrml; 
    
    SetCoordIndex ( me : mutable; aCoordIndex : HArray1OfInteger from TColStd );
    CoordIndex ( me )  returns HArray1OfInteger from TColStd;
    
    SetMaterialIndex ( me : mutable; aMaterialIndex : HArray1OfInteger from TColStd );
    MaterialIndex ( me )  returns HArray1OfInteger from TColStd;
    
    SetNormalIndex ( me : mutable; aNormalIndex : HArray1OfInteger from TColStd );
    NormalIndex ( me )  returns HArray1OfInteger from TColStd;
    
    SetTextureCoordIndex ( me : mutable; 
    	aTextureCoordIndex : HArray1OfInteger from TColStd );
    TextureCoordIndex ( me )  returns HArray1OfInteger from TColStd;
   
    Print  ( me; anOStream: in out OStream from Standard) returns OStream from Standard;
    ---C++:  return  & 

fields

    myCoordIndex        : HArray1OfInteger from TColStd;  -- Coordinate indices
    myMaterialIndex     : HArray1OfInteger from TColStd;  -- Material indices
    myNormalIndex       : HArray1OfInteger from TColStd;  -- Surface normal indices
    myTextureCoordIndex : HArray1OfInteger from TColStd;  -- Texture Coordinate indices

end IndexedFaceSet;
