-- Created on: 1998-10-29
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Hctxff2d from TopOpeBRep inherits TShared from  MMgt

uses

    Shape from TopoDS,
    Face from TopoDS,
    HSurface from BRepAdaptor,
    Surface from BRepAdaptor,
    SurfaceType from GeomAbs

is

    Create returns mutable Hctxff2d from TopOpeBRep;
    SetFaces(me:mutable; F1,F2:Face);
    SetHSurfaces(me:mutable; S1,S2:HSurface from BRepAdaptor);
    SetHSurfacesPrivate(me:mutable) is private;
    SetTolerances(me:mutable;Tol1,Tol2:Real);
    GetTolerances(me;Tol1,Tol2:out Real);
    GetMaxTolerance(me) returns Real;
    Face(me;I:Integer) returns Face;---C++ : return const &
    HSurface(me;I:Integer) returns HSurface from BRepAdaptor;
    SurfacesSameOriented(me) returns Boolean;
    FacesSameOriented(me) returns Boolean;
    FaceSameOrientedWithRef(me;I:Integer) returns Boolean;

fields

    myFace1 : Face from TopoDS;
    mySurface1 : HSurface from BRepAdaptor;
    mySurfaceType1 : SurfaceType from GeomAbs;
    myf1surf1F_sameoriented : Boolean;

    myFace2 : Face from TopoDS;
    mySurface2 : HSurface from BRepAdaptor;
    mySurfaceType2 : SurfaceType from GeomAbs;
    myf2surf1F_sameoriented : Boolean;

    mySurfacesSameOriented : Boolean;
    myFacesSameOriented : Boolean;
    
    myTol1,myTol2 : Real;
    
end Hctxff2d from TopOpeBRep;
