-- Created on: 2012-03-23
-- Created by: DBV
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package QABugs
uses
    Draw,
    TCollection, 
    gp, 
    PrsMgr, 
    Prs3d,
    Quantity,
    SelectMgr,
    AIS
is 
    class  MyText;
    class  PresentableObject;
    
    Commands(DI : in out Interpretor from Draw);
    Commands_1(DI : in out Interpretor from Draw);
    Commands_2(DI : in out Interpretor from Draw);
    Commands_3(DI : in out Interpretor from Draw);
    Commands_4(DI : in out Interpretor from Draw);
    Commands_5(DI : in out Interpretor from Draw);
    Commands_6(DI : in out Interpretor from Draw);
    Commands_7(DI : in out Interpretor from Draw);
    Commands_8(DI : in out Interpretor from Draw);
    Commands_9(DI : in out Interpretor from Draw);
    Commands_10(DI : in out Interpretor from Draw);
    Commands_11(DI : in out Interpretor from Draw);
    Commands_12(DI : in out Interpretor from Draw);
    Commands_13(DI : in out Interpretor from Draw);
    Commands_14(DI : in out Interpretor from Draw);
    Commands_15(DI : in out Interpretor from Draw);
    Commands_16(DI : in out Interpretor from Draw);
    Commands_17(DI : in out Interpretor from Draw);
    Commands_18(DI : in out Interpretor from Draw);
    Commands_19(DI : in out Interpretor from Draw);
end;
