-- File:	IGESDimen_ToolDimensionDisplayData.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolDimensionDisplayData  from IGESDimen

    ---Purpose : Tool to work on a DimensionDisplayData. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses DimensionDisplayData from IGESDimen,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolDimensionDisplayData;
    ---Purpose : Returns a ToolDimensionDisplayData, ready to work


    ReadOwnParams (me; ent : mutable DimensionDisplayData;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : DimensionDisplayData;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : DimensionDisplayData;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a DimensionDisplayData <ent>, from
    --           its specific (own) parameters

    OwnCorrect (me; ent : mutable DimensionDisplayData) returns Boolean  is static;
    ---Purpose : Sets automatic unambiguous Correction on a DimensionDisplayData
    --           (NbPropertyValues forced to 14)

    DirChecker (me; ent : DimensionDisplayData) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : DimensionDisplayData;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : DimensionDisplayData; entto : mutable DimensionDisplayData;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : DimensionDisplayData;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolDimensionDisplayData;
