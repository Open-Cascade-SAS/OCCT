-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class GlobalUncertaintyAssignedContext from StepRepr 

inherits RepresentationContext from StepRepr 

uses

	HArray1OfUncertaintyMeasureWithUnit from StepBasic, 
	UncertaintyMeasureWithUnit from StepBasic, 
	HAsciiString from TCollection
is

	Create returns mutable GlobalUncertaintyAssignedContext;
	---Purpose: Returns a GlobalUncertaintyAssignedContext


	Init (me : mutable;
	      aContextIdentifier : mutable HAsciiString from TCollection;
	      aContextType : mutable HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      aContextIdentifier : mutable HAsciiString from TCollection;
	      aContextType : mutable HAsciiString from TCollection;
	      aUncertainty : mutable HArray1OfUncertaintyMeasureWithUnit from StepBasic) is virtual;

	-- Specific Methods for Field Data Access --

	SetUncertainty(me : mutable; aUncertainty : mutable HArray1OfUncertaintyMeasureWithUnit);
	Uncertainty (me) returns mutable HArray1OfUncertaintyMeasureWithUnit;
	UncertaintyValue (me; num : Integer) returns mutable UncertaintyMeasureWithUnit;
	NbUncertainty (me) returns Integer;

fields

	uncertainty : HArray1OfUncertaintyMeasureWithUnit from StepBasic;

end GlobalUncertaintyAssignedContext;
