-- File:        PresentationView.cdl
-- Created:     Fri Dec  1 11:11:25 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class PresentationView from StepVisual 

inherits PresentationRepresentation from StepVisual 

uses

	HAsciiString from TCollection, 
	HArray1OfRepresentationItem from StepRepr,
	RepresentationContext from StepRepr
is

	Create returns mutable PresentationView;
	---Purpose: Returns a PresentationView


end PresentationView;
