-- Created on: 1997-01-22
-- Created by: Mister rmi
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Driver from FWOSDriver  inherits MetaDataDriver from CDF
uses
    MetaData from CDM,Document from CDM,
    ExtendedString from TCollection,
    ExtendedString from TCollection
is
    Create
    returns mutable Driver from FWOSDriver;
    ---Purpose: initializes the MetaDatadriver with its specific name.


    	
    Find(me: mutable; aFolder, aName, aVersion: ExtendedString from TCollection)
    returns Boolean from Standard;
    ---Purpose: indicate whether a file exists corresponding to the folder and the name
    
    HasReadPermission(me: mutable; aFolder, aName, aVersion: ExtendedString from TCollection)
    returns Boolean from Standard;

    
    MetaData(me: mutable; aFolder, aName, aVersion: ExtendedString from TCollection)
    returns MetaData from CDM
    is  private;
    
    CreateMetaData(me: mutable; aDocument: Document from CDM;
    	         aFileName: ExtendedString from TCollection)
    returns  MetaData from CDM
    is  private;
    
    FindFolder(me: mutable; aFolder: ExtendedString from TCollection)
    returns Boolean from Standard;


   DefaultFolder(me: mutable) returns ExtendedString from TCollection;
   
   BuildFileName(me: mutable; aDocument: Document from CDM)
   returns ExtendedString from TCollection;
    
   Concatenate(myclass; aFolder,aName:  ExtendedString from TCollection)
   returns ExtendedString from TCollection
   is private;


   BuildMetaData(me: mutable; aFileName: ExtendedString from TCollection)
   returns MetaData from CDM
   is  private;

   SetName(me: mutable; aDocument: Document from CDM; aName: ExtendedString from TCollection)
   returns ExtendedString from TCollection
   is redefined;
   
end Driver from FWOSDriver;
