-- Created on: 2000-08-15
-- Created by: data exchange team
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package MXCAFDoc 

	---Purpose: 

uses
    TopLoc,
    PTopLoc,
    TDF,
    PDF,
    MDF,
    MDataStd,
    CDM

is
    class DocumentToolRetrievalDriver;
    class DocumentToolStorageDriver;
    class ColorToolRetrievalDriver;
    class ColorToolStorageDriver;
    class ShapeToolRetrievalDriver;
    class ShapeToolStorageDriver;

    class LayerToolRetrievalDriver;
    class LayerToolStorageDriver;
    
    class LocationStorageDriver;
    class LocationRetrievalDriver;
    class ColorStorageDriver;
    class ColorRetrievalDriver;
    class VolumeStorageDriver;
    class VolumeRetrievalDriver;
    class AreaStorageDriver;
    class AreaRetrievalDriver;
    class CentroidStorageDriver;
    class CentroidRetrievalDriver;
    
    class GraphNodeStorageDriver;
    class GraphNodeRetrievalDriver;

    class DatumStorageDriver;
    class DatumRetrievalDriver;
    class DimTolStorageDriver;
    class DimTolRetrievalDriver;
    class DimTolToolRetrievalDriver;
    class DimTolToolStorageDriver;
    class MaterialStorageDriver;
    class MaterialRetrievalDriver;
    class MaterialToolRetrievalDriver;
    class MaterialToolStorageDriver;

    AddStorageDrivers(aDriverSeq : ASDriverHSequence from MDF; theMsgDriver : MessageDriver from CDM);
	---Purpose: Adds the attribute storage drivers to <aDriverSeq>.


    AddRetrievalDrivers(aDriverSeq : ARDriverHSequence from MDF; theMsgDriver : MessageDriver from CDM);
	---Purpose: Adds the attribute retrieval drivers to <aDriverSeq>.


end MXCAFDoc;
