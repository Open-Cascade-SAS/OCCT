-- File:        CurveOnSurface.cdl
-- Created:     Fri Dec  1 11:11:10 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993



class CurveOnSurface from StepGeom inherits SelectType from StepData

	-- <CurveOnSurface> is an EXPRESS Select Type construct translation.
	-- it gathers : Pcurve, SurfaceCurve, CompositeCurveOnSurface

uses

	Pcurve,
	SurfaceCurve,
	CompositeCurveOnSurface
is

	Create returns CurveOnSurface;
	---Purpose : Returns a CurveOnSurface SelectType

	CaseNum (me; ent : Transient) returns Integer;
	---Purpose: Recognizes a CurveOnSurface Kind Entity that is :
	--        1 -> Pcurve
	--        2 -> SurfaceCurve
	--        3 -> CompositeCurveOnSurface
	--        0 else

	Pcurve (me) returns any Pcurve;
	---Purpose : returns Value as a Pcurve (Null if another type)

	SurfaceCurve (me) returns any SurfaceCurve;
	---Purpose : returns Value as a SurfaceCurve (Null if another type)

	CompositeCurveOnSurface (me) returns any CompositeCurveOnSurface;
	---Purpose : returns Value as a CompositeCurveOnSurface (Null if another type)


end CurveOnSurface;

