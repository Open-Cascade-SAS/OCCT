-- Created on: 1998-02-27
-- Created by: Christian CAILLET
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class ModifEditForm  from IFSelect  inherits Modifier

    ---Purpose : This modifier applies an EditForm on the entities selected

uses CString, AsciiString from TCollection,
     InterfaceModel, CopyTool, Protocol from Interface, ContextModif,
     EditForm

is

    Create (editform : EditForm) returns mutable ModifEditForm;
    ---Purpose : Creates a ModifEditForm. It may not change the graph

    EditForm (me) returns EditForm;
    ---Purpose : Returns the EditForm

    Perform (me; ctx  : in out ContextModif;
    	     target   : mutable InterfaceModel;
    	     protocol : Protocol from Interface;
    	     TC       : in out CopyTool);
    ---Purpose : Acts by applying an EditForm to entities, selected or all model

    Label (me) returns AsciiString from TCollection;
    ---Purpose : Returns Label as "Apply EditForm <+ label of EditForm>"

fields

    theedit : EditForm;

end ModifEditForm;
