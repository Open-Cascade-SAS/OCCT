-- Created on: 2003-06-04
-- Created by: Galina KULIKOVA
-- Copyright (c) 2003-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class GeometricToleranceRelationship from StepDimTol
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity GeometricToleranceRelationship

uses
    HAsciiString from TCollection,
    GeometricTolerance from StepDimTol

is
    Create returns GeometricToleranceRelationship from StepDimTol;
	---Purpose: Empty constructor

    Init (me: mutable; aName: HAsciiString from TCollection;
                       aDescription: HAsciiString from TCollection;
                       aRelatingGeometricTolerance: GeometricTolerance from StepDimTol;
                       aRelatedGeometricTolerance: GeometricTolerance from StepDimTol);
	---Purpose: Initialize all fields (own and inherited)

    Name (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Name
    SetName (me: mutable; Name: HAsciiString from TCollection);
	---Purpose: Set field Name

    Description (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Description
    SetDescription (me: mutable; Description: HAsciiString from TCollection);
	---Purpose: Set field Description

    RelatingGeometricTolerance (me) returns GeometricTolerance from StepDimTol;
	---Purpose: Returns field RelatingGeometricTolerance
    SetRelatingGeometricTolerance (me: mutable; RelatingGeometricTolerance: GeometricTolerance from StepDimTol);
	---Purpose: Set field RelatingGeometricTolerance

    RelatedGeometricTolerance (me) returns GeometricTolerance from StepDimTol;
	---Purpose: Returns field RelatedGeometricTolerance
    SetRelatedGeometricTolerance (me: mutable; RelatedGeometricTolerance: GeometricTolerance from StepDimTol);
	---Purpose: Set field RelatedGeometricTolerance

fields
    theName: HAsciiString from TCollection;
    theDescription: HAsciiString from TCollection;
    theRelatingGeometricTolerance: GeometricTolerance from StepDimTol;
    theRelatedGeometricTolerance: GeometricTolerance from StepDimTol;

end GeometricToleranceRelationship;
