-- Created on: 2007-08-22
-- Created by: Sergey ZARITCHNY
-- Copyright (c) 2007-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class IntPackedMap from PDataStd inherits Attribute from PDF

	---Purpose: Persistance attribute of  TDataStd_IntPackedMap  

uses   
    HArray1OfInteger  from  PColStd


is
    Create returns mutable  IntPackedMap from  PDataStd;

    Init (me : mutable; theLow,  theUp:  Integer  from Standard);
    ---Purpose: Inits the internal container
    --  if  (upper  -  lower)  ==  0  and (upper  |  lower) == 0, the corresponding  
    --  array is empty (not requested)
     
    IsEmpty (me)
    ---Purpose: Returns true if the internal container is empty
    returns Boolean from Standard;  

    Upper  (me)
     ---Purpose: Returns an upper bound of the internal container
    returns Integer from Standard;   

    Lower  (me)
     ---Purpose: Returns a lower bound of the internal container
    returns Integer from Standard;   
    
    GetValue (me; theIndex : Integer from Standard)  
    returns Integer from Standard;
        
    SetValue (me : mutable; theIndex : Integer from Standard;  
    	    	    	    theValue : Integer from Standard);
    
fields 

    myIntValues      :  HArray1OfInteger from PColStd;   
    
end IntPackedMap;
