-- Created on: 2002-12-14
-- Created by: data exchange team
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class DegreeOfFreedom from StepFEA
inherits SelectType from StepData

    ---Purpose: Representation of STEP SELECT type DegreeOfFreedom

uses
    SelectMember from StepData,
    EnumeratedDegreeOfFreedom from StepFEA,
    HAsciiString from TCollection

is
    Create returns DegreeOfFreedom from StepFEA;
	---Purpose: Empty constructor
	
    CaseNum (me; ent: Transient) returns Integer;
	---Purpose: Recognizes a kind of CurveElementFreedom select type
	--          return 0

    CaseMem (me; ent: SelectMember from StepData) returns Integer is redefined;
	---Purpose: Recognizes a items of select member CurveElementFreedomMember
	--          1 -> EnumeratedCurveElementFreedom
	--          2 -> ApplicationDefinedDegreeOfFreedom
	--          0 else
	
    NewMember(me) returns SelectMember from StepData is redefined;
	---Purpose: Returns a new select member the type CurveElementFreedomMember

    SetEnumeratedDegreeOfFreedom (me:in out; aVal: EnumeratedDegreeOfFreedom from StepFEA);
	---Purpose: Returns Value as EnumeratedDegreeOfFreedom (or Null if another type)
	
    EnumeratedDegreeOfFreedom (me) returns EnumeratedDegreeOfFreedom from StepFEA;
    	---Purpose: Returns Value as EnumeratedDegreeOfFreedom (or Null if another type)
	
    SetApplicationDefinedDegreeOfFreedom(me: in out; aVal :HAsciiString from TCollection);
	---Purpose: Set Value for ApplicationDefinedDegreeOfFreedom

    ApplicationDefinedDegreeOfFreedom (me) returns HAsciiString from TCollection;
	---Purpose: Returns Value as ApplicationDefinedDegreeOfFreedom (or Null if another type)

end DegreeOfFreedom;
