-- Created on: 1993-08-16
-- Created by: Bruno DUMORTIER
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class Chronometer from Draw inherits Drawable3D from Draw

	---Purpose: Class to store chronometer variables.

uses

    Timer from OSD,
    Display from Draw,
    Interpretor from Draw

is

    Create returns mutable Chronometer from Draw;
    
    
    Timer(me : mutable) returns Timer from OSD
	---C++: return &
    is static;

    DrawOn(me; dis : in out Display);
	---Purpose: Does nothhing,
    
    Copy(me) returns mutable Drawable3D from Draw
	---Purpose: For variable copy.
    is redefined;
	
    Dump(me; S : in out OStream)
	---Purpose: For variable dump.
    is redefined;

    Whatis(me;  I : in out Interpretor from Draw)
	---Purpose: For variable whatis command.
    is redefined;

fields

    myTimer : Timer from OSD;

end Chronometer;
