-- Created on: 2002-12-12
-- Created by: data exchange team
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class CurveElementIntervalConstant from StepFEA
inherits CurveElementInterval from StepFEA

    ---Purpose: Representation of STEP entity CurveElementIntervalConstant

uses
    CurveElementLocation from StepFEA,
    EulerAngles from StepBasic,
    CurveElementSectionDefinition from StepElement

is
    Create returns CurveElementIntervalConstant from StepFEA;
	---Purpose: Empty constructor

    Init (me: mutable; aCurveElementInterval_FinishPosition: CurveElementLocation from StepFEA;
                       aCurveElementInterval_EuAngles: EulerAngles from StepBasic;
                       aSection: CurveElementSectionDefinition from StepElement);
	---Purpose: Initialize all fields (own and inherited)

    Section (me) returns CurveElementSectionDefinition from StepElement;
	---Purpose: Returns field Section
    SetSection (me: mutable; Section: CurveElementSectionDefinition from StepElement);
	---Purpose: Set field Section

fields
    theSection: CurveElementSectionDefinition from StepElement;

end CurveElementIntervalConstant;
