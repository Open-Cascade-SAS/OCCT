-- File:        PointOnCurve.cdl
-- Created:     Mon Dec  4 12:02:29 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWPointOnCurve from RWStepGeom

	---Purpose : Read & Write Module for PointOnCurve

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     PointOnCurve from StepGeom,
     EntityIterator from Interface

is

	Create returns RWPointOnCurve;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable PointOnCurve from StepGeom);

	WriteStep (me; SW : in out StepWriter; ent : PointOnCurve from StepGeom);

	Share(me; ent : PointOnCurve from StepGeom; iter : in out EntityIterator);

end RWPointOnCurve;
