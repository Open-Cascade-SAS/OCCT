-- Created on: 1993-03-10
-- Created by: JCV
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Plane from Geom inherits ElementarySurface from Geom

        ---Purpose : Describes a plane in 3D space.
    	-- A plane is positioned in space by a coordinate system
    	-- (a gp_Ax3 object) such that the plane is defined by
    	-- the origin, "X Direction" and "Y Direction" of this
    	-- coordinate system.
    	-- This coordinate system is the "local coordinate
    	-- system" of the plane. The following apply:
    	-- - Its "X Direction" and "Y Direction" are respectively
    	--   the u and v parametric directions of the plane.
    	-- - Its origin is the origin of the u and v parameters
    	--   (also called the "origin" of the plane).
    	-- - Its "main Direction" is a vector normal to the plane.
    	--   This normal vector gives the orientation of the
    	--   plane only if the local coordinate system is "direct".
    	--   (The orientation of the plane is always defined by
  	--   the "X Direction" and the "Y Direction" of its local
    	--   coordinate system.)
    	--   The parametric equation of the plane is:
    	-- P(u, v) = O + u*XDir + v*YDir
    	-- where O, XDir and YDir are respectively the
    	-- origin, the "X Direction" and the "Y Direction" of the
    	-- local coordinate system of the plane.
    	-- The parametric range of the two parameters u and v
    	-- is ] -infinity, +infinity [.
        

uses Ax1      from gp,
     Ax3      from gp,
     Dir      from gp,
     Lin      from gp,
     Pln      from gp, 
     Pnt      from gp, 
     Trsf     from gp, 
     Vec      from gp,
     GTrsf2d  from gp,
     Curve    from Geom,
     Geometry from Geom
     
raises ConstructionError from Standard,
       RangeError        from Standard


is



  Create (A3 : Ax3)    returns mutable Plane;
        ---Purpose :
        --  Creates a plane located in 3D space with an axis placement
        --  three axis.  The "ZDirection" of "A3" is the direction normal
        --  to the plane.  The "Location" point of "A3" is the origin of
        --  the plane. The "XDirection" and "YDirection" of "A3" define
        --  the directions of the U isoparametric and V isoparametric
        --  curves.


  Create (Pl : Pln)  returns mutable Plane;
        ---Purpose :
        --  Creates a plane from a non transient plane from package gp.


  Create (P : Pnt; V : Dir)    returns mutable Plane;
        ---Purpose :
        --  P is the "Location" point or origin of the plane.
        --  V is the direction normal to the plane.


  Create (A, B, C ,D : Real)   returns mutable Plane
        ---Purpose :
        --  Creates a plane from its cartesian equation :
        --  Ax + By + Cz + D = 0.0
     raises ConstructionError;
        ---Purpose :
        --  Raised if Sqrt (A*A + B*B + C*C) <= Resolution from gp
  

  SetPln (me : mutable; Pl : Pln);
        ---Purpose :
        --  Set <me> so that <me> has the same geometric properties as Pl.


  Pln (me)  returns Pln
        ---Purpose : Converts this plane into a gp_Pln plane.
         is static;

  
  UReverse (me : mutable)
        ---Purpose : 
        -- Changes the orientation of this plane in the u (or v)
    	-- parametric direction. The bounds of the plane are not
    	-- changed but the given parametric direction is
    	-- reversed. Hence the orientation of the surface is reversed.
  is redefined;

  UReversedParameter (me; U : Real ) returns Real;
	---Purpose: Computes the u  parameter on the modified
    	-- plane, produced when reversing the u 
    	-- parametric of this plane, for any point of u parameter U  on this plane.
    	-- In the case of a plane, these methods return - -U.

  VReverse (me : mutable)
        ---Purpose : 
        -- Changes the orientation of this plane in the u (or v)
    	-- parametric direction. The bounds of the plane are not
    	-- changed but the given parametric direction is
    	-- reversed. Hence the orientation of the surface is reversed.
  is redefined;
  

  VReversedParameter (me; V : Real ) returns Real;
	---Purpose: Computes the v parameter on the modified
    	-- plane, produced when reversing the  v
    	-- parametric of this plane, for any point of v parameter V on this plane.
    	-- In the case of a plane, these methods return -V.
  
  
  TransformParameters(me; U,V : in out Real; T : Trsf from gp)
	---Purpose: Computes the  parameters on the  transformed  surface for
	--          the transform of the point of parameters U,V on <me>.
	--          me->Transformed(T)->Value(U',V')
	--          is the same point as
	--          me->Value(U,V).Transformed(T)
	--          Where U',V' are the new values of U,V after calling
	--          me->TranformParameters(U,V,T)
	--          This methods multiplies U and V by T.ScaleFactor()
     is redefined;  

  ParametricTransformation(me; T : Trsf from gp) returns GTrsf2d from gp
	---Purpose: Returns a 2d transformation  used to find the  new
	--          parameters of a point on the transformed surface.
	--          me->Transformed(T)->Value(U',V')
	--          is the same point as
	--          me->Value(U,V).Transformed(T)
	--          Where U',V' are  obtained by transforming U,V with
	--          th 2d transformation returned by
	--          me->ParametricTransformation(T)
	--          This  methods  returns  a scale  centered  on  the
	--          origin with T.ScaleFactor
     is redefined;  

  Bounds (me; U1, U2, V1, V2 : out Real);
        ---Purpose : Returns the parametric bounds U1, U2, V1 and V2 of this plane.
    	-- Because a plane is an infinite surface, the following is always true:
    	-- - U1 = V1 =   Standard_Real::RealFirst()
    	-- - U2 = V2 =   Standard_Real::RealLast().


  Coefficients (me; A, B, C, D : out Real);
        ---Purpose :
        --  Computes the normalized coefficients of the plane's 
        --  cartesian equation : Ax + By + Cz + D = 0.0


  IsUClosed (me)  returns Boolean;
        ---Purpose : return False


  IsVClosed (me)  returns Boolean;
        ---Purpose : return False


  IsUPeriodic (me)   returns Boolean;
        ---Purpose : return False.


  IsVPeriodic (me)  returns Boolean;
        ---Purpose : return False.


  UIso (me; U : Real)   returns mutable Curve;
        ---Purpose :
        --  Computes the U isoparametric curve.
        --  This is a Line parallel to the YAxis of the plane.


  VIso (me; V : Real)   returns mutable Curve;
        ---Purpose :
        --  Computes the V isoparametric curve.
        --  This is a Line parallel to the XAxis of the plane.


  D0 (me; U, V : Real; P : out Pnt);
        ---Purpose :
        --  Computes the point P (U, V) on <me>.
        --  P = O + U * XDir + V * YDir.
        --  where O is the "Location" point of the plane, XDir the 
        --  "XDirection" and YDir the "YDirection" of the plane's local
        --  coordinate system.


  D1 (me; U, V : Real; P : out Pnt; D1U, D1V : out Vec);
        ---Purpose :
        --  Computes the current point and the first derivatives in the
        --  directions U and V.


  D2 (me; U, V : Real; P : out Pnt; D1U, D1V, D2U, D2V, D2UV : out Vec);
        ---Purpose :
        --  Computes the current point, the first and the second 
        --  derivatives in the directions U and V.


  D3 (me; U, V : Real; P : out Pnt;  
      D1U, D1V, D2U, D2V, D2UV, D3U, D3V, D3UUV, D3UVV :out Vec);
        ---Purpose :
        --  Computes the current point, the first,the second and the 
        --  third derivatives in the directions U and V.


  DN (me; U, V : Real; Nu, Nv : Integer)   returns Vec
        ---Purpose :
        --  Computes the derivative of order Nu in the direction u 
        --  and Nv in the direction v.
     raises RangeError;
        ---Purpose : Raised if Nu + Nv < 1 or Nu < 0 or Nv < 0.



  Transform (me : mutable; T : Trsf);

    	---Purpose: Applies the transformation T to this plane.
        
  Copy (me)  returns mutable like me;

    	---Purpose: Creates a new object which is a copy of this plane.
end;

