-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Shell from StepShape inherits SelectType from StepData

	-- <Shell> is an EXPRESS Select Type construct translation.
	-- it gathers : OpenShell, ClosedShell

uses

	OpenShell,
	ClosedShell
is

	Create returns Shell;
	---Purpose : Returns a Shell SelectType

	CaseNum (me; ent : Transient) returns Integer;
	---Purpose: Recognizes a Shell Kind Entity that is :
	--        1 -> OpenShell
	--        2 -> ClosedShell
	--        0 else

	OpenShell (me) returns any OpenShell;
	---Purpose : returns Value as a OpenShell (Null if another type)

	ClosedShell (me) returns any ClosedShell;
	---Purpose : returns Value as a ClosedShell (Null if another type)


end Shell;

