-- Created on: 2000-01-26
-- Created by: Denis PASCAL
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class ChildNodeIterator from TDataStd 

	---Purpose:  Iterates on the  ChildStepren step of  a step, at the
	--           first level  only.   It  is possible  to ask  the
	--          iterator to explore all the sub step levels of the
	--          given one, with the option "allLevels".

uses TreeNode from TDataStd

is

    Create
    	returns ChildNodeIterator from TDataStd;
    	---Purpose: Creates an empty iterator.
    
    Create(aTreeNode : TreeNode from TDataStd;
    	   allLevels : Boolean from Standard = Standard_False)
    	returns ChildNodeIterator from TDataStd;
    	---Purpose: Iterates on the ChildStepren of the given Step. If
    	--          <allLevels> option is set to true, it explores not
    	--          only the first, but all the sub Step levels.
    
    Initialize(me : in out;
    	       aTreeNode : TreeNode from TDataStd;
    	       allLevels : Boolean from Standard = Standard_False);
    	---Purpose: Initializes the iteration on  the Children Step of
    	--          the  given Step. If <allLevels>  option is  set to
    	--          true, it explores not  only the first, but all the
    	--          sub Step levels.
    
    More(me) returns Boolean;
    	---C++: inline
	---Purpose: Returns True if there is a current Item in the
	--          iteration.
    
    Next(me : in out);
    	---Purpose: Move to the next Item 
    
    NextBrother(me : in out);
    	---Purpose: Move to the next Brother. If there is none, go up
    	--          etc. This method is interesting only with
    	--          "allLevels" behavior, because it avoids to explore
    	--          the current Step ChildStepren.
    
    Value(me) returns TreeNode from TDataStd;
    	---C++: inline
	---Purpose: Returns the current item; a null Step if there is
	--          no one.

fields

    myNode       : TreeNode from TDataStd;
    myFirstLevel : Integer  from Standard;

end ChildNodeIterator;





