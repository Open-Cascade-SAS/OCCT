-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class OrganizationalAddress from StepBasic 

inherits Address from StepBasic 

uses

	HArray1OfOrganization from StepBasic, 
	HAsciiString from TCollection, 
	Organization from StepBasic
is

	Create returns mutable OrganizationalAddress;
	---Purpose: Returns a OrganizationalAddress


	Init (me : mutable;
	      hasAinternalLocation : Boolean from Standard;
	      aInternalLocation : mutable HAsciiString from TCollection;
	      hasAstreetNumber : Boolean from Standard;
	      aStreetNumber : mutable HAsciiString from TCollection;
	      hasAstreet : Boolean from Standard;
	      aStreet : mutable HAsciiString from TCollection;
	      hasApostalBox : Boolean from Standard;
	      aPostalBox : mutable HAsciiString from TCollection;
	      hasAtown : Boolean from Standard;
	      aTown : mutable HAsciiString from TCollection;
	      hasAregion : Boolean from Standard;
	      aRegion : mutable HAsciiString from TCollection;
	      hasApostalCode : Boolean from Standard;
	      aPostalCode : mutable HAsciiString from TCollection;
	      hasAcountry : Boolean from Standard;
	      aCountry : mutable HAsciiString from TCollection;
	      hasAfacsimileNumber : Boolean from Standard;
	      aFacsimileNumber : mutable HAsciiString from TCollection;
	      hasAtelephoneNumber : Boolean from Standard;
	      aTelephoneNumber : mutable HAsciiString from TCollection;
	      hasAelectronicMailAddress : Boolean from Standard;
	      aElectronicMailAddress : mutable HAsciiString from TCollection;
	      hasAtelexNumber : Boolean from Standard;
	      aTelexNumber : mutable HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      hasAinternalLocation : Boolean from Standard;
	      aInternalLocation : mutable HAsciiString from TCollection;
	      hasAstreetNumber : Boolean from Standard;
	      aStreetNumber : mutable HAsciiString from TCollection;
	      hasAstreet : Boolean from Standard;
	      aStreet : mutable HAsciiString from TCollection;
	      hasApostalBox : Boolean from Standard;
	      aPostalBox : mutable HAsciiString from TCollection;
	      hasAtown : Boolean from Standard;
	      aTown : mutable HAsciiString from TCollection;
	      hasAregion : Boolean from Standard;
	      aRegion : mutable HAsciiString from TCollection;
	      hasApostalCode : Boolean from Standard;
	      aPostalCode : mutable HAsciiString from TCollection;
	      hasAcountry : Boolean from Standard;
	      aCountry : mutable HAsciiString from TCollection;
	      hasAfacsimileNumber : Boolean from Standard;
	      aFacsimileNumber : mutable HAsciiString from TCollection;
	      hasAtelephoneNumber : Boolean from Standard;
	      aTelephoneNumber : mutable HAsciiString from TCollection;
	      hasAelectronicMailAddress : Boolean from Standard;
	      aElectronicMailAddress : mutable HAsciiString from TCollection;
	      hasAtelexNumber : Boolean from Standard;
	      aTelexNumber : mutable HAsciiString from TCollection;
	      aOrganizations : mutable HArray1OfOrganization from StepBasic;
	      aDescription : mutable HAsciiString from TCollection) is virtual;

	-- Specific Methods for Field Data Access --

	SetOrganizations(me : mutable; aOrganizations : mutable HArray1OfOrganization);
	Organizations (me) returns mutable HArray1OfOrganization;
	OrganizationsValue (me; num : Integer) returns mutable Organization;
	NbOrganizations (me) returns Integer;
	SetDescription(me : mutable; aDescription : mutable HAsciiString);
	Description (me) returns mutable HAsciiString;

fields

	organizations : HArray1OfOrganization from StepBasic;
	description : HAsciiString from TCollection;

end OrganizationalAddress;
