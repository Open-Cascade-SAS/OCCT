-- Created on: 1997-12-15
-- Created by: Philippe MANGIN
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class  SectionPlacement from  GeomFill

	---Purpose: To place section in sweep Function                   
    	---Level: Advanced

uses 
    LocationLaw  from  GeomFill, 
    Geometry from Geom,
    Curve    from Geom, 
    HCurve   from Adaptor3d, 
    Curve    from GeomAdaptor, 
    ExtPC  from  Extrema,  
    Trsf   from  gp,
    Mat    from  gp, 
    Ax1    from  gp,     
    Vec    from  gp, 
    Pnt    from  gp
     
raises
    NotDone 
    
is
    Create(L  :  LocationLaw  from  GeomFill; 
           Section  :  Geometry  from  Geom)   
    returns   SectionPlacement from  GeomFill; 
     
    SetLocation(me :  in  out;  L  :  LocationLaw  from  GeomFill)  
    ---Purpose: To change the section Law         
    is  static;
	    
    Perform(me:in  out; Tol  :  Real) 
    is  static;    
     
    Perform(me:in  out; Path  :  HCurve  from  Adaptor3d; 
                        Tol  :  Real) 
    is  static;  
     
    Perform(me:in  out; ParamOnPath  :  Real;
                        Tol  :  Real) 
    is  static;   
     
    IsDone(me)   
    returns  Boolean;  
     
    ParameterOnPath(me)  returns  Real; 
     
    ParameterOnSection(me)  returns  Real; 
     
    Distance(me)  returns  Real;  
     
    Angle(me)  returns  Real;
      
    Transformation(me; WithTranslation :  Boolean; 
                   WithCorrection  :  Boolean  =  Standard_False) 
    returns  Trsf  from  gp;
     
    Section(me; WithTranslation  :  Boolean) 
    ---Purpose: Compute the Section, in the coordinate syteme given by
    --          the Location Law.         
    --          If <WithTranslation> contact beetween
    --          <Section> and <Path> is forced.     
    returns  Curve from Geom; 
     
    ModifiedSection(me;  WithTranslation  :  Boolean)  
    ---Purpose: Compute the Section, in the coordinate syteme given by
    --          the Location Law.         
    --          To have the Normal to section equal to the Location
    --          Law Normal.  If <WithTranslation> contact beetween
    --          <Section> and <Path> is forced.
    returns  Curve from Geom; 
     
    SectionAxis(me;  M  :  Mat  from  gp; 
                T,  N,  BN  :  out  Vec  from  gp)  is private; 
		 
    Choix(me;  Dist,  Angle  :  Real)   
    returns  Boolean   
    is  private; 
    
fields
  done    :  Boolean;
  isplan  :  Boolean; 
  TheAxe  :  Ax1  from  gp; 
  Gabarit :  Real;
  myLaw :  LocationLaw  from  GeomFill;
  myAdpSection  :  Curve  from  GeomAdaptor;   
  mySection  :  Curve  from  Geom;  
  SecParam,  PathParam,  Dist,  AngleMax  :  Real; 
  myExt        :  ExtPC  from  Extrema;  
  
  myIsPoint : Boolean from Standard; 
  myPoint   : Pnt     from gp;
  
end ;
