-- Created on: 1996-01-02
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Shell from BRepCheck inherits Result from BRepCheck

	---Purpose: 

uses Shape  from TopoDS,
     Shell  from TopoDS, 
     ListOfShape from TopTools,
     IndexedDataMapOfShapeListOfShape  from  TopTools,
     Status from BRepCheck

is

    Create(S: Shell from TopoDS)
    
    	returns Shell from BRepCheck;


    InContext(me: mutable; ContextShape: Shape from TopoDS);
    


    Minimum(me: mutable);
    

    
    Blind(me: mutable);


    Closed(me: mutable; Update: Boolean from Standard = Standard_False)
	---Purpose: Checks if the oriented  faces of the shell  give a
	--          closed shell.    If the  wire is  closed,  returns
	--          BRepCheck_NoError.If      <Update>     is  set  to
	--          Standard_True, registers the status in the list.
    	returns Status from BRepCheck
	is static;


    Orientation(me: mutable; Update: Boolean from Standard = Standard_False)
	---Purpose: Checks if the   oriented faces  of  the shell  are
	--          correctly oriented.  An internal  call is  made to
	--          the  method  Closed.   If  <Update>    is set   to
	--          Standard_True, registers the status in the list.
    	returns Status from BRepCheck
	is static;


    SetUnorientable(me: mutable)
    
    	is static;


    IsUnorientable(me)
    
    	returns Boolean from Standard
	is static;


    NbConnectedSet (me: mutable; theSets : in out ListOfShape from TopTools)
    
    	returns Integer from Standard;


fields

    myNbori : Integer from Standard;
    myCdone : Boolean from Standard;
    myCstat : Status  from BRepCheck;
    myOdone : Boolean from Standard;
    myOstat : Status  from BRepCheck;
    myMapEF : IndexedDataMapOfShapeListOfShape  from  TopTools;

end Shell;
