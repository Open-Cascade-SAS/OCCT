-- File:        Placement.cdl
-- Created:     Fri Dec  1 11:11:24 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class Placement from StepGeom 

inherits GeometricRepresentationItem from StepGeom 

uses

	CartesianPoint from StepGeom, 
	HAsciiString from TCollection
is

	Create returns mutable Placement;
	---Purpose: Returns a Placement


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aLocation : mutable CartesianPoint from StepGeom) is virtual;

	-- Specific Methods for Field Data Access --

	SetLocation(me : mutable; aLocation : mutable CartesianPoint);
	Location (me) returns mutable CartesianPoint;

fields

	location : CartesianPoint from StepGeom;

end Placement;
