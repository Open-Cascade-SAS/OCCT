-- Created on: 1995-10-24
-- Created by: Mister rmi
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Polygon3D from PPoly inherits Persistent from Standard

    	---Purpose: This class represents a 3d Polygon3D.
    	--          
    	--          It is defined by an array of 3d nodes values.
    	--          If the Polygon3D is closed, the point will be
    	--          repeated.


uses HArray1OfPnt  from PColgp,
     HArray1OfReal from PColStd

is

    Create(Nodes: HArray1OfPnt from PColgp;
    	   Defl : Real from Standard) 
    returns mutable Polygon3D from PPoly;
    	---Purpose: Defaults with allocation of nodes.

    Create(Nodes      : HArray1OfPnt  from PColgp;
           Parameters : HArray1OfReal from PColStd;
    	   Defl       : Real          from Standard) 
    returns mutable Polygon3D from PPoly;
    	---Purpose: Defaults with allocation of nodes + Parameters
    

    Deflection(me) returns Real;

    Deflection(me : mutable; Defl : Real from Standard);
    

    NbNodes(me) returns Integer;
    
    Nodes(me) returns HArray1OfPnt from PColgp;

    Nodes(me : mutable; Nodes : HArray1OfPnt from PColgp);
    

    HasParameters(me) returns Boolean from Standard;

    Parameters(me : mutable; Parameters : HArray1OfReal from PColStd);
    	---Purpose: Sets the value of myParameters

    Parameters(me) returns HArray1OfReal from PColStd;
	---Purpose: Reference on the parameters values.
    
fields

    myDeflection : Real          from Standard;
    myNodes      : HArray1OfPnt  from PColgp;
    myParameters : HArray1OfReal from PColStd;
    	-- myParameters is Optional (Pointer can be Null)
    
end Polygon3D;
