-- File:	BOPTools_CheckResult.cdl
-- Created:	Thu Sep  2 16:18:42 2004
-- Author:	Oleg FEDYAEV
--		<ofv@opencascade.com>
---Copyright:	 Open Cascade 2004

class CheckResult from BOPTools
    ---Purpose: contains information about faulty shapes
    --          and faulty types
uses 
    
    Shape       from TopoDS,
    ListOfShape from TopTools,
    CheckStatus from BOPTools,
    Geometry    from Geom

is

    Create
    	returns CheckResult;
    ---Purpose: empty constructor

    AddShape(me: in out; TheShape: Shape from TopoDS);
    ---Purpose: adds a shape with faulty to a list

    GetShapes(me)
    	returns ListOfShape from TopTools;
    ---C++: return const &
    ---Purpose: gets access to faulty shapes in a list const

    SetCheckStatus(me:in out; TheStatus: CheckStatus from BOPTools);
    ---Purpose: sets faulty status for shapes

    GetCheckStatus(me)
    	returns  CheckStatus from BOPTools;
    ---Purpose: gets faulty status for shapes

    SetInterferenceGeometry(me: in out; TheGeometry: Geometry from Geom);
    ---Purpose: sets an attached geometry to faulty shapes if any

    GetInterferenceGeometry(me)
    	returns Geometry from Geom;
    ---C++: return const &
    ---Purpose: gets an attached geometry to shapes if any

fields

    myStatus   : CheckStatus from BOPTools;
    myShapes   : ListOfShape from TopTools;
    myGeometry : Geometry    from Geom;

end CheckResult;
