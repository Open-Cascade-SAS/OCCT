-- Created on: 1996-01-09
-- Created by: Denis PASCAL
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package DrawDim 

	---Purpose: This package provides Drawable Dimensions. 	
	--          
	--          The classes PlanarDimension and subclasses provide
	--            services  to  build  drawable dimensions between
	--          point line and circle in a given 3d plane.
	--          
	--           The   classes  Dimension and   subclasses provide
	--            services  to build  drawable  dimensions between
	--          plane and cylindrical surfaces.


uses Draw, gp, TColgp, TopoDS, TCollection

is



    deferred class Dimension;
    
    ---Purpose: Dimension between planes and cylinder
    --          =====================================
    
    	class Angle;
	class Distance;
	class Radius;

    
    ---Purpose: Dimensions between point, line and circle ON a plane
    --          ====================================================

    	deferred class PlanarDimension;
	
      	    class PlanarAngle;
      	    class PlanarDistance;
      	    class PlanarRadius; 
    	    class PlanarDiameter;

    ---Purpose: Commands
    --          ========

    DrawShapeName (ashape : Shape from TopoDS; aname : CString);
    
    AllCommands (I : in out Interpretor from Draw);
    
    PlanarDimensionCommands (I : in out Interpretor from Draw);

    ---Purpose: tools
    --          =====

    Nearest (aShape : Shape from TopoDS; apoint : Pnt from gp)
    returns Pnt from gp;

    Lin (e : Edge from TopoDS; l           : in out Lin from gp; 
                               infinite    : in out Boolean from Standard;
                               first, last : in out Real from Standard)
    ---Purpose: false if <e> is not a linear edge
    returns Boolean from Standard;    

    Circ (e : Edge from TopoDS; l : in out Circ from gp; first, last : in out Real from Standard)
    ---Purpose: false if <e> is not a circular edge
    returns Boolean from Standard;

    Pln (f : Face from TopoDS; p : in out Pln from gp)    
    ---Purpose: false if <f> is not a planar face
    returns Boolean from Standard;
    
end DrawDim;



