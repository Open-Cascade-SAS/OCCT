-- Created on: 2001-04-24
-- Created by: Christian CAILLET
-- Copyright (c) 2001-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class MeasureQualification  from StepShape    inherits TShared

    ---Purpose : Added for Dimensional Tolerances

uses
    HAsciiString from TCollection,
    MeasureWithUnit from StepBasic,
    ValueQualifier from StepShape,
    HArray1OfValueQualifier from StepShape

is

    Create returns mutable MeasureQualification;

    Init (me : mutable; name : HAsciiString from TCollection;
    	    description : HAsciiString from TCollection;
	    qualified_measure : MeasureWithUnit from StepBasic;
	    qualifiers : HArray1OfValueQualifier from StepShape);

    Name (me) returns HAsciiString from TCollection;
    SetName (me : mutable; name : HAsciiString from TCollection);

    Description (me) returns HAsciiString from TCollection;
    SetDescription (me : mutable; description : HAsciiString from TCollection);

    QualifiedMeasure (me) returns MeasureWithUnit from StepBasic;
    SetQualifiedMeasure (me : mutable; qualified_measure : MeasureWithUnit from StepBasic);

    Qualifiers (me) returns HArray1OfValueQualifier from StepShape;
    NbQualifiers (me) returns Integer;
    SetQualifiers (me : mutable; qualifiers : HArray1OfValueQualifier from StepShape);
    QualifiersValue (me; num : Integer) returns ValueQualifier from StepShape;
    SetQualifiersValue (me : mutable; num : Integer; aqualifier : ValueQualifier from StepShape);

fields

    theName : HAsciiString from TCollection;
    theDescription : HAsciiString from TCollection;
    theQualifiedMeasure : MeasureWithUnit from StepBasic;
    theQualifiers : HArray1OfValueQualifier from StepShape;

end MeasureQualification;
