-- File:	MDataStd_NamedDataRetrievalDriver.cdl
-- Created:	Wed Jun 27 17:19:10 2007
-- Author:	Sergey ZARITCHNY
--		<szy@friendox>
---Copyright:	Open CASCADE 2007


class NamedDataRetrievalDriver from MDataStd inherits ARDriver from MDF

	---Purpose: 

uses
    RRelocationTable from MDF,
    Attribute        from TDF,
    Attribute        from PDF, 
    MessageDriver    from CDM

is
    Create(theMessageDriver : MessageDriver from CDM)
    returns mutable NamedDataRetrievalDriver from MDataStd;

    VersionNumber(me) returns Integer from Standard;

    SourceType(me) returns Type from Standard;

    NewEmpty (me) returns mutable Attribute from TDF;

    Paste(me;
    	  Source     :         Attribute from PDF;
    	  Target     : mutable Attribute from TDF;
    	  RelocTable : RRelocationTable from MDF);

end NamedDataRetrievalDriver;
