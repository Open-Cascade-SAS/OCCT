-- Created on: 1994-11-03
-- Created by: Marie Jose MARTZ
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class Actor from IGESToBRep
    inherits ActorOfTransientProcess  from Transfer

    ---Purpose : This class performs the transfer of an Entity from
    --           IGESToBRep
    --           
    --           I.E. for each type of Entity, it invokes the appropriate Tool
    --           then returns the Binder which contains the Result

uses TransientProcess, Binder, InterfaceModel from Interface

is

    Create  returns mutable Actor from IGESToBRep;

    SetModel (me : mutable; model : InterfaceModel from Interface);
    
    SetContinuity (me : mutable; continuity : Integer from Standard = 0);
    ---Purpose   By default continuity = 0
    --           if continuity = 1 : try C1
    --           if continuity = 2 : try C2
    
    GetContinuity (me) returns Integer from Standard;
    ---Purpose : Return "thecontinuity"

    Recognize (me : mutable; start : Transient) returns Boolean  is redefined;

    Transfer (me : mutable; start : Transient; TP : mutable TransientProcess)
    	returns mutable Binder  is redefined;

    UsedTolerance (me) returns Real;
    ---Purpose : Returns the tolerance which was actually used, either from
    --           the file or from statics

fields

    themodel      : InterfaceModel from Interface;
    thecontinuity : Integer;
    theeps        : Real;

end Actor;
