-- Created on: 1997-08-07
-- Created by: VAUTHIER Jean-Claude
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- modified     Sergey Zaritchny


class PlacementRetrievalDriver from MDataXtd  inherits ARDriver from MDF

	---Purpose: 

uses RRelocationTable from MDF,
     Attribute        from PDF,
     Attribute        from TDF, 
     MessageDriver    from CDM

is


    Create(theMessageDriver : MessageDriver from CDM)  -- Version 0
    returns mutable PlacementRetrievalDriver from MDataXtd;
    

    VersionNumber(me) returns Integer from Standard;
	---Purpose: Returns the version number from which the driver
	--          is available: 0.

    SourceType(me) returns Type from Standard;
	---Purpose: Returns the type: Placement from PDataXtd.

    NewEmpty (me)  returns mutable Attribute from TDF;


    Paste(me;
    	  Source     :         Attribute from PDF;
    	  Target     : mutable Attribute from TDF;
    	  RelocTable : RRelocationTable  from MDF);

end PlacementRetrievalDriver;
