-- Created on: 1991-10-10
-- Created by: Jean Claude VAUTHIER
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.





class CylinderToBSplineSurface  from Convert

        --- Purpose :
        --  This algorithm converts a bounded cylinder into a rational 
        --  B-spline surface. The cylinder is a Cylinder from package gp. 
        --  The parametrization of the cylinder is  :
        --  P (U, V) = Loc + V * Zdir + Radius * (Xdir*Cos(U) + Ydir*Sin(U)) 
        --  where Loc is the location point of the cylinder, Xdir, Ydir and
        --  Zdir are the normalized directions of the local cartesian
        --  coordinate system of the cylinder (Zdir is the direction of the
        --  cylinder's axis). The U parametrization range is U [0, 2PI].
        --- KeyWords :
        --  Convert, Cylinder, BSplineSurface.

inherits ElementarySurfaceToBSplineSurface


uses Cylinder from gp

raises DomainError from Standard

is

  Create (Cyl : Cylinder; U1, U2, V1, V2 : Real)
     returns CylinderToBSplineSurface
       --- Purpose : 
       --  The equivalent B-splineSurface as the same orientation as the 
       --  cylinder in the U and V parametric directions.
     raises DomainError;
        --- Purpose :
        --  Raised if U1 = U2 or U1 = U2 + 2.0 * Pi
        --  Raised if V1 = V2.


  Create (Cyl : Cylinder; V1, V2 : Real)
     returns CylinderToBSplineSurface
       --- Purpose : 
       --  The equivalent B-splineSurface as the same orientation as the
       --  cylinder in the U and V parametric directions.
     raises DomainError;
        --- Purpose :
        --  Raised if V1 = V2.


end CylinderToBSplineSurface;


