-- Created on: 1996-01-08
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



deferred class ProjectedWires from LocOpe inherits TShared from MMgt

	---Purpose: 

uses Face   from TopoDS,
     Wire   from TopoDS,
     Edge   from TopoDS,
     Vertex from TopoDS

is

    InitEdgeIterator(me: mutable)
    
    	is deferred;


    MoreEdge(me: mutable)
    	returns Boolean from Standard
	is deferred;


    Edge(me: mutable)
    	returns Edge from TopoDS
	is deferred;


    OnFace(me: mutable)
	---Purpose: Returns the face of the shape on which the current
	--          edge is projected.
    	returns Face from TopoDS
	is deferred;

    
    OnEdge(me: mutable; E: out Edge from TopoDS)
	---Purpose: If the   current  edge is  projected  on  an edge,
	--          returns <Standard_True> and sets the value of <E>.
	--          Otherwise, returns <Standard_False>.
    	returns Boolean from Standard
	is deferred;


    NextEdge(me: mutable)
    
    	is deferred;


    OnVertex(me: mutable; Vwire :     Vertex from TopoDS;
    	                  Vshape: out Vertex from TopoDS)
			  
	returns Boolean from Standard
	is deferred;


    OnEdge(me: mutable; V: Vertex from TopoDS;
                        E: out Edge from TopoDS;
			P: out Real from Standard)
	---Purpose: If the vertex <V> lies on  an edge of the original
	--          shape,  returns     <Standard_True> and   sets the
	--          concerned edge in  <E>,  and the parameter on  the
	--          edge in <P>.
	--          Else returns <Standard_False>.
	returns Boolean from Standard
	is deferred;


end ProjectedWires;
