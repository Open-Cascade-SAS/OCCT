-- Created on: 2002-10-29
-- Created by: Michael SAZONOV
-- Copyright (c) 2002-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



package BinDrivers

uses
    Standard,
    TDF,
    TCollection,
    TColStd,
    CDM,
    PCDM,
    Storage,
    BinObjMgt,
    BinMDF,
    BinLDrivers

is

    class DocumentStorageDriver;
    class DocumentRetrievalDriver;

    Factory (theGUID : GUID from Standard) returns Transient from Standard;

    AttributeDrivers (MsgDrv : MessageDriver from CDM)
    	returns ADriverTable from BinMDF;
    	---Purpose: Creates the table of drivers of types supported

    StorageVersion returns AsciiString from TCollection;
        ---Purpose: returns "1"
    
end BinDrivers;
