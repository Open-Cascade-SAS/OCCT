-- Created on: 1994-02-17
-- Created by: Bruno DUMORTIER
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.





class Profiler from GeomFill

	---Purpose: Evaluation of the common BSplineProfile of a group
	--          of curves  from Geom. All the curves will have the
	--          same  degree,  the same knot-vector, so  the  same
	--          number of poles.


uses
    Array1OfReal    from TColStd,
    Array1OfInteger from TColStd,
    Array1OfPnt     from TColgp,
    Curve           from Geom,
    SequenceOfCurve from TColGeom


raises
    NotDone     from StdFail,
    DomainError from Standard

is
    Create returns Profiler from GeomFill;
    
    Delete(me:out) is virtual;
    ---C++: alias "Standard_EXPORT virtual ~GeomFill_Profiler(){Delete() ; }"
    
    AddCurve( me    : in out;
              Curve : in Curve from Geom)
    is static;
    
    Perform(me   : in out ;
            PTol : in Real from Standard)
	---Purpose: Converts all curves to BSplineCurves.
	--          Set them to the common profile.
	--          <PTol> is used to compare 2 knots.
    is virtual;
    
    Degree(me) returns Integer from Standard
    raises 
    	NotDone from StdFail
	---Purpose: Raises if not yet perform
    is static;
    
    IsPeriodic(me) returns Boolean from Standard
	---C++: inline
    is static;
    
    NbPoles(me) returns Integer from Standard
    raises 
    	NotDone from StdFail
	---Purpose: Raises if not yet perform
    is static;
    
    Poles(me; Index : in     Integer     from Standard;
    	      Poles : in out Array1OfPnt from TColgp)
    	---Purpose: returns in <Poles> the  poles  of the BSplineCurve
    	--          from index <Index> adjusting to the current profile.
    raises 
    	NotDone     from StdFail,
	---Purpose: Raises if not yet perform
    	DomainError from Standard
	---Purpose: Raises if <Index> not in the range [1,NbCurves]
	--          if  the  length  of  <Poles>  is  not  equal  to
	--          NbPoles().
    is static;
    
    Weights(me; Index   : in     Integer      from Standard;
    	        Weights : in out Array1OfReal from TColStd)
    	---Purpose: returns in <Weights> the weights of the BSplineCurve
    	--          from index <Index> adjusting to the current profile.
    raises 
    	NotDone from StdFail,
	---Purpose: Raises if not yet perform
    	DomainError from Standard
	---Purpose: Raises if <Index> not in the range [1,NbCurves] or
	--          if  the  length  of  <Weights>  is  not  equal  to
	--          NbPoles().
    is static;
    
    NbKnots(me) returns Integer from Standard
    raises 
    	NotDone from StdFail
	---Purpose: Raises if not yet perform
    is static;
    
    KnotsAndMults(me;
                  Knots : in out Array1OfReal    from TColStd;
		  Mults : in out Array1OfInteger from TColStd)
    raises 
    	NotDone from StdFail,
	---Purpose: Raises if not yet perform
    	DomainError from Standard
	---Purpose: Raises if  the lengthes of <Knots> and <Mults> are
	--          not equal to NbKnots().
    is static;
    
    Curve(me; Index : Integer from Standard) 
    returns Curve from Geom
    	---C++: return const&
    	---C++: inline
    is static;
    
    
fields
    mySequence   : SequenceOfCurve from TColGeom is protected;
    myIsDone     : Boolean         from Standard is protected;
    myIsPeriodic : Boolean         from Standard is protected;

end Profiler;
