-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class UniformCurveAndRationalBSplineCurve from StepGeom 

inherits BSplineCurve from StepGeom 


	--- This classe is an implementation of EXPRESS
	--  ANDOR Subtype Declaration.
uses

	UniformCurve from StepGeom, 
	RationalBSplineCurve from StepGeom, 
	HAsciiString from TCollection, 
	Integer from Standard, 
	HArray1OfCartesianPoint from StepGeom, 
	BSplineCurveForm from StepGeom, 
	Logical from StepData, 
	HArray1OfReal from TColStd, 
	Real from Standard
is

	Create returns mutable UniformCurveAndRationalBSplineCurve;
	---Purpose: Returns a UniformCurveAndRationalBSplineCurve


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aDegree : Integer from Standard;
	      aControlPointsList : mutable HArray1OfCartesianPoint from StepGeom;
	      aCurveForm : BSplineCurveForm from StepGeom;
	      aClosedCurve : Logical from StepData;
	      aSelfIntersect : Logical from StepData) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aDegree : Integer from Standard;
	      aControlPointsList : mutable HArray1OfCartesianPoint from StepGeom;
	      aCurveForm : BSplineCurveForm from StepGeom;
	      aClosedCurve : Logical from StepData;
	      aSelfIntersect : Logical from StepData;
	      aUniformCurve : mutable UniformCurve from StepGeom;
	      aRationalBSplineCurve : mutable RationalBSplineCurve from StepGeom) is virtual;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aDegree : Integer from Standard;
	      aControlPointsList : mutable HArray1OfCartesianPoint from StepGeom;
	      aCurveForm : BSplineCurveForm from StepGeom;
	      aClosedCurve : Logical from StepData;
	      aSelfIntersect : Logical from StepData;
	      aWeightsData : mutable HArray1OfReal from TColStd) is virtual;

	-- Specific Methods for Field Data Access --

	SetUniformCurve(me : mutable; aUniformCurve : mutable UniformCurve);
	UniformCurve (me) returns mutable UniformCurve;
	SetRationalBSplineCurve(me : mutable; aRationalBSplineCurve : mutable RationalBSplineCurve);
	RationalBSplineCurve (me) returns mutable RationalBSplineCurve;

	-- Specific Methods for ANDOR Field Data Access --

	SetWeightsData(me : mutable; aWeightsData : mutable HArray1OfReal);
	WeightsData (me) returns mutable HArray1OfReal;
	WeightsDataValue (me; num : Integer) returns Real;
	NbWeightsData (me) returns Integer;

	-- Specific Methods for ANDOR Field Data Access --


fields

	uniformCurve : UniformCurve from StepGeom;
	rationalBSplineCurve : RationalBSplineCurve from StepGeom;

end UniformCurveAndRationalBSplineCurve;
