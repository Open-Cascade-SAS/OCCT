-- File:	TopoDSToStep_Builder.cdl
-- Created:	Fri Nov 25 08:31:25 1994
-- Author:	Frederic MAUPAS
--		<fma@stylox>
---Copyright:	 Matra Datavision 1994


class Builder from TopoDSToStep
    inherits Root from TopoDSToStep

    ---Purpose: This builder Class provides services to build
    --          a ProSTEP Shape model from a Cas.Cad BRep.                 

uses

    FinderProcess                 from Transfer,
    Shape                         from TopoDS,
    Tool                          from TopoDSToStep,
    BuilderError                  from TopoDSToStep,
    TopologicalRepresentationItem from StepShape

raises NotDone from StdFail 
    
is 

--  -----------------------------------------------------------
--  Constructor
--  -----------------------------------------------------------

    Create returns Builder from TopoDSToStep;
    
    Create(S           : Shape from TopoDS;
           T           : in out Tool from TopoDSToStep;
           FP          : mutable FinderProcess from Transfer)
    	returns Builder from TopoDSToStep;
    
    Init(me          : in out;
         S           : Shape from TopoDS;
         T           : in out Tool from TopoDSToStep;
         FP          : mutable FinderProcess from Transfer);
    
--  -----------------------------------------------------------    
--  Get the Result
--  -----------------------------------------------------------

    Error(me) returns BuilderError from TopoDSToStep;
    
    Value (me) returns TopologicalRepresentationItem from StepShape
    	raises NotDone
    	is static;
    	---C++: return const &

fields

    myResult : TopologicalRepresentationItem from StepShape;
    
    myError  : BuilderError                  from TopoDSToStep;

end Builder;
