-- Created on: 1996-12-16
-- Created by: Remi Lequette
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Builder from TNaming  

	---Purpose: A tool to create and maintain topological attributes. 
    	-- Constructor creates an empty
    	-- TNaming_NamedShape attribute at the given
    	-- label. It allows adding "old shape" and "new
    	-- shape" pairs with the specified evolution to this
    	-- named shape. One evolution type per one
    	-- builder must be used.
        
uses
    Shape                        from TopoDS,
    Label                        from TDF,
    Data                         from TDF, 
    NamedShape                   from TNaming,	
    UsedShapes                   from TNaming
    
raises
    ConstructionError            from Standard
is

	Create (aLabel : Label from TDF) returns Builder from TNaming;
	    ---Purpose:  Create an   Builder.   
	    --  Warning:  Before Addition copies the current Value, and clear 
    	

	---Category: To Load Shape Evolution
	--           =======================
      
    	Generated(me : in out; newShape : Shape from TopoDS);
	    ---Purpose:  Records the shape newShape which was
    	    -- generated during a topological construction.
    	    --  As an example, consider the case of a face
    	    --  generated in construction of a box.
	    
	Generated(me : in out; oldShape, newShape : Shape from TopoDS);
	    ---Purpose: Records the shape newShape which was
    	    --  generated from the shape oldShape during a topological construction.
    	    -- As an example, consider the case of a face
    	    -- generated from an edge in construction of a prism.
    

	---Category: Load Modifications.

	Delete(me : in out; oldShape : Shape from TopoDS);
	    ---Purpose:  Records the shape oldShape which was deleted from the current label.
    	    -- As an example, consider the case of a face removed by a Boolean operation.
	    
	Modify(me : in out; oldShape, newShape : Shape from TopoDS);
	    ---Purpose:  Records the shape newShape which is a
    	    -- modification of the shape oldShape.
    	    -- As an example, consider the case of a face split
    	    --  or merged in a Boolean operation.
	    --          
	
    	---Category: Load Selection.
    	Select (me : in out; aShape, inShape : Shape from TopoDS);
	    ---Purpose:   Add a  Shape to the current label ,  This Shape is
	    --          unmodified.  Used for example  to define a set
	    --          of shapes under a label.
			      

        ---Category: Querying

    	NamedShape(me) returns NamedShape from TNaming;
	    ---Purpose: Returns the NamedShape which has been built or is under construction.  

fields

    myShapes: UsedShapes from TNaming; 
    myAtt   : NamedShape from TNaming;
end Builder;
