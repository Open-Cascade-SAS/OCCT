-- Created on: 1993-01-09
-- Created by: CKY / Contract Toubro-Larsen ( Anand NATRAJAN )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class ExternalRefLibName from IGESBasic  inherits IGESEntity

        ---Purpose: defines ExternalRefLibName, Type <416> Form <4>
        --          in package IGESBasic
        --          Used when it is assumed that a copy of the subfigure
        --          exists in native form in a library on the receiving 
        --          system

uses

        HAsciiString from TCollection

is

        Create returns mutable ExternalRefLibName;

        -- Specific Methods pertaining to the class

        Init (me : mutable; aLibName, anExtName : HAsciiString);
        ---Purpose : This method is used to set the fields of the class
        --           ExternalRefLibName
        --       - aLibName  : Name of library in which ExtName resides
        --       - anExtName : External Reference Entity Symbolic Name

        LibraryName (me) returns HAsciiString from TCollection;
        ---Purpose : returns name of library in which External Reference Entity
        -- Symbolic Name resides

        ReferenceName (me) returns HAsciiString from TCollection;
        ---Purpose : returns External Reference Entity Symbolic Name

fields

--
-- Class    : IGESBasic_ExternalRefLibName
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class ExternalRefLibName.
--
-- Reminder : A ExternalRefLibName instance is defined by :
--            - Name of library in which name resides
--            - External Reference Entity Symbolic Name

        theLibName              : HAsciiString from TCollection;
        theExtRefEntitySymbName : HAsciiString from TCollection;

end ExternalRefLibName;
