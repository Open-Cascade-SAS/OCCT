-- Created on: 1999-03-09
-- Created by: Roman LYGIN
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



private class TrsfModification from ShapeCustom inherits TrsfModification from BRepTools

	---Purpose: Complements BRepTools_TrsfModification to provide reversible
	--          scaling regarding tolerances.
	--          Uses actual tolerances (attached to the shapes) not ones
	--          returned by BRep_Tool::Tolerance to work with tolerances
    	--          lower than Precision::Confusion.

uses
    Face     from TopoDS,
    Edge     from TopoDS,
    Vertex   from TopoDS,
    Location from TopLoc,
    Shape    from GeomAbs,
     
    Surface  from Geom,
    Curve    from Geom,
    Curve    from Geom2d,
     
    Trsf     from gp,
    Pnt      from gp

is
    Create (T: Trsf from gp) returns mutable TrsfModification from ShapeCustom;
    	---Purpose: Empty constructor
    
    NewSurface (me: mutable; F       :     Face     from TopoDS;
                             S       : out Surface  from Geom;
		             L       : out Location from TopLoc;
		             Tol     : out Real     from Standard;
                             RevWires: out Boolean from Standard;
                             RevFace : out Boolean from Standard)
    returns Boolean from Standard;
      	---Purpose: Calls inherited method.
	--          Sets <Tol> as actual tolerance of <F> multiplied with scale
	--          factor.

    NewCurve (me: mutable; E  :     Edge     from TopoDS;
                           C  : out Curve    from Geom;
		           L  : out Location from TopLoc;
		           Tol: out Real     from Standard)
    returns Boolean from Standard;
      	---Purpose: Calls inherited method.
	--          Sets <Tol> as actual tolerance of <E> multiplied with scale
	--          factor.

    NewPoint (me: mutable; V  :     Vertex   from TopoDS;
                           P  : out Pnt      from gp;
		           Tol: out Real     from Standard)
    returns Boolean from Standard;
      	---Purpose: Calls inherited method.
	--          Sets <Tol> as actual tolerance of <V> multiplied with scale
	--          factor.

    NewCurve2d (me: mutable;  E    :     Edge     from TopoDS;
                              F    :     Face     from TopoDS;
                              NewE :     Edge     from TopoDS;
                              NewF :     Face     from TopoDS;
                              C    : out Curve    from Geom2d;
		              Tol  : out Real     from Standard)
    returns Boolean from Standard;
      	---Purpose: Calls inherited method.
	--          Sets <Tol> as actual tolerance of <E> multiplied with scale
	--          factor.

    NewParameter (me: mutable; V  :     Vertex   from TopoDS;
                               E  :     Edge     from TopoDS;
                               P  : out Real     from Standard;
  		               Tol: out Real     from Standard)
    returns Boolean from Standard;
      	---Purpose: Calls inherited method.
	--          Sets <Tol> as actual tolerance of <V> multiplied with scale
	--          factor.

end TrsfModification;
