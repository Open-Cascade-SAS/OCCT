-- File:        FillAreaStyleColour.cdl
-- Created:     Mon Dec  4 12:02:27 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWFillAreaStyleColour from RWStepVisual

	---Purpose : Read & Write Module for FillAreaStyleColour

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     FillAreaStyleColour from StepVisual,
     EntityIterator from Interface

is

	Create returns RWFillAreaStyleColour;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable FillAreaStyleColour from StepVisual);

	WriteStep (me; SW : in out StepWriter; ent : FillAreaStyleColour from StepVisual);

	Share(me; ent : FillAreaStyleColour from StepVisual; iter : in out EntityIterator);

end RWFillAreaStyleColour;
