-- Created on: 1993-09-01
-- Created by: Laurent PAINNOT
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class FunctionTool from AppCont


uses Function        from AppCont,
     Pnt             from gp,
     Pnt2d           from gp,
     Vec             from gp,
     Vec2d           from gp,
     Array1OfPnt     from TColgp,
     Array1OfPnt2d   from TColgp,
     Array1OfVec     from TColgp,
     Array1OfVec2d   from TColgp

is
    
    FirstParameter(myclass; C: Function from AppCont) returns Real;
    	---Purpose: returns the first parameter of the Function.

    LastParameter(myclass; C: Function from AppCont) returns Real;
    	---Purpose: returns the last parameter of the Function.

    NbP2d(myclass; C: Function from AppCont) returns Integer;
    	---Purpose: Returns 0.


    NbP3d(myclass; C: Function from AppCont) returns Integer;
    	---Purpose: Returns 1. (the approximation will be done only for one 
    	--          function.


    Value(myclass; C: Function from AppCont; U: Real; tabPt: out Array1OfPnt);
    	---Purpose: <tabP> is an array of only 1 element, the point value at
    	--          the parameter <U>.


    D1(myclass; C: Function from AppCont; U: Real; tabV: out Array1OfVec)
    returns Boolean;
    	---Purpose: <tabV> is an array of only 1 element, the derivative 
    	--          value at the parameter <U>.


    ----------------------------------------------------------
    -- the following methods won t be called by the algorithms
    -- but the description must exist in the tool.
    ----------------------------------------------------------



    Value(myclass; C: Function from AppCont;U: Real; 
    	  tabPt2d: out Array1OfPnt2d);
    
    Value(myclass; C: Function from AppCont; U: Real; 
    	  tabPt: out Array1OfPnt;
    	  tabPt2d: out Array1OfPnt2d);


    D1(myclass;C: Function from AppCont;U: Real; 
    	     tabV2d: out Array1OfVec2d)
    returns Boolean;


    D1(myclass; C: Function from AppCont; U: Real; 
    	     tabV: out Array1OfVec;
	     tabV2d: out Array1OfVec2d)
    returns Boolean;


end FunctionTool;    
    
