-- File:	IGESBasic_ToolOrderedGroupWithoutBackP.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolOrderedGroupWithoutBackP  from IGESBasic

    ---Purpose : Tool to work on a OrderedGroupWithoutBackP. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses OrderedGroupWithoutBackP from IGESBasic,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolOrderedGroupWithoutBackP;
    ---Purpose : Returns a ToolOrderedGroupWithoutBackP, ready to work


    ReadOwnParams (me; ent : mutable OrderedGroupWithoutBackP;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : OrderedGroupWithoutBackP;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : OrderedGroupWithoutBackP;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a OrderedGroupWithoutBackP <ent>, from
    --           its specific (own) parameters

    OwnCorrect (me; ent : mutable OrderedGroupWithoutBackP) returns Boolean  is static;
    ---Purpose : Sets automatic unambiguous Correction on an OrderedGroupWithoutBackP
    --           (Null Elements are removed from list)

    DirChecker (me; ent : OrderedGroupWithoutBackP) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : OrderedGroupWithoutBackP;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : OrderedGroupWithoutBackP; entto : mutable OrderedGroupWithoutBackP;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : OrderedGroupWithoutBackP;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolOrderedGroupWithoutBackP;
