-- Created on: 1992-03-26
-- Created by: Herve LEGRAND
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package GeomLProp

    ---Purpose: These global functions compute the degree of
    --          continuity of a 3D curve built by concatenation of two
    --          other curves (or portions of curves) at their junction point.

uses Standard, gp, Geom, GeomAbs, LProp

is
    
    private  class CurveTool; 
    private  class SurfaceTool;
					    
    class CLProps from GeomLProp 
            instantiates CLProps from LProp(Curve      from Geom,
	                                    Vec        from gp,
					    Pnt        from gp,
					    Dir        from gp,
					    CurveTool  from GeomLProp); 
					     

    class SLProps from GeomLProp 
            instantiates SLProps from LProp(Surface     from Geom,
	                                    SurfaceTool from GeomLProp); 

    
    Continuity(C1,C2 : Curve from Geom;
    	       u1,u2 : Real from Standard;
    	       r1,r2 : Boolean from Standard;
               tl,ta : Real from Standard) 
    ---Purpose: Computes the regularity at the junction between C1 and
    --          C2. The booleans r1 and r2 are true if the curves must
    --          be taken reversed.  The point u1 on C1 and the point
    --          u2 on C2 must be confused.
    --          tl and ta are the linear and angular tolerance used two
    --          compare the derivative.
    returns Shape from GeomAbs;

    
    Continuity(C1,C2 : Curve from Geom;
    	       u1,u2 : Real from Standard;
    	       r1,r2 : Boolean from Standard) 
    ---Purpose: The  same  as  preciding   but   using  the   standard
    --          tolerances from package Precision.
    returns Shape from GeomAbs;

end GeomLProp;    




