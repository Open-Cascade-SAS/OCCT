-- Created on: 1996-12-17
-- Created by: Yves FRICAUD
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

private class RefShape from TNaming 

uses
   Label       from TDF,
   NamedShape  from TNaming, 	
   Shape       from TopoDS,
   PtrNode     from TNaming     

is
    Create returns RefShape from TNaming;
	---C++: inline    
    
    Create (S : Shape from TopoDS) returns RefShape from TNaming;
	---C++: inline    
    
    Shape    (me : in out; S    : Shape    from TopoDS);
    	---C++: inline
    
    FirstUse (me : in out; aPtr : PtrNode from TNaming);
	---C++: inline

    ---Category: Querying

    FirstUse (me) returns PtrNode from TNaming;
	---C++: inline    
    
    Shape (me) returns Shape    from TopoDS;
	---C++: return const&
    	---C++: inline

    Label (me) returns Label from TDF;
    
    NamedShape (me) returns NamedShape from TNaming;

	    
fields

    myShape      : Shape    from TopoDS;
    myFirstUse   : PtrNode  from TNaming;	

end RefShape;
