-- File:	MDataStd_IntPackedMapRetrievalDriver.cdl
-- Created:	Thu Aug 23 10:20:22 2007
-- Author:	Sergey ZARITCHNY
--		<sergey.zaritchny@opencascade.com>
---Copyright:	Open CasCade SA 2007


class IntPackedMapRetrievalDriver from MDataStd inherits ARDriver from MDF

	---Purpose: Retrieval driver of IntPackedMap attribute

uses
    RRelocationTable from MDF,
    Attribute        from PDF,
    Attribute        from TDF, 
    MessageDriver    from CDM 

is
    Create(theMessageDriver : MessageDriver from CDM)  -- Version 0
    returns mutable IntPackedMapRetrievalDriver from MDataStd;
    

    VersionNumber(me) returns Integer from Standard;
	---Purpose: Returns the version number from which the driver
	--          is available: 0.

    SourceType(me) returns Type from Standard;
	---Purpose: Returns the type: IntPackedMap from PDataStd.

    NewEmpty (me)  returns mutable Attribute from TDF;


    Paste(me;
    	  Source     :         Attribute from PDF;
    	  Target     : mutable Attribute from TDF;
    	  RelocTable : RRelocationTable  from MDF);

end IntPackedMapRetrievalDriver;
