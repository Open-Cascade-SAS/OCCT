-- Created on: 1994-05-31
-- Created by: Modelistation
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class IGESTypeForm from IGESSelect    inherits Signature  from IFSelect

    ---Purpose : IGESTypeForm is a Signature specific to the IGES Norm :
    --           it gives the signature under two possible forms :
    --           - as "mmm nnn", with "mmm" as IGES Type Number, and "nnn"
    --             as IGES From Number (even if = 0)  [Default]
    --           - as "mmm" alone, which gives only the IGES Type Number

uses CString, Transient, InterfaceModel

is

    Create (withform : Boolean = Standard_True) returns mutable IGESTypeForm;
    ---Purpose : Creates a Signature for IGES Type & Form Numbers
    --           If <withform> is False, for IGES Type Number only

    SetForm (me : mutable; withform : Boolean);
    ---Purpose : Changes the mode for giving the Form Number

    Value (me; ent : any Transient; model : InterfaceModel) returns CString;
    ---Purpose : Returns the signature for IGES, "mmm nnn" or "mmm" according
    --           creation choice (Type & Form or Type only)

fields

    theform : Boolean;

end IGESTypeForm;
