-- File:        LayeredItem.cdl
-- Created:     Fri Dec  1 11:11:11 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993



class LayeredItem from StepVisual inherits SelectType from StepData

	-- <LayeredItem> is an EXPRESS Select Type construct translation.
	-- it gathers : PresentationRepresentation, RepresentationItem

uses

	PresentationRepresentation,
	RepresentationItem from StepRepr
is

	Create returns LayeredItem;
	---Purpose : Returns a LayeredItem SelectType

	CaseNum (me; ent : Transient) returns Integer;
	---Purpose: Recognizes a LayeredItem Kind Entity that is :
	--        1 -> PresentationRepresentation
	--        2 -> RepresentationItem
	--        0 else

	PresentationRepresentation (me) returns any PresentationRepresentation;
	---Purpose : returns Value as a PresentationRepresentation (Null if another type)

	RepresentationItem (me) returns any RepresentationItem;
	---Purpose : returns Value as a RepresentationItem (Null if another type)


end LayeredItem;

