-- Created on: 1994-05-31
-- Created by: Christian CAILLET
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SelectVisibleStatus  from IGESSelect  inherits SelectExtract

    ---Purpose : This selection looks at Blank Status of IGES Entities
    --           Direct  selection keeps Visible Entities (Blank = 0),
    --           Reverse selection keeps Blanked Entities (Blank = 1)


uses AsciiString from TCollection, Transient, InterfaceModel

is

    Create returns mutable SelectVisibleStatus;
    ---Purpose : Creates a SelectVisibleStatus

    Sort (me; rank : Integer; ent : Transient; model : InterfaceModel)
    	returns Boolean;
    ---Purpose : Returns True if <ent> is an IGES Entity with Blank Status = 0

    ExtractLabel (me) returns AsciiString from TCollection;
    ---Purpose : Returns the Selection criterium : "IGES Entity, Status Visible"

end SelectVisibleStatus;
