-- Created on: 1998-11-13
-- Created by: Jean-Michel BOULCOURT
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package BRepProj

        ---Purpose:     The BRepProj    package  provides   Projection
        --            Algorithms     like  Cylindrical    and  Conical
        --          Projections.  Those algorithms have been put in an
        --          independant package   instead of  BRepAlgo   (like
        --          NormalProjection) because of cyclic reference with
        --          BRepFill. So this package is not available for
        --          the moment to BRepFill.
        --          

uses
    gp, 
    TopoDS,     
    TopTools
	      
is

    
    class  Projection; 
        ---Purpose: provides  conical  and  cylindrical projections of  
        --          Edge  or Wire  on  a Shape from TopoDS. The result  
        --          will be a Edge  or  Wire  from  TopoDS.    
	

end BRepProj;
