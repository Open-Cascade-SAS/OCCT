-- File:	RWStepFEA_RWCurveElementLocation.cdl
-- Created:	Thu Dec 12 17:51:04 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWCurveElementLocation from RWStepFEA

    ---Purpose: Read & Write tool for CurveElementLocation

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    CurveElementLocation from StepFEA

is
    Create returns RWCurveElementLocation from RWStepFEA;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : CurveElementLocation from StepFEA);
	---Purpose: Reads CurveElementLocation

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: CurveElementLocation from StepFEA);
	---Purpose: Writes CurveElementLocation

    Share (me; ent : CurveElementLocation from StepFEA;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWCurveElementLocation;
