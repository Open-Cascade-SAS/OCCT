-- Created on: 1999-04-14
-- Created by: Roman LYGIN
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SplitCurve2dContinuity from ShapeUpgrade inherits SplitCurve2d from ShapeUpgrade

    	---Purpose: Corrects/splits a 2d curve with a continuity criterion.
    	--  Tolerance is used to correct the curve at a knot that respects
    	--  geometrically the criterion, in order to reduce the
    	--  multiplicity of the knot.

uses

    Curve from Geom2d,
    Shape from GeomAbs

is

    Create returns SplitCurve2dContinuity from ShapeUpgrade;
        ---Purpose: Empty constructor.
	
    SetCriterion (me: mutable; Criterion: Shape from GeomAbs);
    	---Purpose: Sets criterion for splitting.
	
    SetTolerance (me: mutable; Tol: Real);
    	---Purpose: Sets tolerance.
	
    
    Compute(me: mutable) is redefined;
    	---Purpose: Calculates points for correction/splitting of the curve
    


fields

    myCriterion: Shape from GeomAbs;
    myCont     : Integer;
    myTolerance: Real;
    
end SplitCurve2dContinuity;
