-- Created on: 1997-04-24
-- Created by: Yves FRICAUD
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class SameShapeIterator from TNaming 

	---Purpose:  To iterate on   all  the label which contained  a
	--          given shape.

uses
    Shape       from TopoDS,
    UsedShapes  from TNaming,
    Iterator    from TNaming,
    Label       from TDF,
    PtrNode     from TNaming 	

raises
     NoMoreObject from Standard,
     NoSuchObject from Standard 

is

    Create(aShape      : Shape     from TopoDS; 
    	   Shapes      : UsedShapes from TNaming)
    returns SameShapeIterator from TNaming 
    is private;    

    Create(aShape      : Shape     from TopoDS; 
    	   access      : Label from TDF)
    returns SameShapeIterator from TNaming;
    
    More(me) returns Boolean;
    	---C++: inline
    
    Next(me : in out)
    raises
       NoMoreObject from Standard;
       
    Label(me) returns Label from TDF
    raises
	NoSuchObject from Standard;
	
fields
    myNode  : PtrNode from TNaming;	
    myIsNew   : Boolean from Standard;

friends

    class Tool from TNaming
    
end SameShapeIterator;
