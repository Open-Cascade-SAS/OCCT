-- Created on: 2003-09-29
-- Created by: Alexander SOLOVYOV and Sergey LITONIN
-- Copyright (c) 2003-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class SensitiveFace from MeshVS inherits SensitiveFace from Select3D

	---Purpose: This class provides custom sensitive face, which will be selected if it center is in rectangle.

uses
  EntityOwner from SelectBasics,

  Array1OfPnt from TColgp,

  TypeOfSensitivity from Select3D,
  Projector         from Select3D,

  Pnt   from gp,
  Pnt2d from gp,

  Array1OfPnt2d from TColgp,

  Box2d from Bnd

is

  Create ( theOwner    : EntityOwner from SelectBasics;
           thePoints   : Array1OfPnt from TColgp;
           theSensType : TypeOfSensitivity from Select3D = Select3D_TOS_INTERIOR )
    returns mutable SensitiveFace from MeshVS;

  Project( me: mutable; aProjector : Projector from Select3D ) is redefined;

  Matches  ( me: mutable; XMin, YMin, XMax, YMax: Real;
             aTol: Real ) returns Boolean is redefined;

  Matches  ( me: mutable; Polyline: Array1OfPnt2d from TColgp;
              aBox:Box2d; aTol: Real ) returns Boolean is redefined;

fields
  myCentre      : Pnt   from gp is protected;
  myProjCentre  : Pnt2d from gp is protected;

end SensitiveFace;
