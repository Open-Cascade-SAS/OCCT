-- File:	StepElement_CurveElementFreedom.cdl
-- Created:	Tue Dec 10 18:12:57 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V2.0
-- Copyright:	Open CASCADE 2002

class CurveElementFreedom from StepElement
inherits SelectType from StepData

    ---Purpose: Representation of STEP SELECT type CurveElementFreedom

uses
    SelectMember from StepData,
    EnumeratedCurveElementFreedom from StepElement,
    HAsciiString from TCollection

is
    Create returns CurveElementFreedom from StepElement;
	---Purpose: Empty constructor

    CaseNum (me; ent: Transient) returns Integer;
	---Purpose: Recognizes a kind of CurveElementFreedom select type
	--          return 0 

    CaseMem (me; ent: SelectMember from StepData) returns Integer is redefined;
	---Purpose: Recognizes a items of select member CurveElementFreedomMember
	--          1 -> EnumeratedCurveElementFreedom
	--          2 -> ApplicationDefinedDegreeOfFreedom
	--          0 else


     NewMember(me) returns SelectMember from StepData is redefined;
	---Purpose: Returns a new select member the type CurveElementFreedomMember

    SetEnumeratedCurveElementFreedom(me: in out; aVal :EnumeratedCurveElementFreedom from StepElement);
	---Purpose: Set Value for EnumeratedCurveElementFreedom

    EnumeratedCurveElementFreedom (me) returns EnumeratedCurveElementFreedom from StepElement;
	---Purpose: Returns Value as EnumeratedCurveElementFreedom (or Null if another type)

    SetApplicationDefinedDegreeOfFreedom(me: in out; aVal :HAsciiString from TCollection);
	---Purpose: Set Value for ApplicationDefinedDegreeOfFreedom

    ApplicationDefinedDegreeOfFreedom (me) returns HAsciiString from TCollection;
	---Purpose: Returns Value as ApplicationDefinedDegreeOfFreedom (or Null if another type)

end CurveElementFreedom;
