-- Created on: 1998-08-03
-- Created by: Christian CAILLET
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ToVRML  from XSDRAWSTLVRML

    ---Purpose : Writes a Shape to a File in VRML Format

uses CString, OStream, AsciiString from TCollection, Shape from TopoDS

is

    Create returns ToVRML;

    EmissiveColorRed   (me : in out) returns Real;
    ---C++ : return &
    EmissiveColorGreen (me : in out) returns Real;
    ---C++ : return &
    EmissiveColorBlue  (me : in out) returns Real;
    ---C++ : return &
    DiffuseColorRed    (me : in out) returns Real;
    ---C++ : return &
    DiffuseColorGreen  (me : in out) returns Real;
    ---C++ : return &
    DiffuseColorBlue   (me : in out) returns Real;
    ---C++ : return &
    Transparency       (me : in out) returns Real;
    ---C++ : return &
    AmbientIntensity   (me : in out) returns Real;
    ---C++ : return &
    SpecularColorRed   (me : in out) returns Real;
    ---C++ : return &
    SpecularColorGreen (me : in out) returns Real;
    ---C++ : return &
    SpecularColorBlue  (me : in out) returns Real;
    ---C++ : return &
    Shininess          (me : in out) returns Real;
    ---C++ : return &
    Texture            (me : in out) returns AsciiString;
    ---C++ : return &
    CreaseAngle        (me : in out) returns Real;
    ---C++ : return &
    Deflection         (me : in out) returns Real;
    ---C++ : return &


    Write (me; shape : Shape from TopoDS; filename : CString) returns Boolean;
    ---Purpose : conversion of a Shape into VRML format for 3d visualisation

fields

  myEmissiveColorRed   : Real;  -- def 0.3
  myEmissiveColorGreen : Real;  -- def 0.3
  myEmissiveColorBlue  : Real;  -- def 0.3
  myDiffuseColorRed    : Real;  -- def 0.3
  myDiffuseColorGreen  : Real;  -- def 0.3
  myDiffuseColorBlue   : Real;  -- def 0.5
  myTransparency       : Real;  -- def 0.0
  myAmbientIntensity   : Real;  -- def 0.3
  mySpecularColorRed   : Real;  -- def 0.7
  mySpecularColorGreen : Real;  -- def 0.7
  mySpecularColorBlue  : Real;  -- def 0.8
  myShininess          : Real;  -- def 0.1
  myTexture            : AsciiString;  -- def " [] "
  myCreaseAngle        : Real;  -- def 1.57
  myDeflection         : Real;  -- def 0.005

end ToVRML;
