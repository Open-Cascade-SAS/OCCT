-- Created on: 1998-03-04
-- Created by: Julia Gerasimova
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class BadEdgeFilter from AIS inherits Filter from SelectMgr

	---Purpose: A Class

uses

    EntityOwner                    from SelectMgr,
    Edge                           from TopoDS,
    DataMapOfIntegerListOfShape    from TopTools,    
    ShapeEnum                      from TopAbs
    
is
    Create
    returns mutable BadEdgeFilter from AIS;
    	--- Purpose: Constructs an empty filter object for bad edges.   
    ActsOn( me; aType : ShapeEnum from TopAbs )
    returns Boolean from Standard
    is redefined;
    
    IsOk( me; EO : EntityOwner from SelectMgr )
    returns Boolean from Standard is redefined virtual;

    SetContour( me : mutable ; Index : Integer from Standard );
    	---Purpose: sets  <myContour> with  current  contour. used  by
    	--          IsOk.

    AddEdge( me: mutable ; anEdge : Edge from TopoDS;
    	    	    	   Index : Integer from Standard );
    	---Purpose:  Adds an  edge  to the list  of non-selectionnable
    	--          edges.

    RemoveEdges( me: mutable ; Index : Integer from Standard );
    	---Purpose: removes from the  list of non-selectionnable edges
    	--          all edges in the contour <Index>.

fields

    myBadEdges : DataMapOfIntegerListOfShape from TopTools;
    myContour  : Integer                     from Standard;

end BadEdgeFilter;
