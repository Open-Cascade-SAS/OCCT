-- Created on: 1999-06-18
-- Created by: Sergei ZERTCHANINOV
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class FaceConnect  from ShapeFix

    ---Purpose : Rebuilds connectivity between faces in shell

uses 
    DataMapOfShapeListOfShape from TopTools,
    Face from TopoDS, Shell from TopoDS

is

    Create returns FaceConnect from ShapeFix;

    Add (me : in out; aFirst : Face from TopoDS; aSecond : Face from TopoDS)
    returns Boolean from Standard;
    ---Purpose : 

    Build (me : in out; shell : Shell from TopoDS;
    	   sewtoler : Real from Standard; fixtoler : Real from Standard)
    returns Shell from TopoDS;
    ---Purpose : 

    Clear (me : in out);
    ---Purpose : Clears internal data structure

fields

    myConnected    : DataMapOfShapeListOfShape from TopTools;
    	-- Map of pairs (face, list of connected faces) - to store connectivity info
    myOriFreeEdges : DataMapOfShapeListOfShape from TopTools;
    	-- Map of pairs (face, list of original free edges)
    myResFreeEdges : DataMapOfShapeListOfShape from TopTools;
    	-- Map of pairs (free edge, list of result free edges)
    myResSharEdges : DataMapOfShapeListOfShape from TopTools;
    	-- Map of pairs (free edge, list of result shared edges)

end FaceConnect;
