-- Created on: 1993-03-23
-- Created by: BBL,JLF
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Modified:    DCB (20-OCT-98)
--              Define Name()/SetName() as deferred.

deferred class AlienImageData from AlienImage inherits AlienImage

        ---Version: 0.0

        ---Purpose: This class defines an Alien image.
        -- Alien Image is X11 . xwd image or SGI .rgb image for examples

        ---Keywords:
        ---Warning:
        ---References:

uses
  AsciiString    from TCollection

is
        Initialize ;

        SetName( me : in out mutable;
                 aName : in AsciiString from TCollection)
        is virtual;
        ---Level: Public
        ---Purpose: Set Image name .

        Name( me : in immutable ) returns AsciiString from TCollection
        is virtual;
        ---C++: return const &
        ---Level: Public
        ---Purpose: get Image name .

fields
  myName:      AsciiString from TCollection is protected;

end AlienImageData;
 
