-- Created on: 2007-05-29
-- Created by: Vlad Romashko
-- Copyright (c) 2007-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Tick from TDataStd inherits Attribute from TDF

    ---Purpose: Defines a boolean attribute.
    --          If it exists at a label - true,
    --          Otherwise - false.

uses 

    Attribute         from TDF,
    Label             from TDF,
    GUID              from Standard,
    Integer           from Standard,
    DataSet           from TDF,
    RelocationTable   from TDF

is

    ---Purpose: Static methods
    --          ==============

    GetID (myclass)   
    ---C++: return const &  
    returns GUID from Standard;


    Set (myclass; label : Label from TDF)  
    ---Purpose: Find, or create, a Tick attribute.
    returns Tick from TDataStd;  


    ---Purpose: Tick methods
    --          ============

    Create
    returns mutable Tick from TDataStd;


    ---Category: Inherited methods
    --           =================

    ID (me)
    ---C++: return const & 
    returns GUID from Standard;

    Restore (me: mutable; With : Attribute from TDF);

    NewEmpty (me)
    returns mutable Attribute from TDF;

    Paste (me; Into : mutable Attribute from TDF;
	       RT   : mutable RelocationTable from TDF);    

    Dump (me; anOS : in out OStream from Standard)
    returns OStream from Standard
    is redefined;
    ---C++: return &


end Tick;
