-- File:        CameraModelD2.cdl
-- Created:     Mon Dec  4 12:02:24 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWCameraModelD2 from RWStepVisual

	---Purpose : Read & Write Module for CameraModelD2

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     CameraModelD2 from StepVisual,
     EntityIterator from Interface

is

	Create returns RWCameraModelD2;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable CameraModelD2 from StepVisual);

	WriteStep (me; SW : in out StepWriter; ent : CameraModelD2 from StepVisual);

	Share(me; ent : CameraModelD2 from StepVisual; iter : in out EntityIterator);

end RWCameraModelD2;
