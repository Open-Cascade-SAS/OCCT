-- Created on: 1999-11-26
-- Created by: Andrey BETENEV
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0

class RWCcDesignPersonAndOrganizationAssignment from RWStepAP203

    ---Purpose: Read & Write tool for CcDesignPersonAndOrganizationAssignment

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    CcDesignPersonAndOrganizationAssignment from StepAP203

is
    Create returns RWCcDesignPersonAndOrganizationAssignment from RWStepAP203;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : CcDesignPersonAndOrganizationAssignment from StepAP203);
	---Purpose: Reads CcDesignPersonAndOrganizationAssignment

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: CcDesignPersonAndOrganizationAssignment from StepAP203);
	---Purpose: Writes CcDesignPersonAndOrganizationAssignment

    Share (me; ent : CcDesignPersonAndOrganizationAssignment from StepAP203;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWCcDesignPersonAndOrganizationAssignment;
