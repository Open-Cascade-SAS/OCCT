-- Created on: 1992-12-15
-- Created by: Jean Louis FRENKEL
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



generic class WFShape from Prs3d 
     (FacePresentation   as any;        -- as WFRestrictedFace  from Prs3d
      CurvePresentation  as any;        -- as Curve             from Prs3d 
      PointPresentation  as any)        -- as Point             from Prs3d

inherits Root from Prs3d

uses
    Shape            from TopoDS,
    HSequenceOfShape from TopTools,
    Presentation     from Prs3d,
    Drawer           from Prs3d,
    Length           from Quantity
    
is
    Add(myclass; aPresentation: Presentation from Prs3d;
    	    	 aShape       : Shape        from TopoDS;
                 aDrawer      : Drawer       from Prs3d);
		 

    PickCurve(myclass; X,Y,Z     : Length from Quantity;
    	               aDistance : Length from Quantity;
                       aShape    : Shape  from TopoDS;
    	               aDrawer   : Drawer from Prs3d)
    returns HSequenceOfShape from TopTools;


    PickPatch(myclass; X,Y,Z     : Length from Quantity;
    	               aDistance : Length from Quantity;
                       aShape    : Shape  from TopoDS; 
    	               aDrawer   : Drawer from Prs3d)
    returns HSequenceOfShape from TopTools;
		   

end WFShape from Prs3d;
