-- Created on: 1992-07-28
-- Created by: Christian CAILLET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package Dico

    ---Purpose : Defines alphanumeric dictionaries and iterators on them
    --           Those are generic classes (Iterator is nested in Dictionary)
    --           Three default instantiations are offered :
    --           with Integer and Handle Objects (Persistent and Transient)

uses TCollection, MMgt, Standard

is

    generic class Dictionary,Iterator,StackItem;

    class DictionaryOfInteger    instantiates Dictionary (Integer);
    class DictionaryOfTransient  instantiates Dictionary (Transient);


end Dico;
