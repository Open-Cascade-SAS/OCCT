-- File:        FacetedBrepAndBrepWithVoids.cdl
-- Created:     Fri Jun 17 11:44:53 1994
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWFacetedBrepAndBrepWithVoids from RWStepShape

	---Purpose : Read & Write Module for FacetedBrepAndBrepWithVoids

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     FacetedBrepAndBrepWithVoids from StepShape,
     EntityIterator from Interface

is

	Create returns RWFacetedBrepAndBrepWithVoids;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable FacetedBrepAndBrepWithVoids from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : FacetedBrepAndBrepWithVoids from StepShape);

	Share(me; ent : FacetedBrepAndBrepWithVoids from StepShape; iter : in out EntityIterator);

end RWFacetedBrepAndBrepWithVoids;
