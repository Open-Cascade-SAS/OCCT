-- Created on: 1993-10-22
-- Created by: Gilles DEBARBOUILLE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class UnitsSystem from Units 
inherits

        TShared from MMgt  
	---Purpose: This class  allows  the  user  to  define his  own
	--          system of units.
  
uses

    AsciiString        from TCollection,
    HSequenceOfInteger from TColStd,
    QuantitiesSequence from Units
    


	
raises NoSuchUnit from Units,NoSuchType from Units

is

    Create returns mutable UnitsSystem from Units;
    
    ---Level: Public 
    
    ---Purpose: Returns an instance of UnitsSystem initialized to the 
    --          S.I. units system.

    Create(aName: CString from Standard;Verbose: Boolean from Standard = Standard_False)
    returns mutable UnitsSystem from Units;

    ---Level: Public 

    ---Purpose: Returns an instance of UnitsSystem initialized to the 
    --          S.I. units system upgraded by the base system units decription
    --	 	file.
    --          Attempts to find the four following files:
    --          $CSF_`aName`Defaults/.aName
    --          $CSF_`aName`SiteDefaults/.aName
    --          $CSF_`aName`GroupDefaults/.aName
    --          $CSF_`aName`UserDefaults/.aName
    --		See : Resource_Manager for the description of this file.
 
    QuantitiesSequence(me) returns QuantitiesSequence from Units;
    
    ---Level: Internal 
    
    ---Purpose: Returns the sequence of refined quantities.
    
    ActiveUnitsSequence(me) returns HSequenceOfInteger from TColStd;
    
    ---Level: Advanced 
    
    ---Purpose: Returns a sequence of integer in correspondance with 
    --          the sequence of quantities, which indicates, for each 
    --          redefined quantity, the index into the sequence of 
    --          units, of the active unit.
    
    Specify(me : mutable ; aquantity , aunit : CString)
    raises NoSuchType from Units
    ---Level: Public 
    
    ---Purpose: Specifies for <aquantity> the unit <aunit> used.

    is static;
    
    Remove(me : mutable ; aquantity , aunit : CString)
    
    ---Level: Public 
    
    ---Purpose: Removes for <aquantity> the unit <aunit> used.

    is static;
    
    Activate(me : mutable ; aquantity , aunit : CString)
    
    ---Level: Public 
    
    ---Purpose: Specifies for <aquantity> the unit <aunit> used.

    is static;

    Activates(me : mutable)
    
    ---Level: Public 
    
    ---Purpose: Activates the first unit of all defined system quantities

    is static;
    
    ActiveUnit(me ; aquantity : CString) returns AsciiString from TCollection
    
    ---Level: Public 
    
    ---Purpose: Returns for <aquantity> the active unit.

    is static;
    
    ConvertValueToUserSystem(me ; aquantity : CString ;
                                  avalue    : Real ;
                                  aunit     : CString) returns Real
    
    ---Level: Public 
    
    ---Purpose: Converts a real value <avalue> from the unit <aunit> 
    --          belonging to the physical dimensions <aquantity> to 
    --          the corresponding unit of the user system.

    is static;
    
    ConvertSIValueToUserSystem(me ; aquantity : CString ; avalue : Real) returns Real
    
    ---Level: Public 
    
    ---Purpose: Converts the real value <avalue> from the S.I. system 
    --          of units to the user system of units. <aquantity> is 
    --          the physical dimensions of the measurement.

    is static;
    
    ConvertUserSystemValueToSI(me ; aquantity : CString ; avalue : Real) returns Real

    ---Level: Public 
    
    ---Purpose: Converts the real value <avalue> from the user system 
    --          of units to the S.I. system of units. <aquantity> is 
    --          the physical dimensions of the measurement.

    is static;
    
    Dump(me)

    ---Level: Internal
    
    is static;

    IsEmpty(me) returns Boolean from Standard
    
    ---Level: Internal
    
    ---Purpose: Returns TRUE if no units has been defined in the system. 

    is static;

fields

    thequantitiessequence  : QuantitiesSequence from Units;
    theactiveunitssequence : HSequenceOfInteger from TColStd;

end UnitsSystem;
