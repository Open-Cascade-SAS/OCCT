-- Created on: 1994-11-14
-- Created by: Bruno DUMORTIER
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


private class MultiLineTool from BRepFill

    ---Purpose: private  class   used  to  instantiate the  continuous
    --          approximations routines.

uses
     Pnt           from gp,
     Pnt2d         from gp,
     Vec           from gp,
     Vec2d         from gp,
     Array1OfPnt   from TColgp,
     Array1OfPnt2d from TColgp,
     Array1OfVec   from TColgp,
     Array1OfVec2d from TColgp,
     MultiLine     from BRepFill

is
    
    FirstParameter(myclass; ML: MultiLine from BRepFill) 
    	---Purpose: returns the first parameter of the Line.
    returns Real from  Standard;


    LastParameter(myclass; ML: MultiLine from BRepFill) 
    	---Purpose: returns the last parameter of the Line.
    returns Real from Standard;


    NbP2d(myclass; ML: MultiLine from BRepFill) 
    	---Purpose: Returns the number of 2d points of a MLine
    returns Integer from Standard;


    NbP3d(myclass; ML: MultiLine from BRepFill) 
    	---Purpose: Returns the number of 3d points of a MLine.
    returns Integer from Standard;


    Value(myclass; ML   :     MultiLine   from BRepFill; 
    	    	   U    :     Real        from Standard; 
    	    	   tabPt: out Array1OfPnt from TColgp);
    	---Purpose: returns the 3d points of the multipoint <MPointIndex>
    	--          when only 3d points exist.


    Value(myclass; ML     :     MultiLine     from BRepFill; 
    	    	   U      :     Real          from Standard; 
                   tabPt2d: out Array1OfPnt2d from TColgp);
    	---Purpose: returns the 2d points of the multipoint <MPointIndex>
    	--          when only 2d points exist.


    Value(myclass; ML     :     MultiLine     from BRepFill;
    	    	   U      :     Real          from Standard; 
            	   tabPt  : out Array1OfPnt   from TColgp;
    	    	   tabPt2d: out Array1OfPnt2d from TColgp);
    	---Purpose: returns the 3d and 2d points of the multipoint 
    	--          <MPointIndex>.


    D1(myclass; ML  :     MultiLine   from BRepFill;
    	    	U   :     Real        from Standard; 
    	    	tabV: out Array1OfVec from TColgp)
    returns Boolean from Standard;
    	---Purpose: returns the 3d derivative values of the multipoint 
    	--          <MPointIndex> when only 3d points exist.
    	--          returns False if the derivative cannot be computed.


    D1(myclass; ML    :     MultiLine     from BRepFill; 
    	        U     :     Real          from Standard; 
    	        tabV2d: out Array1OfVec2d from TColgp)
    returns Boolean from Standard;
    	---Purpose: returns the 2d derivative values of the multipoint 
    	--          <MPointIndex> only when 2d points exist.
    	--          returns False if the derivative cannot be computed.


    D1(myclass; ML    :     MultiLine     from BRepFill; 
    	    	U     :     Real          from Standard; 
             	tabV  : out Array1OfVec   from TColgp; 
    	    	tabV2d: out Array1OfVec2d from TColgp)
    returns Boolean from Standard;
    	---Purpose: returns the 3d and 2d derivative values of the 
    	--          multipoint <MPointIndex>.
    	--          returns False if the derivative cannot be computed.

end MultiLineTool;    
    
