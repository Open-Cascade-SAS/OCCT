-- Created on: 2008-03-28
-- Created by: Sergey ZARITCHNY
-- Copyright (c) 2008-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class RealArrayRetrievalDriver_1 from MDataStd inherits ARDriver from MDF

	---Purpose: Retrieval  driver of RealArray attribute supporting 
	--          delta mechanism by default

uses
    RRelocationTable from MDF,
     Attribute        from TDF,
     Attribute        from PDF, 
     MessageDriver    from CDM
is

    Create(theMessageDriver : MessageDriver from CDM)  
    returns mutable RealArrayRetrievalDriver_1 from MDataStd;


    VersionNumber(me) returns Integer from Standard;
	---Purpose: Returns the version number from which the driver
	--          is available: 1.

    SourceType(me) returns Type from Standard;
	---Purpose: Returns the type: RealArray from PDataStd.

    NewEmpty (me) returns mutable Attribute from TDF;


    Paste(me;
    	  Source     :         Attribute from PDF;
    	  Target     : mutable Attribute from TDF;
    	  RelocTable : RRelocationTable from MDF);


end RealArrayRetrievalDriver_1;


