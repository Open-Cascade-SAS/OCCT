-- Created on: 1994-09-23
-- Created by: Yves FRICAUD
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class CutCurve from MAT2d 

	---Purpose: Cuts a curve at the extremas of curvature
	--          and at the inflections. Constructs a trimmed
	--          Curve for each interval.

uses
    Curve           from Geom2d,
    TrimmedCurve    from Geom2d,
    SequenceOfCurve from TColGeom2d,
    Side            from MAT
    
raises 
    OutOfRange from Standard
    
is
    Create;
    
    Create  (C : Curve from Geom2d) returns CutCurve from MAT2d;
    
    Perform (me : in out; C : Curve from Geom2d) 	    
	---Purpose: Cuts a curve at the extremas of curvature
	--          and at the inflections.
    is static;
    
    Perform (me : in out; C : Curve from Geom2d; aSide : Side from MAT)
    	---Purpose: Cuts a curve at the inflections, and at the extremas
    	--          of curvature where the concavity is on <aSide>. 
    is static;
    
    PerformInf (me : in out; C : Curve from Geom2d)    	
    	---Purpose: Cuts a curve at the inflections.
    is static;
    
    UnModified (me) returns Boolean from Standard
    	---Purpose: Returns True if the curve is not cut.
    is static;
    

    NbCurves (me) returns Integer from Standard
    	---Purpose: Returns the number of curves.
    	--          it's allways greatest than 2.    
    	--          
    	raises
    	    OutOfRange from Standard
	    ---Purpose: raises if the Curve is UnModified;        
    is static;
    

    Value (me ; Index : Integer from Standard) returns TrimmedCurve from Geom2d
	---Purpose: Returns the Indexth curve.    
        raises
    	    OutOfRange from Standard
	    ---Purpose: raises if Index not in the range [1,NbCurves()]
    is static;

    
fields
    theCurves : SequenceOfCurve from TColGeom2d;
    
end CutCurve;
