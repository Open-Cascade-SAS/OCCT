-- Created on: 1991-02-22
-- Created by: Jean Claude Vauthier
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package CPnts 

        --- Purpose :  
        --  This package  contains   the definition  of  the geometric
        --  algorithms   used to  compute  characteristic  points   on
        --  parametrized curves in 3d or 2d space. 
        --  This package defines the external geometric entities, with
        --  their requirements, used in the algorithms.

uses math, gp, StdFail, Adaptor3d  ,  Adaptor2d

is


   imported RealFunction;
    ---Purpose: typedef Standard_Real (*CPnts_RealFunction)
    --          (const Standard_Real, const Standard_Address)
    --          
    --          A pointer on a function for MyGaussFunction

   private class MyGaussFunction;
       ---Purpose: for implementation, compute values for Gauss

   private class MyRootFunction;
       ---Purpose: for implementation,  compute Length  and Derivative
       --          of the curve for Newton.

   class  AbscissaPoint;
       ---Purpose:  
       -- This algorithm computes a point and its parameter 
       -- as the distance between this and a given point is the abscissa

   class UniformDeflection;
        --- Purpose : This Algorithm computes a distribution of points 
        --  with a given chordal deviation on a parametrized curve.

end CPnts;








