-- Created on: 1993-06-14
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class BuilderON from TopOpeBRepBuild

uses

    PBuilder from TopOpeBRepBuild,
    PGTopo from TopOpeBRepBuild,
    PWireEdgeSet from TopOpeBRepBuild,
    ListOfShape from TopTools,
    Shape from TopoDS,
    Interference from TopOpeBRepDS,
    ListOfInterference from TopOpeBRepDS,
    Plos from TopOpeBRepTool

is
    -- BuilderON3d
    --------------
    Create returns BuilderON;
    Create(PB:PBuilder;F:Shape;PG:PGTopo;PLSclass:Plos;PWES:PWireEdgeSet) returns BuilderON;
    Perform(me:in out;PB:PBuilder;F:Shape;PG:PGTopo;PLSclass:Plos;PWES:PWireEdgeSet) is static;

    -- private
    GFillONCheckI(me;I:Interference) returns Boolean;
    GFillONPartsWES1(me:in out;I:Interference);
    GFillONPartsWES2(me:in out;I:Interference;EspON:Shape);


    -- BuilderON2d
    --------------
    Perform2d(me:in out;PB:PBuilder;F:Shape;PG:PGTopo;PLSclass:Plos;PWES:PWireEdgeSet) is static;
    
    -- private
    GFillONParts2dWES2(me:in out;I:Interference;EspON:Shape);
    
fields

    myPB : PBuilder from TopOpeBRepBuild;
    myPG : PGTopo from TopOpeBRepBuild;
    myPLSclass : Plos from TopOpeBRepTool;
    myPWES : PWireEdgeSet from TopOpeBRepBuild;
    myFace : Shape from TopoDS;
    
    myFEI : ListOfInterference from TopOpeBRepDS; --BuilderON2d 
    
end BuilderON from TopOpeBRepBuild;
