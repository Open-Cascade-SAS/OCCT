-- Created on: 1993-03-24
-- Created by: JCV
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Direction  from Geom2d inherits Vector from Geom2d 

        --- Purpose :
        --  The class Direction specifies a vector that is never null.
        --  It is a unit vector.


uses  Dir2d    from gp,
      Pnt2d    from gp, 
      Trsf2d   from gp,
      Vec2d    from gp,
      Geometry from Geom2d

raises ConstructionError from Standard

is


  Create (X, Y :Real)  returns Direction
        --- Purpose : Creates a unit vector with it 2 cartesian coordinates.
     raises ConstructionError;
        --- Purpose : 
        --  Raised if Sqrt( X*X + Y*Y) <= Resolution from gp.

  Create (V : Dir2d) returns Direction;
        --- Purpose : Creates a persistent copy of <me>.


  
  SetCoord (me : mutable; X, Y : Real)
        --- Purpose : Assigns the coordinates X and Y to this unit vector,
    	-- then normalizes it.
    	-- Exceptions
    	-- Standard_ConstructionError if Sqrt(X*X +
    	-- Y*Y) is less than or equal to gp::Resolution().
     raises ConstructionError;
     

  SetDir2d (me : mutable; V : Dir2d);
        --- Purpose : Converts the gp_Dir2d unit vector V into this unit vector.


  SetX (me : mutable; X : Real)
        --- Purpose : 
    	-- Assigns a value to the X coordinate of this unit vector, then normalizes it.
    	-- Exceptions
    	-- Standard_ConstructionError if the value assigned
    	-- causes the magnitude of the vector to become less
    	-- than or equal to gp::Resolution().
     raises ConstructionError;
    

  SetY (me : mutable; Y : Real)
        --- Purpose : Assigns a value to the Y coordinate of this unit vector, then normalizes it.
    	-- Exceptions
    	-- Standard_ConstructionError if the value assigned
    	-- causes the magnitude of the vector to become less
    	-- than or equal to gp::Resolution().
     raises ConstructionError;
       

  Dir2d (me) returns Dir2d;
        --- Purpose : Converts this unit vector into a gp_Dir2d unit vector.
      

  Magnitude (me)   returns Real;
        --- Purpose : returns 1.0


  SquareMagnitude (me)   returns Real;
        --- Purpose : returns 1.0


  Crossed (me; Other : Vector)  returns Real;
        --- Purpose : Computes the cross product between <me> and <Other>.
        ---C++: alias operator ^
     

  Transform (me : mutable; T : Trsf2d);

    	---Purpose: Applies the transformation T to this unit vector, then normalizes it.


  Copy (me)  returns like me;
    	---Purpose: Creates a new object which is a copy of this unit vector.     
end;

