-- Created on: 1995-08-09
-- Created by: Arnaud BOUZY
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Point from AIS inherits InteractiveObject from AIS

	---Purpose: Constructs point datums to be used in construction of
    	-- composite shapes. The datum is displayed as the plus marker +.

uses 
    Point                 from Geom,
    TypeOfMarker          from Aspect,
    Presentation          from Prs3d,
    PresentationManager3d from PrsMgr,
    NameOfColor           from Quantity,
    Color			  from Quantity,
    Selection             from SelectMgr,
    Projector             from Prs3d,
    Transformation        from Geom,
    Vertex                from TopoDS,
    KindOfInteractive     from AIS   


is
    Create(aComponent : Point from Geom) 
    returns Point from AIS;
    	---Purpose:
    	-- Initializes the point aComponent from which the point
    	-- datum will be built.

    Signature(me) returns Integer from Standard is redefined;
   	 ---Purpose: Returns index 1, the default index for a point.
   	 ---C++: inline

    Type(me) returns KindOfInteractive from AIS is redefined;
    	---Purpose: Indicates that a point is a datum.
        ---C++: inline

    Component(me: mutable) returns Point from Geom 
    is static;
    	---Purpose: Returns the component specified in SetComponent.
    SetComponent(me: mutable;aComponent:Point from Geom )
    is static;
    	---Purpose: Constructs an instance of the point aComponent.
    AcceptDisplayMode(me;aMode:Integer from Standard) returns Boolean from  Standard is redefined static;
    	---Purpose: Returns true if the display mode selected is valid for point datums.

    Compute(me            : mutable;
    	    aPresentationManager: PresentationManager3d from PrsMgr;
    	    aPresentation : Presentation from Prs3d;
    	    aMode         : Integer from Standard = 0) 
    is redefined virtual protected;
    
    Compute(me:mutable;
    	        aProjector: Projector from Prs3d;
                aPresentation: Presentation from Prs3d)
    is redefined static private;

    Compute(me            : mutable;
            aProjector    : Projector from Prs3d;
            aTrsf         : Transformation from Geom;
            aPresentation : Presentation from Prs3d)
    is redefined;
    	---Purpose: computes the presentation according to a point of view
    	--          given by <aProjector>.
    	--          To be Used when the associated degenerated Presentations
    	--          have been transformed by <aTrsf> which is not a Pure
   	--          Translation. The HLR Prs can't be deducted automatically
    	--          WARNING :<aTrsf> must be applied
    	--           to the object to display before computation  !!!

-- Methods from SelectableObject

    ComputeSelection(me         : mutable;
    	    	     aSelection : Selection from SelectMgr;
    	    	     aMode      : Integer from Standard )is private;

-- Methods from InteractiveObject

    SetColor(me :mutable; aColor : NameOfColor from Quantity) 
    is redefined static;
    	---Purpose: Allows you to provide settings for the cp;pr aColor.
    SetColor(me :mutable; aColor : Color from Quantity) 
    is redefined static;

    UnsetColor(me:mutable) is redefined static;
    	---Purpose: Allows you to remove color settings.
    SetMarker(me:mutable; aType : TypeOfMarker from Aspect);
    	---Purpose: Allows you to provide settings for a marker. These include
    	-- -   type of marker,
    	-- -   marker color,
    	-- -   scale factor.    
    
    UnsetMarker(me:mutable);
    	---Purpose: Removes the marker settings.    
    HasMarker(me) returns Boolean from Standard;
    	---Purpose: Returns true if the point datum has a marker.
    	---C++: inline

    Vertex(me) returns Vertex from TopoDS;
    	---Purpose: Converts a point into a vertex.
    UpdatePointValues(me:mutable) is private;
    	---Level: Internal 
		   


fields

    myComponent   : Point from Geom;
    myHasTOM      : Boolean from Standard; 
    myTOM         : TypeOfMarker from Aspect;    
end Point;
