-- Created on: 1993-07-06
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.





class MakeVertex from BRepBuilderAPI inherits MakeShape from BRepBuilderAPI

	---Purpose: Describes functions to build BRepBuilder vertices directly
    	-- from 3D geometric points. A vertex built using a
    	-- MakeVertex object is only composed of a 3D point and
    	-- a default precision value (Precision::Confusion()).
    	-- Later on, 2D representations can be added, for example,
    	-- when inserting a vertex in an edge.
    	-- A MakeVertex object provides a framework for:
    	-- -   defining and implementing the construction of a vertex, and
    	-- -   consulting the result.

uses
    Pnt        from gp,
    Vertex     from TopoDS,
    MakeVertex from BRepLib

is
    Create (P : Pnt from gp) 
	---Purpose: Constructs a vertex from point P.
    	-- Example create a vertex from a 3D point.
    	-- gp_Pnt P(0,0,10);
    	-- TopoDS_Vertex V = BRepBuilderAPI_MakeVertex(P);
    returns MakeVertex from BRepBuilderAPI;
    
    Vertex(me) returns Vertex from TopoDS
	---C++: return const &
	---C++: alias "Standard_EXPORT operator TopoDS_Vertex() const;"
    	---Purpose: Returns the constructed vertex.
    is static;
    
fields

    myMakeVertex : MakeVertex from BRepLib;	   
	       

end MakeVertex;
