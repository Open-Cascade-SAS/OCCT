-- Created on: 1993-07-06
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class Curve3D from PBRep inherits GCurve from PBRep

	---Purpose: Representation of a curve by a 3D curve.

uses

    Location from PTopLoc,
    Curve    from PGeom

is

    Create(C  : Curve    from PGeom;
    	   CF : Real     from Standard;
	   CL : Real     from Standard;
    	   L  : Location from PTopLoc) 
    returns mutable Curve3D from PBRep;
    	---Purpose : CF is curve first param
    	--           CL is curve last param
    	--           As far as they can't be computed from a Persistent Curve
    	--          they are given in the Curve3D constructor

    Curve3D(me) returns Curve from PGeom
    is static;

    IsCurve3D(me) returns Boolean
	 ---Purpose: Returns True.
    is redefined;
	
fields
    
    myCurve3D : Curve from PGeom;

end Curve3D;
