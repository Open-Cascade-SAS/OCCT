-- Created on: 1999-09-16
-- Created by: Edward AGAPOV
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class ExtPExtS from Extrema 
		    
	---Purpose: It calculates all the extremum (minimum and
	--          maximum) distances between a point and a linear
	--          extrusion surface.
		    
uses
    POnSurf from Extrema,
    GenExtPS from Extrema,
    FuncExtPS from Extrema,
    
    HCurve from Adaptor3d,
    SurfacePtr from Adaptor3d, 
    SurfaceOfLinearExtrusion from Adaptor3d,
    
    Ax2 from gp,
    Vec from gp,
    Pnt from gp

raises 
    NotDone from StdFail,
    OutOfRange


is
    Create returns ExtPExtS;

    Create (P: Pnt; S: SurfaceOfLinearExtrusion from Adaptor3d; 
		    Umin, Usup, Vmin, Vsup: Real; 
		    TolU,TolV: Real) 
		    returns ExtPExtS;
    ---Purpose: It calculates all the distances between a point 
    --          from gp and a Surface.
    
    Create (P: Pnt; S: SurfaceOfLinearExtrusion from Adaptor3d; 
		    TolU,TolV: Real) 
		    returns ExtPExtS;
    ---Purpose: It calculates all the distances between a point 
    --          from gp and a Surface.

    Initialize(me: in out; S: SurfaceOfLinearExtrusion from Adaptor3d;
    			   Uinf, Usup, Vinf, Vsup: Real;
			   TolU, TolV: Real)
    ---Purpose: Initializes the fields of the algorithm.
		    is static;

    Perform(me: in out; P: Pnt)
		    is static;
    
    IsDone (me) returns Boolean
    ---Purpose: Returns True if the distances are found.
    		    is static;
    
    NbExt (me) returns Integer
    ---Purpose: Returns the number of extremum distances.
    		    raises  NotDone from StdFail
	    	-- if IsDone(me)=False.
    		    is static;

    SquareDistance (me; N: Integer) returns Real
    ---Purpose: Returns the value of the Nth resulting square distance.
    		    raises  NotDone from StdFail,
    	    	-- if IsDone(me)=False.
    	        OutOfRange
		-- if N < 1 or N > NbPoints(me).
    		    is static;

    Point (me; N: Integer) returns POnSurf
    ---C++: return const &
    ---Purpose: Returns the point of the Nth resulting distance.
    		    raises  NotDone from StdFail,
    	    	-- if IsDone(me)=False.
    	        OutOfRange
		-- if N < 1 or N > NbPoints(me).
    		    is static;

    --- Private methods
    
    MakePreciser (me; U : in out Real from Standard;
		      P : Pnt from gp;
		      isMin : Boolean from Standard;
		      OrtogSection: Ax2 from gp) is static private;

fields
    myuinf   : Real from Standard;
    myusup   : Real from Standard;
    mytolu   : Real from Standard;
    myvinf   : Real from Standard;
    myvsup   : Real from Standard;
    mytolv   : Real from Standard;
    
    myF	        : FuncExtPS  from Extrema;
    myC         : HCurve     from Adaptor3d; 
    myS	        : SurfacePtr from Adaptor3d;
    myDirection : Vec        from gp;
    myPosition  : Ax2        from gp;
    myExtPS     : GenExtPS   from Extrema;
    
    myIsAnalyticallyComputable : Boolean  from Standard;

    myDone : Boolean from Standard;
    myNbExt: Integer from Standard;
    mySqDist: Real    from Standard [4];
    myPoint: POnSurf from Extrema  [4];
    
end ExtPExtS;
