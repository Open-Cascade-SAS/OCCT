-- Created on: 1993-06-07
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ArcFunction from IntPatch

inherits FunctionWithDerivative from math

uses
     HCurve2d      from Adaptor2d,
     HSurface      from Adaptor3d,
     Pnt           from gp,
     SequenceOfPnt from TColgp,
     Quadric       from IntSurf

is

    Create
    
    	returns ArcFunction from IntPatch;


    SetQuadric(me: in out; Q: Quadric from IntSurf)
    
	---C++: inline
    	is static;


    Set(me: in out; A: HCurve2d from Adaptor2d)
    
	---C++: inline
    	is static;


    Set(me: in out; S: HSurface from Adaptor3d)
    
	---C++: inline
    	is static;


    Value(me: in out; X: Real from Standard; F: out Real from Standard)
    
    	returns Boolean from Standard;
    

    Derivative(me: in out; X: Real from Standard; D: out Real from Standard)
    
    	returns Boolean from Standard;
    

    Values(me: in out; X: Real from Standard; F,D: out Real from Standard)
    
    	returns Boolean from Standard;
    

    NbSamples(me)
    
    	returns Integer from Standard
	is static;


    GetStateNumber(me: in out)

    	returns Integer from Standard
    	is redefined;
	
	
    Valpoint(me; Index: Integer from Standard)
    
    	returns Pnt from gp
	---C++: return const&
	---C++: inline
	is static;
    
    Quadric(me) 
    	returns Quadric from IntSurf
	---C++: return const&
	---C++: inline
	is static;
       
    Arc(me)
   	returns HCurve2d from Adaptor2d
	---C++: return const&
	---C++: inline
	is static;
       
    Surface(me)
   	returns HSurface from Adaptor3d
	---C++: return const&
	---C++: inline
	is static;
	    
fields

    myArc  : HCurve2d      from Adaptor2d;
    mySurf : HSurface      from Adaptor3d;
    myQuad : Quadric       from IntSurf;
    ptsol  : Pnt           from gp;
    seqpt  : SequenceOfPnt from TColgp;

end ArcFunction;
