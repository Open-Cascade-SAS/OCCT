-- File:        SurfaceStyleSilhouette.cdl
-- Created:     Fri Dec  1 11:11:28 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class SurfaceStyleSilhouette from StepVisual 

inherits TShared from MMgt

uses

	CurveStyle from StepVisual
is

	Create returns mutable SurfaceStyleSilhouette;
	---Purpose: Returns a SurfaceStyleSilhouette

	Init (me : mutable;
	      aStyleOfSilhouette : mutable CurveStyle from StepVisual) is virtual;

	-- Specific Methods for Field Data Access --

	SetStyleOfSilhouette(me : mutable; aStyleOfSilhouette : mutable CurveStyle);
	StyleOfSilhouette (me) returns mutable CurveStyle;

fields

	styleOfSilhouette : CurveStyle from StepVisual;

end SurfaceStyleSilhouette;
