-- Created on: 1997-10-29
-- Created by: Roman BORISOV
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Assembly from FEmTool

	---Purpose: Assemble and solve system from (one dimensional) Finite Elements  

uses 
    Array2OfInteger  from  TColStd, 
    HAssemblyTable  from  FEmTool, 
    Matrix  from  math, 
    Vector  from  math,	     
    ProfileMatrix  from  FEmTool, 
    SeqOfLinConstr  from  FEmTool, 
    SequenceOfReal  from  TColStd 
    
raises   
        NotDone  from  StdFail, 
        DimensionError, 
	DomainError
is 
    Create(Dependence :  Array2OfInteger  from  TColStd; 
           Table      :  HAssemblyTable  from  FEmTool)   
    returns  Assembly from FEmTool; 
     
    NullifyMatrix(me : in  out); 
    ---Purpose: Nullify all Matrix 's Coefficient
           
    AddMatrix(me  : in  out;   
              Element    :  Integer; 
	      Dimension1 :  Integer; 
	      Dimension2 :  Integer; 
              Mat  :  Matrix  from  math)
    ---Purpose: Add an elementary Matrix in the assembly Matrix 
    	raises  DomainError; --  if  Dependence(Dimension1,Dimension2)  is  False
              
    NullifyVector(me : in  out);                
    ---Purpose:  Nullify  all  Coordinate of  assembly  Vector (second member)
     
    AddVector(me  :  in  out; 
              Element    :  Integer; 
	      Dimension  :  Integer; 
              Vec  :  Vector  from  math);  
    ---Purpose: Add an elementary Vector in the assembly Vector (second member)     

    ResetConstraint(me : in  out);                
    ---Purpose: Delete all Constraints.
    
    NullifyConstraint(me : in  out);                
    ---Purpose: Nullify all Constraints.   
     
    AddConstraint(me : in  out; 
            IndexofConstraint :  Integer;
            Element           :  Integer; 
            Dimension         :  Integer;	     
            LinearForm        :  Vector  from  math;
            Value             :  Real); 
	         
     
    Solve(me  :  in  out)  returns  Boolean; 
    ---Purpose: Solve the assembly system         
    --          Returns Standard_False if the computation failed.
     
    Solution(me;  Solution : out  Vector  from  math) 
    raises  NotDone  from  StdFail;  -- if the system is not solved.  
     
    NbGlobVar(me) 
    returns  Integer; 
     
    GetAssemblyTable(me;  AssTable  :  out  HAssemblyTable  from  FEmTool);
	      
fields  
    myDepTable  :  Array2OfInteger;
    myRefTable  :  HAssemblyTable; 
    IsSolved    :  Boolean;
    H           :  ProfileMatrix  from  FEmTool;  
    B	        :  Vector  from  math;
    GHGt        :  ProfileMatrix  from  FEmTool; 
    G	        :  SeqOfLinConstr  from  FEmTool; 
    C           :  SequenceOfReal  from  TColStd;     
end Assembly;

