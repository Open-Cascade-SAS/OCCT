-- Created on: 1995-03-10
-- Created by: Remi LEQUETTE
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Box from Draw inherits Drawable3D from Draw

	---Purpose: 

uses Pnt from gp,
    Color from Draw,
    Display from Draw

is

    Create(p1,p2 : Pnt; col : Color)
    returns mutable Box;
    
    DrawOn(me; dis : in out Display);
    
    First(me) returns Pnt from gp
	---C++: return const&
    is static;

    First(me : mutable; P : Pnt from gp)
    is static;

    Last(me) returns Pnt from gp
	---C++: return const&
    is static;

    Last(me : mutable; P : Pnt from gp)
    is static;

fields

    myFirst : Pnt;
    myLast  : Pnt;
    myColor : Color;
    
end Box;
