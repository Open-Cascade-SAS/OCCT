-- Created on: 2008-09-01
-- Created by: Vladislav ROMASHKO
-- Copyright (c) 2008-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

private class SplitData from Voxel

    ---Purpose: A container of split information.
    --          An instance of this class is used as a slice 
    --          in inner representation of recursive octtree voxels.

is

    Create
    ---Purpose: An empty constructor.
    returns SplitData from Voxel;

    GetValues(me : in out)
    ---Purpose: Gives access to the values.
    ---C++: return &
    returns Address from Standard;

    GetSplitData(me : in out)
    ---Purpose: Gives access to the next split data.
    ---C++: return &
    returns Address from Standard;

fields

    myValues    : Address from Standard;
    mySplitData : Address from Standard;
    
end SplitData;

