-- File:	DrawDim_Radius.cdl
-- Created:	Mon Apr 21 13:36:26 1997
-- Author:	Denis PASCAL
--		<dp@dingox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1997



class Radius from DrawDim inherits Dimension from DrawDim

	---Purpose: 

uses Face    from TopoDS,
     Display from Draw

is

    Create (cylinder : Face from TopoDS)
    returns mutable Radius from DrawDim;
    
    Cylinder (me) returns Face from TopoDS;
    ---C++: return const&

    Cylinder (me : mutable; face : Face from TopoDS);    

    DrawOn (me; dis : in out Display);
    
fields

    myCylinder : Face from TopoDS;
    
end Radius;

