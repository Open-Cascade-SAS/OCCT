-- Created by: Peter KURNEV
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement. 

 
class BOP from BOPAlgo  
    inherits Builder from BOPAlgo
 
---Purpose: 

uses 
    ShapeEnum from TopAbs,
    Shape from TopoDS,   
    ListOfShape from TopTools, 
    --
    BaseAllocator from BOPCol,  
    ListOfShape from BOPCol, 
    MapOfShape  from BOPCol, 
    IndexedDataMapOfShapeListOfShape from BOPCol, 
    --
    Operation  from BOPAlgo, 
    PaveFiller from BOPAlgo 

--raises

is
    Create 
    ---Purpose:  Empty constructor     
        returns BOP from BOPAlgo;  
    ---C++: alias "Standard_EXPORT virtual ~BOPAlgo_BOP();"  
      
    Create (theAllocator: BaseAllocator from BOPCol)
        returns BOP from BOPAlgo; 
	 
    Clear(me:out) 
    is redefined; 
    ---Purpose:  Clears internal fields and arguments   
     
    AddTool (me:out;  
            theShape: Shape from TopoDS) 
    ---Purpose:  Adds Tool argument of the operation    	     
        is virtual;  
        
    SetTools (me:out;
            theShapes: ListOfShape from TopTools)
        is virtual;  
         
    SetTools (me:out;
            theShapes: ListOfShape from BOPCol)
        is virtual; 
 
    SetOperation(me:out;  
            theOperation: Operation from BOPAlgo); 
	 
    Operation(me) 
        returns Operation from BOPAlgo; 
    -- 
    Perform(me:out) 
        is redefined;  
    --
    --  protected methods 
    -- 
    CheckData(me:out) 
        is redefined protected; 

    Prepare(me:out)  
        is redefined protected; 
    ---Purpose:  Provides preparing actions 

    PerformInternal1(me:out; 
            thePF:PaveFiller from BOPAlgo) 
        is redefined protected;   
    ---Purpose:  Performs calculations using prepared Filler 
    --           object <thePF>          	 
     
    BuildResult(me:out; 
            theType: ShapeEnum from TopAbs) 
        is redefined protected;     
     
    BuildShape(me:out) 
        is protected; 
 
    BuildRC(me:out) 
        is protected; 
 
    BuildSolid(me:out) 
        is protected; 
 
    IsBoundSplits(me:out; 
            theS:Shape from TopoDS; 
            theMEF:out IndexedDataMapOfShapeListOfShape from BOPCol)  
        returns Boolean from Standard
        is protected;
 
fields 
    myOperation : Operation from BOPAlgo   is protected; 
    myDims      : Integer from Standard[2] is protected;  
    -- 
    myRC        : Shape from TopoDS        is protected; 
    myTools     : ListOfShape from BOPCol  is protected; 
    myMapTools  : MapOfShape  from BOPCol  is protected;  
    
end BOP;
