-- Created on: 2008-08-28
-- Created by: Vladislav ROMASHKO
-- Copyright (c) 2008-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Reader from Voxel

    ---Purpose: Reads a cube of voxels from disk.
    --          Beware, a caller of the reader is responsible for deletion of the read voxels.

uses

    BoolDS          from Voxel,
    ColorDS         from Voxel,
    FloatDS         from Voxel,
    ExtendedString  from TCollection

is

    Create
    ---Purpose: An empty constructor.
    returns Reader from Voxel;

    Read(me : in out;
    	 file : ExtendedString from TCollection)
    ---Purpose: Reads the voxels from disk
    returns Boolean from Standard;

    IsBoolVoxels(me)
    ---Purpose: Informs the user about the type of voxels he has read.
    returns Boolean from Standard;

    IsColorVoxels(me)
    ---Purpose: Informs the user about the type of voxels he has read.
    returns Boolean from Standard;

    IsFloatVoxels(me)
    ---Purpose: Informs the user about the type of voxels he has read.
    returns Boolean from Standard;

    GetBoolVoxels(me)
    ---Purpose: Returns a pointer to the read 1bit voxels.
    returns Address from Standard;

    GetColorVoxels(me)
    ---Purpose: Returns a pointer to the read 4bit voxels.
    returns Address from Standard;

    GetFloatVoxels(me)
    ---Purpose: Returns a pointer to the read 4bytes voxels.
    returns Address from Standard;


    ---Private area
    -- ============

    ReadBoolAsciiVoxels(me : in out;
    	    	    	file : ExtendedString from TCollection)
    ---Purpose: Reads 1bit voxels from disk in ASCII format.
    returns Boolean from Standard
    is private;

    ReadColorAsciiVoxels(me : in out;
    	    	     	 file : ExtendedString from TCollection)
    ---Purpose: Reads 4bit voxels from disk in ASCII format.
    returns Boolean from Standard
    is private;

    ReadFloatAsciiVoxels(me : in out;
    	    	    	 file : ExtendedString from TCollection)
    ---Purpose: Reads 4bytes voxels from disk in ASCII format.
    returns Boolean from Standard
    is private;

    ReadBoolBinaryVoxels(me : in out;
    	    	    	 file : ExtendedString from TCollection)
    ---Purpose: Reads 1bit voxels from disk in BINARY format.
    returns Boolean from Standard
    is private;

    ReadColorBinaryVoxels(me : in out;
    	    	     	  file : ExtendedString from TCollection)
    ---Purpose: Reads 4bit voxels from disk in BINARY format.
    returns Boolean from Standard
    is private;

    ReadFloatBinaryVoxels(me : in out;
    	    	    	  file : ExtendedString from TCollection)
    ---Purpose: Reads 4bytes voxels from disk in BINARY format.
    returns Boolean from Standard
    is private;


fields

    myBoolVoxels  : Address from Standard;
    myColorVoxels : Address from Standard;
    myFloatVoxels : Address from Standard;

end Reader;
