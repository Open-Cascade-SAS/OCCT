-- Created on: 1998-01-08
-- Created by: Isabelle GRIGNON
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Document from PCDMShape inherits Document from PCDM


    ---Purpose: This document is used to store a Shape1 from PTopoDS.
    
uses

    Orientation   from TopAbs,
    Shape1        from PTopoDS,
    Location      from PTopLoc
    
is
    Create returns mutable Document from PCDMShape;
    ---Level: Internal 

    Create(T : Shape1 from PTopoDS) returns mutable Document from PCDMShape;
    ---Level: Internal 

    Shape(me) returns Shape1 from PTopoDS
    ---Level: Internal 
    ---C++: return const
    is static;

    Shape(me : mutable; T : Shape1 from PTopoDS)
    ---Level: Internal 
    is static;

fields

    myShape : Shape1 from PTopoDS;

end Document from PCDMShape;
