-- Created on: 1999-03-03
-- Created by: Fabrice SERVANT
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Modified by skv - Thu Sep 25 18:04:05 2003 OCC567 
-- Definition of new pointer to MaillageAffinage 
-- which is used in Intersection class.

package IntPolyh 

	---Purpose:  This   package  provides algorithms    to compute
	--           starting   points for   the     surface  surface
	--           intersection  packages. Those  starting points are
	--           used if   the  two   surfaces are  bi-parametric
	--           surfaces (bezier, nurbs, algorithm surfaces ...)
	--          
    	--  This package provides methods 
    	--     
    	--      to compute meshes on the  two surfaces. The meshes can
    	--      be refined if  necessary.  It is the major improvement
    	--      to  the Intf  package which   gives  the same  kind of
    	--      ressources.
        --
        --      to intersect the two meshes
        --
        --      to give approximated starting-points. Those points are
        --      organised in lines, when  the points belong to a  same
        --      section line, or returned as isolated points when they
        --      can neither  define a  new  line nor  be  linked to an
        --      existant line.
        --      
        --  A  starting-point   contains 3d   information,  parametric
        --  ionformation and  quality criterion. (i.e.   X,Y,Z, U1,V1,
        --  U2,V2,  Incidence).  Incidence  is  a real wich   gives an
        --  estimated   angle    between the two   surfaces  near  the
        --  intersection point.
        --  
        --  

uses
    TCollection,
    TColStd,
    gp, 	      
    Bnd,
    Adaptor3d
 
is 
    imported ArrayOfSectionLines from IntPolyh; 
    imported ArrayOfCouples from IntPolyh; 
    imported ArrayOfEdges from IntPolyh; 
    imported ArrayOfPoints from IntPolyh; 
    imported ArrayOfStartPoints from IntPolyh; 
    imported ArrayOfTangentZones from IntPolyh; 
    imported ArrayOfTriangles from IntPolyh; 
    
    class Intersection;
	---Purpose:  the main   algorithm.  Algorythm   outputs are --
	--            lines  and  points like   discribe   in the last
	--          paragraph.  The Algorythm provides direct acces to
	--            the elements of those   lines  and points. Other
	--          classes  of this package  are for internal use and
	--          only concern the algorithmic part.

    ------------------------------------------------------------
    ----   Internal classes and algorithms 
    ------------------------------------------------------------
    class Couple;
	---Purpose: couple of triangles


    class Point;
    class StartPoint;
    class SeqOfStartPoints instantiates Sequence from TCollection
        (StartPoint from IntPolyh);

    class Edge;
     

    class Triangle;
    
   
    class MaillageAffinage;
    	---Purpose: Provide the algorythms used in the package

    class SectionLine;
    
    
--    class TangentZone; For the moment we use the StartPoint Class
    
    pointer PMaillageAffinage to MaillageAffinage from IntPolyh;
    
end;









