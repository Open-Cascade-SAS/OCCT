-- Created on: 1993-04-06
-- Created by: Philippe DAUTRY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Transformation from PGeom2d inherits Persistent from Standard

        ---Purpose :  The    class Transformation  allows   to  create
        --         Translation, Rotation,   Symmetry,     Scaling  and
        --         complex transformations obtained by  combination of
        --         the  previous elementary   transformations.     The
        --         restriction to  these basic  transformations allows
        --         us to be sure that   an object  will never   change
        --         nature.
        --         
	---See Also : Transformation from Geom2d.


uses Trsf2d from gp

is


  Create returns mutable Transformation from PGeom2d;
        ---Purpose : Creates a transformation with default values.
	---Level: Internal 


  Create (aTrsf : Trsf2d from gp) returns mutable Transformation from PGeom2d;
        ---Purpose :  Creates a transformation with <aTrsf>.
	---Level: Internal 


  Trsf (me : mutable; aTrsf : Trsf2d from gp);
        ---Purpose : Creates a Transformation with <aTrsf>.
	---Level: Internal 


  Trsf (me)  returns Trsf2d from gp;
        ---Purpose : Returns the value of the field trsf.
	---Level: Internal 


fields

  trsf : Trsf2d from gp;

end;
