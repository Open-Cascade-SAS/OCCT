-- Created on: 1999-10-21
-- Created by: Denis PASCAL
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Naming from PNaming inherits Attribute from PDF

	---Purpose: 

uses 
    Name from PNaming
			    
is
    Create
    returns Naming from PNaming;
    
    SetName(me : mutable ; aName : Name from PNaming);

    GetName(me) returns Name from PNaming;

fields

    myName :  Name from PNaming;

end Naming;
