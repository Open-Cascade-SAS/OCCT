-- Created on: 1993-09-01
-- Created by: Laurent PAINNOT
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



deferred class Function from AppCont

    ---Purpose: deferred class describing a continous 3d function f(u)


uses Pnt from gp,
     Vec from gp

is

    Delete(me:out) is virtual;
    ---C++: alias "Standard_EXPORT virtual ~AppCont_Function(){Delete() ; }"
    

    FirstParameter(me) returns Real
    	---Purpose: returns the first parameter of the function.
    is deferred;

    LastParameter(me) returns Real
    	---Purpose: returns the last parameter of the function.
    is deferred;

    Value(me; U: Real) returns Pnt
    	---Purpose: returns the point at parameter <U>.
    is deferred;

    D1(me; U: Real; P: in out Pnt; V: in out Vec) returns Boolean
    	---Purpose: returns the point and the derivative values at
    	--          the parameter <U>.
    is deferred;
    
    
end Function;    
