-- Created on: 1993-11-10
-- Created by: Jean Marc LACHAUME
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Element from Geom2dHatch

uses
    Orientation from TopAbs,
    Curve from Geom2dAdaptor

is


    Create
    
    	returns Element from Geom2dHatch;

    Create (Other : Element from Geom2dHatch) 
    
    	---Purpose: Magic constructor.

	returns Element from Geom2dHatch ;
     

    Create (Curve       : Curve from Geom2dAdaptor ;
    	    Orientation : Orientation from TopAbs = TopAbs_FORWARD)
    
    	---Purpose: Creates an element.

	returns Element from Geom2dHatch ;


    Curve (me)
    
    	---Purpose: Returns the curve associated to the element.

    	---C++: return const &

        returns Curve from Geom2dAdaptor
        is static ;


    ChangeCurve (me : in out)
    
    	---Purpose: Returns the curve associated to the element.

    	---C++: return &

        returns Curve from Geom2dAdaptor
        is static ;


    Orientation (me : in out ; Orientation : Orientation from TopAbs)

    	---Purpose: Sets the orientation of the element.

    	is static ;


    Orientation (me)

    	---Purpose: Returns the orientation of the element.

    	returns Orientation from TopAbs
    	is static ;


fields

    myCurve       : Curve from Geom2dAdaptor ;
    myOrientation : Orientation from TopAbs ;

end Element from Geom2dHatch;
