-- Created on: 1993-05-05
-- Created by: Christian CAILLET
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Protocol  from IGESData  inherits  Protocol from Interface

    ---Purpose : Description of basic Protocol for IGES
    --           This comprises treatement of IGESModel and Recognition of
    --           Undefined-FreeFormat-Entity

uses OStream, Type, InterfaceModel, Check

is

    Create returns mutable Protocol from IGESData;

    NbResources (me) returns Integer;
    ---Purpose : Gives the count of Resource Protocol. Here, none

    Resource (me; num : Integer) returns Protocol from Interface;
    ---Purpose : Returns a Resource, given a rank. Here, none

    TypeNumber (me; atype : any Type) returns Integer;
    ---Purpose : Returns a Case Number, specific of each recognized Type
    --         Here, Undefined and Free Format Entities have the Number 1.

    	-- --    General Services (defined at Norm level)    -- --

    NewModel (me) returns mutable InterfaceModel;
    ---Purpose : Creates an empty Model for IGES Norm

    IsSuitableModel (me; model : InterfaceModel) returns Boolean;
    ---Purpose : Returns True if <model> is a Model of IGES Norm

    UnknownEntity (me) returns mutable Transient;
    ---Purpose : Creates a new Unknown Entity for IGES (UndefinedEntity)

    IsUnknownEntity (me; ent : Transient) returns Boolean;
    ---Purpose : Returns True if <ent> is an Unknown Entity for the Norm, i.e.
    --           Type UndefinedEntity, status Unknown

end Protocol;
