-- Created on: 1996-12-05
-- Created by: Odile Olivier
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class DimensionOwner from AIS inherits EntityOwner from SelectMgr

  ---Purpose: The owner is the entity which makes it possible to link
    -- the sensitive primitives and the reference shapes that
    -- you want to detect. It stocks the various pieces of
    -- information which make it possible to find objects. An
    -- owner has a priority which you can modulate, so as to
    -- make one entity more selectable than another. You
    -- might want to make edges more selectable than
    -- faces, for example. In that case, you could attribute sa
    -- higher priority to the one compared to the other. An
    -- edge, could have priority 5, for example, and a face,
    -- priority 4. The default priority is 5.

uses

    SelectableObject      from SelectMgr,
    PresentationManager   from PrsMgr,
    PresentationManager3d from PrsMgr,
    NameOfColor           from Quantity,
    DimensionDisplayMode  from AIS

is

    Create (theSelObject  : SelectableObject;
            theDisplayMode    : DimensionDisplayMode from AIS;
            thePriority   : Integer from Standard = 0)
    returns mutable DimensionOwner from AIS;
      ---Purpose:
      -- Initializes the dimension owner, theSO, and attributes it
      -- the priority, thePriority.

    SetDisplayMode (me : mutable; theMode : DimensionDisplayMode from AIS);

    DisplayMode (me)
    returns DimensionDisplayMode from AIS;

    HilightWithColor (me       : mutable;
                      thePM    : PresentationManager3d from PrsMgr;
                      theColor : NameOfColor from Quantity;
                      theMode  : Integer  from  Standard = 0)
    is redefined virtual;

    IsHilighted (me;
                 thePM   : PresentationManager from PrsMgr;
                 theMode : Integer  from  Standard  =0)
    returns Boolean from Standard is redefined virtual;
    ---Purpose: Returns true if an object with the selection mode
    -- aMode is highlighted in the presentation manager aPM.

    Hilight(me    : mutable;
            thePM   : PresentationManager from PrsMgr;
            theMode : Integer  from  Standard  =0) is redefined virtual;

    Unhilight(me    : mutable;
              thePM   : PresentationManager from PrsMgr;
              theMode : Integer  from  Standard  =0) is redefined virtual;
    ---Purpose: Removes highlighting from the selected part of dimension.
fields

    myDisplayMode : DimensionDisplayMode from AIS;

end DimensionOwner;
