-- Created on: 1992-08-26
-- Created by: Jean Louis FRENKEL
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Modified:	GG IMP020200 Add Transformation() method


class Presentation from Prs3d inherits Structure from Graphic3d

    	---Purpose: Defines a presentation object which can be displayed,
    	-- highlighted or erased.
    	-- The presentation object stores the results of the
    	-- presentation algorithms as defined in the StdPrs
    	-- classes and the Prs3d classes inheriting Prs3d_Root.
    	-- This presentation object is used to give display
    	-- attributes defined at this level to
    	-- ApplicationInteractiveServices classes at the level above.
      -- A presentation object is attached to a given Viewer.
        
uses
	Array2OfReal		from TColStd,
    DataStructureManager from Graphic3d,
    Structure            from Graphic3d,
    StructureManager     from Graphic3d,
    Group                from Graphic3d,
    Transformation       from Geom,
    NameOfColor          from Quantity,
    Length               from Quantity,
    ShadingAspect        from Prs3d
    
is

  Create (theStructManager : StructureManager from Graphic3d;
          theToInit        : Boolean          from Standard = Standard_True)
  ---Purpose: Constructs a presentation object
  -- if <Init> is false, no color initialization is done.
  returns Presentation from Prs3d;

  Create (theStructManager : StructureManager from Graphic3d;
          thePrs           : Presentation     from Prs3d)
  ---Purpose: Constructs a presentation object.
  returns Presentation from Prs3d;

    Compute(me : mutable; aProjector: DataStructureManager from Graphic3d)
    returns Structure from Graphic3d
    is redefined virtual;

	Compute ( me	: mutable;
		  aProjector	: DataStructureManager from Graphic3d;
		  AMatrix	: Array2OfReal from TColStd )
		returns Structure from Graphic3d is redefined virtual;
	---Level: Advanced
	---Purpose: Returns the new Structure defined for the new visualization
	---Category: Methods to modify the class definition

	Compute ( me	: mutable;
		  aProjector	: DataStructureManager from Graphic3d;
		  aStructure	: in out Structure from Graphic3d )
		is redefined virtual;
	---Level: Advanced
	---Purpose: Returns the new Structure defined for the new visualization
	---Category: Methods to modify the class definition

	Compute ( me	: mutable;
		  aProjector	: DataStructureManager from Graphic3d;
		  AMatrix	: Array2OfReal from TColStd;
		  aStructure	: in out Structure from Graphic3d )
		is redefined virtual;
	---Level: Advanced
	---Purpose: Returns the new Structure defined for the new visualization
	---Category: Methods to modify the class definition

---Category: Global modification methods.
    SetShadingAspect(me: mutable; aShadingAspect: ShadingAspect from Prs3d);

---Category: Transformation methods.
    Transform   (me: mutable; aTransformation: Transformation from Geom);
    Place       (me: mutable; X,Y,Z: Length from Quantity);

    Multiply    (me: mutable; aTransformation: Transformation from Geom); 
    Move        (me: mutable; X,Y,Z: Length from Quantity);
    Transformation   (me) returns Transformation from Geom;

    Connect(me: mutable; aPresentation: Presentation from Prs3d);
    
    Remove (me: mutable; aPresentation: Presentation from Prs3d);
    RemoveAll (me: mutable);

    CurrentGroup(me) returns Group from Graphic3d is static private;

friends

  class Root from Prs3d

end Presentation;
