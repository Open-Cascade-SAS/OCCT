-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SizeSelect from StepBasic   inherits SelectType from StepData

	-- <SizeSelect> is an EXPRESS Select Type construct translation.
	-- it gathers : MeasureWithUnit (Entity), PositiveLengthMeasure (Real)

uses

    SelectMember from StepData

is

    Create returns SizeSelect;
    ---Purpose : Returns a SizeSelect SelectType

    CaseNum (me; ent : Transient) returns Integer;
    ---Purpose: Recognizes a TrimmingSelect Kind Entity that is :
    --        1 -> SizeMember
    --        0 else (i.e. Real)

    NewMember (me) returns SelectMember  is redefined;
    ---Purpose : Returns a SizeMember (POSITIVE_LENGTH_MEASURE) as preferred

    CaseMem (me; ent : SelectMember) returns Integer  is redefined;
    ---Purpose : Recognizes a SelectMember as Real, named as PARAMETER_VALUE
    --            1 -> PositiveLengthMeasure i.e. Real
    --            0 else (i.e. Entity)
	
    SetRealValue (me : in out; aReal : Real from Standard);
	
    RealValue (me) returns Real;
    ---Purpose : returns Value as a Real (Null if another type)
	
end SizeSelect;

