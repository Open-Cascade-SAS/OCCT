-- Created on: 1997-08-13
-- Created by: Jean-Louis Frenkel
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DirectoryIterator from CDF

uses
    Directory from CDF,
    Document from CDM,
    ListIteratorOfListOfDocument from CDM
raises
    NoSuchObject from Standard

is

    Create
    returns DirectoryIterator from CDF;
    ---Purpose: creates an Iterator with the directory 
    --          of the current CDF.

    Create(aDirectory: Directory from CDF) 
    returns  DirectoryIterator from CDF;

    MoreDocument (me: in out) returns Boolean from Standard;
    ---Purpose : Returns True if there are more entries to return
    
    NextDocument (me: in out);
    ---Purpose : Go to the next entry
    --           (if there is not, Value will raise an exception)
    
    Document (me: in out) returns Document from CDM
    ---Purpose : Returns item value of current entry
    raises NoSuchObject  from Standard;

fields

    myIterator: ListIteratorOfListOfDocument from CDM;
end DirectoryIterator from CDF;
