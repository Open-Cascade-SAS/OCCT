-- Created on: 1992-09-28
-- Created by: Remi GILET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class MakeArcOfCircle from GC inherits Root from GC
    	---Purpose: Implements construction algorithms for an
    	-- arc of circle in 3D space. The result is a Geom_TrimmedCurve curve.
    	-- A MakeArcOfCircle object provides a framework for:
    	-- -   defining the construction of the arc of circle,
    	-- -   implementing the construction algorithm, and
    	-- -   consulting the results. In particular, the
    	--   Value function returns the constructed arc of circle.
        
uses Pnt          from gp,
     Circ         from gp,
     Dir          from gp,
     Ax1          from gp,
     Vec          from gp,
     Real         from Standard,
     TrimmedCurve from Geom

raises NotDone from StdFail

is

Create(Circ           : Circ    from gp       ;
       Alpha1, Alpha2 : Real    from Standard ;
       Sense          : Boolean from Standard ) returns MakeArcOfCircle;
    	---Purpose: Make an arc of circle (TrimmedCurve from Geom) from 
    	--          a circle between two angles Alpha1 and Alpha2 
    	--          given in radiians.

Create(Circ  : Circ    from gp       ;
       P     : Pnt     from gp       ;
       Alpha : Real    from Standard ;
       Sense : Boolean from Standard ) returns MakeArcOfCircle;
    	---Purpose: Make an arc of circle (TrimmedCurve from Geom) from 
    	--          a circle between point <P> and the angle Alpha 
    	--          given in radians.

Create(Circ  : Circ    from gp ;
       P1    : Pnt     from gp ;
       P2    : Pnt     from gp ;
       Sense : Boolean from Standard ) returns MakeArcOfCircle;
    	---Purpose: Make an arc of circle (TrimmedCurve from Geom) from 
    	--          a circle between two points P1 and P2.

Create(P1    : Pnt from gp ;
       P2    : Pnt from gp ;
       P3    : Pnt from gp ) 
    returns MakeArcOfCircle;
    	---Purpose: Make an arc of circle (TrimmedCurve from Geom) from 
    	--          three points P1,P2,P3 between two points P1 and P2.

Create(P1    : Pnt from gp ;
       V     : Vec from gp ;
       P2    : Pnt from gp )
    returns MakeArcOfCircle;
    	---Purpose: Make an arc of circle (TrimmedCurve from Geom) from 
    	--          two points P1,P2 and the tangente to the solution at 
    	--          the point P1.
    	-- The orientation of the arc is:
    	-- -   the sense determined by the order of the points P1, P3 and P2;
    	-- -   the sense defined by the vector V; or
    	-- -   for other syntaxes:
    	--   -   the sense of Circ if Sense is true, or
    	--   -   the opposite sense if Sense is false.
    	-- Note: Alpha1, Alpha2 and Alpha are angle values, given in radians.
    	-- Warning
    	-- If an error occurs (that is, when IsDone returns
    	-- false), the Status function returns:
    	-- -   gce_ConfusedPoints if:
    	--   -   any 2 of the 3 points P1, P2 and P3 are coincident, or
    	--   -   P1 and P2 are coincident; or
    	-- -   gce_IntersectionError if:
    	--   -   P1, P2 and P3 are collinear and not coincident, or
    	--   -   the vector defined by the points P1 and
    	--    P2 is collinear with the vector V.
    
Value(me) returns TrimmedCurve from Geom
    raises NotDone
    is static;
    ---Purpose: Returns the constructed arc of circle.
    -- Exceptions StdFail_NotDone if no arc of circle is constructed.
    ---C++: return const&

Operator(me) returns TrimmedCurve from Geom
    is static;
    ---C++: return const&
    ---C++: alias "Standard_EXPORT operator Handle_Geom_TrimmedCurve() const;"

fields

    TheArc : TrimmedCurve from Geom;
    --The solution from Geom.
    
end MakeArcOfCircle;
