-- Created by: NW,JPB,CAL
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


deferred class AspectLine from Aspect
	
inherits

	TShared

	---Purpose: This class allows the definition of a group
	--	    of attributes for the LINE primitive
	--	    The attributes are:
	--		* Colour
	--		* Type
	--		* Thickness
	--	    When any value of the group is modified
	--	    all graphic objects using the group are modified.

uses

	Color		from Quantity,

	TypeOfLine	from Aspect 

raises

	AspectLineDefinitionError	from Aspect

is

	Initialize;
	---Level: Public
	---Purpose: Initialise the constructor for Graphic3d_AspectLine3d.
	--
	-- Default values :
	--		Color = Quantity_NOC_YELLOW;
	--		Type  = Aspect_TOL_SOLID;
	--		Width = 1.0;
	--

	Initialize ( AColor	: Color from Quantity;
		     AType	: TypeOfLine from Aspect;
		     AWidth	: Real from Standard )
	---Level: Public
	---Purpose: Initialise the values for the
	--	    constructor of Graphic3d_AspectLine3d.
	--
	raises AspectLineDefinitionError from Aspect;
	-- if the width is a negative value.

	---------------------------------------------------
	-- Category: Methods to modify the class definition
	---------------------------------------------------

	SetColor ( me		: mutable;
		   AColor	: Color from Quantity );
	---Level: Public
	---Purpose: Modifies the colour of <me>.
	---Category: Methods to modify the class definition

	SetType ( me	: mutable;
		  AType	: TypeOfLine from Aspect );
	---Level: Public
	---Purpose: Modifies the type of <me>.
	---Category: Methods to modify the class definition

	SetWidth ( me		: mutable;
		   AWidth	: Real from Standard )
	---Level: Public
	---Purpose: Modifies the thickness of <me>.
	--  Category: Methods to modify the class definition
	--  Warning: Raises AspectLineDefinitionError if the
	--	    width is a negative value.
	raises AspectLineDefinitionError from Aspect;

	----------------------------
	-- Category: Inquire methods
	----------------------------

	Values ( me;
		 AColor	: out Color from Quantity;
		 AType	: out TypeOfLine from Aspect;
		 AWidth	: out Real from Standard );
	---Level: Public
	---Purpose: Returns the current values of the group <me>.
	---Category: Inquire methods

--

fields

--
-- Class	:	Aspect_AspectLine
--
-- Purpose	:	Declaration of variables specific to
--			drawing lines
--
-- Reminder	:	A line drawing context is defined by:
--			- the colour
--			- the type
--			- the thickness
--

	-- the colour
	MyColor	:	Color from Quantity;

	-- the type
	MyType	:	TypeOfLine from Aspect;

	-- the thickness
	MyWidth	:	Real from Standard;

end AspectLine;
