-- Created on: 1993-03-03
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Location from PTopLoc inherits Storable

	---Purpose: A Storable  composed local coordinate system. Made
	--          with local   coordinate systems raised   to  power
	--          elevation.
	--          
	--          A Location is either :
	--          
	--          * The Identity.
	--          
	--          * The product  of a Datum3D raised  to a power and
	--          an other Location called the next Location.

uses
    Datum3D      from PTopLoc,
    ItemLocation from PTopLoc

raises
    NoSuchObject from Standard

is
    Create returns Location from PTopLoc;
	---Purpose: Creates an Identity Location.
	---Level: Internal 
	
    Create(D : Datum3D from PTopLoc; 
    	   P : Integer from Standard;
	   N : Location from PTopLoc) 
    returns Location from  PTopLoc;
	---Purpose: Creates a location being the product.
	--          N * D ^ P
	---Level: Internal 
    
    IsIdentity(me) returns Boolean from Standard
	---Purpose: True when the location is an identity.
	---Level: Internal 
    is static;
    
    Datum3D(me) returns Datum3D from PTopLoc
	---Purpose: Returns the first Datum. An error is raised if the
	--          location is an identity.
	---Level: Internal 
    raises NoSuchObject from Standard
    is static;

    Power(me)   returns Integer from Standard
	---Purpose: Returns the power elevation of the first datum. An
	--          error is raised if the location is an identity.
	---Level: Internal 
    raises NoSuchObject from Standard
    is static;
    
    Next(me)    returns Location from PTopLoc
	---Purpose: Returns next Location. An error is raised if the
	--          location is an identity.
	---Level: Internal 
    raises NoSuchObject from Standard
    is static;
    
fields
    myData : ItemLocation from PTopLoc;

end Location;
