-- Created on: 1993-02-19
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Curve from BRepAdaptor inherits Curve from Adaptor3d

	---Purpose: The Curve from BRepAdaptor  allows to use  an Edge
	--          of the BRep topology like a 3D curve.
	--          
	--          It has the methods the class Curve from Adaptor3d.
	--          
	--          It  is created or  Initialized  with  an Edge.  It
	--          takes  into account local  coordinate systems.  If
	--          the Edge has a 3D curve it is  use  with priority.
	--          If the edge  has no 3D curve one  of the curves on
	--          surface is used. It is possible to enforce using a
	--          curve on surface by creating  or initialising with
	--          an Edge and a Face.

uses
    Edge               from TopoDS,
    Face               from TopoDS,
    CurveType          from GeomAbs,
    Shape              from GeomAbs,
    HCurve             from Adaptor3d,
    Curve              from GeomAdaptor,
    CurveOnSurface     from Adaptor3d,
    HCurveOnSurface    from Adaptor3d,
    BezierCurve        from Geom,
    BSplineCurve       from Geom,
    Array1OfReal       from TColStd,
    Trsf               from gp,
    Pnt                from gp,
    Vec                from gp,
    Circ               from gp,
    Elips              from gp,
    Hypr               from gp,
    Parab              from gp,
    Lin                from gp

raises
    NullObject   from Standard,
    DomainError  from Standard,
    OutOfRange   from Standard,
    NoSuchObject from Standard

is
    Create returns Curve from BRepAdaptor;
	---Purpose: Creates an undefined Curve with no Edge loaded.
	
    Create(E : Edge from TopoDS) returns Curve from BRepAdaptor;
	---Purpose: Creates a Curve  to  acces to the geometry of edge
	--          <E>.

    Create(E : Edge from TopoDS; F : Face from TopoDS) 
    returns Curve from BRepAdaptor;
	---Purpose: Creates a Curve to acces to  the geometry  of edge
	--          <E>.   The geometry  will   be  computed using the
	--          parametric curve of <E> on the face  <F>. An Error
	--          is  raised if  the edge does  not have a pcurve on
	--          the face.

    Initialize(me : in out; E : Edge from TopoDS)
	---Purpose: Sets  the Curve <me>  to acces to the  geometry of
	--          edge <E>. 
    is static;

    Initialize(me : in out; E : Edge from TopoDS; F : Face from TopoDS) 
	---Purpose: Sets the Curve <me>  to acces to  the  geometry of
	--          edge <E>.  The geometry will be computed using the
	--          parametric curve of <E>  on the face <F>. An Error
	--          is raised if the edge  does not  have a pcurve  on
	--          the face.
    raises DomainError from Standard
    is static;

    Trsf(me) returns Trsf from gp
	---Purpose: Returns the coordinate system of the curve.
	---C++: return const &
    is static;
    
    Is3DCurve(me) returns Boolean
	---Purpose: Returns True if the edge geometry is computed from
	--          a 3D curve.
    is static;
    
    IsCurveOnSurface(me) returns Boolean
	---Purpose: Returns True if the edge geometry is computed from
	--          a pcurve on a surface.
    is static;
    
    Curve(me) returns Curve from GeomAdaptor
	---Purpose: Returns the Curve of  the  edge.
	---C++: return const &
    is static;

    CurveOnSurface(me) returns CurveOnSurface from Adaptor3d
	---Purpose: Returns the CurveOnSurface of the edge.
	---C++: return const &
    is static;
    
    Edge(me) returns Edge from TopoDS
	---Purpose: Returns the edge.
	--          
	---C++: return const &
    is static;
    
    Tolerance(me) returns Real
	---Purpose: Returns the edge tolerance.
	--          
    is static;

    --
    --     Methods of  Curve  from GeomAdaptor.
    --     

   FirstParameter(me) returns Real
   is redefined static;

   LastParameter(me) returns Real
   is redefined static;     

   Continuity(me) returns Shape from GeomAbs
   is redefined static;

   NbIntervals(me; S : Shape from GeomAbs) returns Integer
	---Purpose: Returns  the number  of  intervals for  continuity
	--          <S>. May be one if Continuity(me) >= <S>
   is redefined static;

   Intervals(me; T : in out Array1OfReal from TColStd; 
    	          S : Shape from GeomAbs)
	---Purpose: Stores in <T> the  parameters bounding the intervals
	--          of continuity <S>.
	--          
	--          The array must provide  enough room to  accomodate
	--          for the parameters. i.e. T.Length() > NbIntervals()
   raises
    	OutOfRange from Standard 
   is redefined static;
    
   Trim(me; First, Last, Tol : Real) returns HCurve from Adaptor3d
	---Purpose: Returns    a  curve equivalent   of  <me>  between
	--          parameters <First>  and <Last>. <Tol>  is used  to
	--          test for 3d points confusion.
   raises
    	OutOfRange from Standard
	---Purpose: If <First> >= <Last> 
   is redefined static;
    
   IsClosed(me) returns Boolean
   is redefined static;
    
   IsPeriodic(me) returns Boolean
   is redefined static;

   Period(me) returns Real
    raises
    	DomainError from Standard -- if the curve is not periodic
    is redefined static;

    
   Value(me; U : Real) returns Pnt from gp
        --- Purpose : Computes the point of parameter U on the curve 
   is redefined static;

   D0 (me; U : Real; P : out Pnt from gp)
        --- Purpose : Computes the point of parameter U.
   is redefined static;

   D1 (me; U : Real; P : out Pnt from gp ; V : out Vec from gp)
        --- Purpose : Computes the point of parameter U on the curve
        --  with its first derivative.

     raises 
       DomainError from Standard
        --- Purpose : Raised if the continuity of the current interval
        --  is not C1.
   is redefined static;
    
   D2 (me; U : Real; P : out Pnt from gp; V1, V2 : out Vec from gp)
        --- Purpose :
        --  Returns the point P of parameter U, the first and second
        --  derivatives V1 and V2.
     raises 
       DomainError from Standard
        --- Purpose : Raised if the continuity of the current interval
        --  is not C2.
     is redefined static;

   D3 (me; U : Real; P : out Pnt from gp; V1, V2, V3 : out Vec from gp)
        --- Purpose :
        --  Returns the point P of parameter U, the first, the second 
        --  and the third derivative.
     raises 
    	DomainError from Standard
        --- Purpose : Raised if the continuity of the current interval
        --  is not C3.
    is redefined static;
        
   DN (me; U : Real; N : Integer)   returns Vec from gp
        --- Purpose :
        --  The returned vector gives the value of the derivative for the 
        --  order of derivation N.
     raises  
    	DomainError from Standard,
        --- Purpose : Raised if the continuity of the current interval
        --  is not CN.
        OutOfRange from Standard
        --- Purpose : Raised if N < 1.            
    is redefined static;


   Resolution(me; R3d :Real) returns Real
        ---Purpose : returns the parametric resolution
   is redefined static;   
   

   GetType(me) returns CurveType from GeomAbs
   is redefined static;

   Line(me) returns Lin from gp
    raises NoSuchObject from Standard
   is redefined static;
   
   Circle(me) returns Circ from gp
    raises NoSuchObject from Standard
   is redefined static;

   Ellipse(me) returns Elips from gp
    raises NoSuchObject from Standard
   is redefined static;

   Hyperbola(me) returns  Hypr from gp
    raises NoSuchObject from Standard
   is redefined static;

   Parabola(me) returns Parab from gp
    raises NoSuchObject from Standard
   is redefined static;


   Degree(me) returns Integer
    raises NoSuchObject from Standard
   is redefined static;

   IsRational(me) returns Boolean
     raises 
    	NoSuchObject from Standard
   is redefined static;

   NbPoles(me) returns Integer
    raises NoSuchObject from Standard
   is redefined static;
    
   NbKnots(me) returns Integer
     raises 
    	NoSuchObject from Standard
   is redefined static;


   Bezier(me) returns BezierCurve from Geom
    	---Purpose: 
        --  Warning : 
    	--         This  will    make a copy of the Bezier Curve
    	--         since it applies to it myTsrf . Be carefull when
    	--         using this method
   raises 
    	NoSuchObject from Standard
   is redefined static;
   
   BSpline(me) returns BSplineCurve from Geom
    	---Purpose: 
    --  Warning : 
    	--         This will   make a copy of the BSpline Curve
    	--         since it applies to it myTsrf . Be carefull when
    	--         using this method

   raises 
    	NoSuchObject from Standard
   is redefined static;

fields

   myTrsf    : Trsf              from gp;
   myCurve   : Curve             from GeomAdaptor;
   myConSurf : HCurveOnSurface   from Adaptor3d;
   myEdge    : Edge              from TopoDS;

end Curve;
