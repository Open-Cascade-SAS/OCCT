-- Created on: 1990-12-19
-- Created by: Christophe MARION
-- Copyright (c) 1990-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package TopLoc 

    ---Level : Public. 
    --  All methods of all  classes will be public.

    ---Purpose: The TopLoc package gives ressources to handle 3D local
    --          coordinate systems called Locations.
    --          
    --          A Location  is a composition of  elementary coordinate
    --          systems,  each one is  called a  Datum.   The Location
    --          keeps track of  this composition.
    --          
    
uses
    Standard,
    MMgt,
    TCollection,
    gp

is
    pointer TrsfPtr to Trsf from gp;
    class Datum3D;
    
    private class ItemLocation;
	
    private class SListOfItemLocation;
    private class SListNodeOfItemLocation;
    
    class Location;

    class MapLocationHasher instantiates
    	  MapHasher from TCollection(Location from TopLoc); 
	  
    class MapOfLocation instantiates
    	  Map from TCollection(Location          from TopLoc,
	    	    	       MapLocationHasher from TopLoc);
    	
    class IndexedMapOfLocation instantiates
    	  IndexedMap from TCollection(Location          from TopLoc,
	    	 		      MapLocationHasher from TopLoc);
    	
end TopLoc;




