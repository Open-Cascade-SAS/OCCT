-- Created on: 1993-03-24
-- Created by: Philippe DAUTRY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class CartesianPoint from Geom2d inherits Point from Geom2d

        --- Purpose : Describes a point in 2D space. A
    	-- Geom2d_CartesianPoint is defined by a gp_Pnt2d
    	-- point, with its two Cartesian coordinates X and Y.
     


uses Ax2d       from gp, 
     Pnt2d      from gp,
     Trsf2d     from gp,
     Vec2d      from gp,
     Geometry   from Geom2d

is

  Create (P : Pnt2d)   returns mutable CartesianPoint;
        --- Purpose : Returns a persistent copy of P.


  Create (X, Y : Real)   returns mutable CartesianPoint;



  SetCoord (me : mutable; X, Y : Real);
        --- Purpose : Set <me> to X, Y coordinates.


  SetPnt2d (me : mutable; P : Pnt2d);
        --- Purpose : Set <me> to P.X(), P.Y() coordinates.


  SetX (me : mutable; X : Real);
        --- Purpose : Changes the X coordinate of me.


  SetY (me : mutable; Y : Real);
        --- Purpose : Changes the Y coordinate of me.

 
  Coord (me; X, Y : out Real);
        --- Purpose : Returns the coordinates of <me>.


  Pnt2d (me)  returns Pnt2d;
        --- Purpose :
        --  Returns a non persistent cartesian point with
        --  the same coordinates as <me>.
    	-- -C++: return const&


  X (me)  returns Real;
        --- Purpose : Returns the X coordinate of <me>.


  Y (me)  returns Real;
        --- Purpose : Returns the Y coordinate of <me>.



  Transform (me : mutable; T : Trsf2d);



  Copy (me)  returns mutable like me;
     
fields

  gpPnt2d : Pnt2d;

end;
