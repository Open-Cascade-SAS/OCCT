-- Created on: 1996-10-23
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class FFDumper from TopOpeBRep inherits TShared from MMgt

uses

    DataMapOfShapeInteger from TopTools,
    PFacesFiller from TopOpeBRep,
    LineInter from TopOpeBRep, 
    VPointInter from TopOpeBRep,
    VPointInterIterator from TopOpeBRep,
    Kind from TopOpeBRepDS,    
    Shape from TopoDS,
    Face from TopoDS
    
is 

    Create(PFF:PFacesFiller) returns mutable FFDumper from  TopOpeBRep; 
    Init(me:mutable;PFF:PFacesFiller); 
    DumpLine(me:mutable;I:Integer);
    DumpLine(me:mutable;L:LineInter);
    DumpVP(me:mutable;VP:VPointInter);
    DumpVP(me:mutable;VP:VPointInter;ISI:Integer); 
    ExploreIndex(me;S:Shape;ISI:Integer) returns Integer; 
    DumpDSP(me;VP:VPointInter;GK:Kind;G:Integer;newinDS:Boolean);
    PFacesFillerDummy(me) returns PFacesFiller;

fields

    myPFF:PFacesFiller from TopOpeBRep;
    myF1,myF2:Face from TopoDS;
    myEM1,myEM2:DataMapOfShapeInteger from TopTools; 
    myEn1,myEn2:Integer;
    myLineIndex : Integer;

end FFDumper from TopOpeBRep;
