-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class StyledItem from StepVisual 

inherits RepresentationItem from StepRepr

uses

	HArray1OfPresentationStyleAssignment from StepVisual, 
	PresentationStyleAssignment from StepVisual, 
	HAsciiString from TCollection
is

	Create returns StyledItem;
	---Purpose: Returns a StyledItem


	Init (me : mutable;
	      aName : HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      aName : HAsciiString from TCollection;
	      aStyles : HArray1OfPresentationStyleAssignment from StepVisual;
	      aItem : RepresentationItem from StepRepr) is virtual;

	-- Specific Methods for Field Data Access --

	SetStyles(me : mutable; aStyles : HArray1OfPresentationStyleAssignment);
	Styles (me) returns HArray1OfPresentationStyleAssignment;
	StylesValue (me; num : Integer) returns PresentationStyleAssignment;
	NbStyles (me) returns Integer;
	SetItem(me : mutable; aItem : RepresentationItem);
	Item (me) returns RepresentationItem;

fields

	styles : HArray1OfPresentationStyleAssignment from StepVisual;
	item : RepresentationItem from StepRepr;

end StyledItem;
