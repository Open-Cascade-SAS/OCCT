-- Created on: 1993-03-02
-- Created by: Philippe DAUTRY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ConicalSurface from PGeom inherits ElementarySurface from PGeom

        ---Purpose : This class defines the infinite conical surface .
        -- 
	---See Also : ConicalSurface from Geom.

uses Ax3      from gp

is


  Create returns mutable ConicalSurface from PGeom;
	---Purpose: Creates a ConicalSurface with default values.
    	---Level: Internal 


  Create (aPosition  : Ax3 from gp;
    	  aRadius    : Real from Standard;
    	  aSemiAngle : Real from Standard)
     returns mutable ConicalSurface from PGeom;
	---Purpose: Creates a ConicalSurface with these values.
    	---Level: Internal 


  Radius (me: mutable; aRadius: Real from Standard);
        ---Purpose : Set the field radius with <aRadius>.
    	---Level: Internal 


  Radius (me) returns Real from Standard;
        ---Purpose : Returns the value of the field radius.
    	---Level: Internal 
     
     
  SemiAngle (me : mutable; aSemiAngle : Real from Standard);
        ---Purpose : Set the value of the field semiAngle with <aSemiAngle>.
    	---Level: Internal 


  SemiAngle (me) returns Real from Standard;
        --- Purpose : Returns the value of the field semiAngle.
    	---Level: Internal 


fields

  radius    : Real from Standard;
  semiAngle : Real from Standard;

end;
