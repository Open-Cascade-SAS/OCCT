-- Created on: 2008-05-08
-- Created by: Vladislav ROMASHKO
-- Copyright (c) 2008-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class ColorDS from Voxel inherits DS from Voxel

    ---Purpose: A 3D voxel model keeping 4 bits for each voxel (one of 16 colors).

is

    Create
    ---Purpose: An empty constructor.
    returns ColorDS from Voxel;

    Create(x     : Real    from Standard;
    	   y     : Real    from Standard;
    	   z     : Real    from Standard;
    	   x_len : Real    from Standard;
    	   y_len : Real    from Standard;
    	   z_len : Real    from Standard;
	   nb_x  : Integer from Standard;
	   nb_y  : Integer from Standard;
	   nb_z  : Integer from Standard)
    ---Purpose: A constructor initializing the voxel model.
    --          (x, y, z) - the start point of the box.
    --          (x_len, y_len, z_len) - lengths in x, y and z directions along axes of a co-ordinate system.
    --          (nb_x, nb_y, nb_z) - number of splits (voxels) along x, y and z directions.
    returns ColorDS from Voxel;

    Init(me : in out;
    	 x     : Real    from Standard;
    	 y     : Real    from Standard;
    	 z     : Real    from Standard;
    	 x_len : Real    from Standard;
    	 y_len : Real    from Standard;
    	 z_len : Real    from Standard;
	 nb_x  : Integer from Standard;
	 nb_y  : Integer from Standard;
	 nb_z  : Integer from Standard)
    ---Purpose: Initialization of the voxel model.
    --          (x, y, z) - the start point of the box.
    --          (x_len, y_len, z_len) - lengths in x, y and z directions along axes of a co-ordinate system.
    --          (nb_x, nb_y, nb_z) - number of splits (voxels) along x, y and z directions.
    is redefined virtual;

    Destroy(me : in out);
    ---C++: alias ~
    ---Purpose: A destructor of the voxel model.

    SetZero(me : in out);
    ---Purpose: The method sets all values equal to 0 (false) and
    --          releases the memory.

    Set(me   : in out;
    	ix   : Integer from Standard;
    	iy   : Integer from Standard;
    	iz   : Integer from Standard;
	data : Byte    from Standard);
    ---Purpose: Defines a value for voxel with co-ordinates (ix, iy, iz).
    --          Only the first four bits are used!
    --          Initial state of the model is so that all voxels have value 0x0000,
    --          and this data doesn't occupy memory.
    --          Memory for data is allocating during setting non-zero values (0x0101, for example).

    Get(me;
    	ix : Integer from Standard;
    	iy : Integer from Standard;
    	iz : Integer from Standard)
    ---Purpose: Returns the value of voxel with co-ordinates (ix, iy, iz).
    returns Byte from Standard;

end ColorDS;
