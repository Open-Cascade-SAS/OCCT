-- File:	BOPTools_InterferencePool.cdl
-- Created:	Fri Jan 26 12:00:38 2001
-- Author:	Peter KURNEV
--		<pkv@irinox>
---Copyright:	 Matra Datavision 2001


class InterferencePool from BOPTools 

	---Purpose:  
    	--  Class for storing information about  
    	--- results of all interferences for all shapes 

uses 
    ShapesDataStructure  from BooleanOperations, 
    PShapesDataStructure from BooleanOperations,  
    KindOfInterference   from BooleanOperations, 
    
    CArray1OfInterferenceLine from BOPTools, 
    CArray1OfSSInterference   from BOPTools,
    CArray1OfESInterference   from BOPTools,
    CArray1OfVSInterference   from BOPTools, 
    CArray1OfEEInterference   from BOPTools, 
    CArray1OfVEInterference   from BOPTools, 
    CArray1OfVVInterference   from BOPTools, 
    PShapeShapeInterference   from BOPTools 
is 
    Create  
    	returns InterferencePool from BOPTools ; 
    	---Purpose:  
    	--- Empty constructor 
    	---
    Create  (aDS:ShapesDataStructure from BooleanOperations)
    	returns InterferencePool from BOPTools ;  
    	---Purpose:   
    	--- Constructor 
    	---
    SetDS  (me:out;aDS:ShapesDataStructure from BooleanOperations); 
    	---Purpose:  
    	--- Modifier  
    	---
    DS(me) 
    	returns  PShapesDataStructure from BooleanOperations; 
    	---Purpose:  
    	--- Selector  
    	---
    HasInterference  (me; 
    	     anInd  :Integer from Standard) 
	returns Boolean from Standard;  
    	---Purpose: 
    	--- Returns  TRUE if the shape with DS_index  <anInd> 
    	--- has at least one  interference with non-empty result            
    	---
    IsComputed     (me;   
    	     anInd1  :  Integer from Standard;
    	     anInd2  :  Integer from Standard) 
	returns Boolean from Standard;  
    	---Purpose: 
    	--- Returns  TRUE if the interference between shapes  
    	--- <anInd1> and <anInd2> has already been computed.           
    	---
    SortTypes      (me;   
    	    	anInd1:in out Integer from Standard; 
                anInd2:in out Integer from Standard); 
    	---Purpose: 
    	--- Sorts types of shapes <anInd1> and <anInd2> in increasing order 
    	---
    InterferenceType  (me;   
    	    	anInd1: Integer from Standard; 
    	    	anInd2: Integer from Standard) 
    	returns KindOfInterference from BooleanOperations;  
    	---Purpose: 
    	--- Gets the type of interference in accordance with the types of  
    	--- shapes  <anInd1> and <anInd2>
    	---
    AddInterference   (me:out;   
    	    	anInd1:  Integer from Standard;
    	    	anInd2:  Integer from Standard; 
                aType:   KindOfInterference from BooleanOperations; 
	    	anIndex: Integer from Standard);  
    	---Purpose: 
    	--- Adds the info about interference in InterferenceLine-s for  
    	--- shapes  <anInd1> and <anInd2>
    	---
    InterferenceTable (me) 
    	returns  CArray1OfInterferenceLine from BOPTools; 
    	---C++:  return  const& 
    	---Purpose: 
    	--- Returns the reference to complete array of interference line-s 
    	---
    SSInterferences (me:out)  
	returns CArray1OfSSInterference   from BOPTools; 
    	---C++:  return  & 
    	---Purpose: 
    	--- Returns the reference to array Of F/F interferences 
    	---
    ESInterferences (me:out)  
	returns CArray1OfESInterference   from BOPTools; 
    	---C++:  return  & 
    	---Purpose: 
    	--- Returns the reference to array Of E/F interferences 
    	---
    VSInterferences (me:out)  
	returns CArray1OfVSInterference   from BOPTools; 
    	---C++:  return  &
    	---Purpose: 
    	--- Returns the reference to array Of V/F interferences 
    	---
    EEInterferences (me:out)  
	returns CArray1OfEEInterference   from BOPTools; 
    	---C++:  return  &  
    	---Purpose: 
    	--- Returns the reference to arrray Of E/E interferences 
    	---
    VEInterferences (me:out)  
	returns CArray1OfVEInterference   from BOPTools; 
    	---C++:  return  &  	 	
    	---Purpose: 
    	--- Returns the reference to arrray Of  V/E interferences 
    	---
    VVInterferences (me:out)  
	returns CArray1OfVVInterference   from BOPTools; 
    	---C++:  return  &  	 	
    	---Purpose: 
    	--- Returns the reference to arrray Of  V/V interferences 
    	---
    -------------- 
    SSInterfs (me)  
	returns CArray1OfSSInterference   from BOPTools; 
    	---C++:  return const & 
     
    ESInterfs (me)  
	returns CArray1OfESInterference   from BOPTools; 
    	---C++:  return const & 
     
    VSInterfs (me)  
	returns CArray1OfVSInterference   from BOPTools; 
    	---C++:  return const &
     
    EEInterfs (me)  
	returns CArray1OfEEInterference   from BOPTools; 
    	---C++:  return const &  
	    
    VEInterfs (me)  
	returns CArray1OfVEInterference   from BOPTools; 
    	---C++:  return const &  	 	
		 
    VVInterfs (me)  
	returns CArray1OfVVInterference   from BOPTools; 
    	---C++:  return const & 
     

    GetInterference (me; 
    	    anIndex:  Integer from Standard; 
            aType  :  KindOfInterference from BooleanOperations) 
	returns PShapeShapeInterference from BOPTools; 


fields 
 
    myDS               :  PShapesDataStructure from BooleanOperations;  
    myNbSourceShapes   :  Integer  from  Standard;  
    
    myInterferenceTable:  CArray1OfInterferenceLine from BOPTools; 
    mySSInterferences  :  CArray1OfSSInterference   from BOPTools;
    myESInterferences  :  CArray1OfESInterference   from BOPTools;
    myVSInterferences  :  CArray1OfVSInterference   from BOPTools;
    myEEInterferences  :  CArray1OfEEInterference   from BOPTools;
    myVEInterferences  :  CArray1OfVEInterference   from BOPTools;
    myVVInterferences  :  CArray1OfVVInterference   from BOPTools;

end InterferencePool;
