-- Created on: 1993-01-13
-- Created by: CKY / Contract Toubro-Larsen ( Deepak PRABHU )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MacroDef from IGESDefs  inherits IGESEntity

        ---Purpose: defines IGES Macro Definition Entity, Type <306> Form <0>
        --          in package IGESDefs
        --          This Class specifies the action of a specific MACRO.
        --          After specification MACRO can be used as necessary
        --          by means of MACRO class instance entity.

uses

        HAsciiString          from TCollection,
        HArray1OfHAsciiString from Interface

raises OutOfRange

is

        Create returns mutable MacroDef;

        -- Specific methods for the entity

        Init (me             : mutable;
              macro          : HAsciiString;
              entityTypeID   : Integer;
              langStatements : HArray1OfHAsciiString;
              endMacro       : HAsciiString);
        ---Purpose : This method is used to set the fields of the class
        --           MacroDef
        --       - macro          : MACRO
        --       - entityTypeID   : Entity Type ID
        --       - langStatements : Language Statements
        --       - endMacro       : END MACRO

        NbStatements(me) returns Integer;
        ---Purpose : returns the number of language statements

        MACRO(me) returns HAsciiString from TCollection;
        ---Purpose : returns the MACRO(Literal)

        EntityTypeID(me) returns Integer;
        ---Purpose : returns the Entity Type ID

        LanguageStatement(me ; StatNum : Integer) 
        returns HAsciiString from TCollection
        raises OutOfRange;
        -- returns the StatNum'th statement
        -- raises exception if StatNum <= 0 or StatNum > NbStatements()

        ENDMACRO(me) returns HAsciiString from TCollection;
        ---Purpose : returns the ENDM(Literal)

fields

--
--  Class    : IGESDefs_MacroDef
--
--  Purpose  : Declaration of variables specific to MacroDef
--
--  Reminder : An MacroDef Entity specifies the action of a
--             specific MACRO. It consists of only language
--             statements in the parameter data.

        theMACRO          : HAsciiString;
        theEntityTypeID   : Integer;
        theLangStatements : HArray1OfHAsciiString;
        theENDMACRO       : HAsciiString;

end MacroDef;
