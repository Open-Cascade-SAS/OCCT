-- Created on: 1998-06-03
-- Created by: data exchange team
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Surface from ShapeCustom 

    ---Purpose: Converts a surface to the analitical form with given 
    --          precision. Conversion is done only the surface is bspline
    --          of bezier and this can be approximed by some analytical
    --          surface with that precision.

uses
    Surface from Geom

is

    Create returns Surface from ShapeCustom;
    
    Create (S: Surface from Geom) returns Surface from ShapeCustom;

    Init (me: in out; S: Surface from Geom);

    Gap (me) returns Real;
    ---C++: inline
    	---Purpose: Returns maximal deviation of converted surface from the original 
	--          one computed by last call to ConvertToAnalytical

    ConvertToAnalytical (me: in out; tol: Real;
    	    	    	    	     substitute: Boolean)
    returns Surface from Geom;
    	---Purpose: Tries to convert the Surface to an Analytic form
    	--          Returns the result
    	--          Works only if the Surface is BSpline or Bezier.
    	--          Else, or in case of failure, returns a Null Handle
    	--
    	--          If <substitute> is True, the new surface replaces the actual
    	--          one in <me>
    	--
    	--          It works by analysing the case which can apply, creating the
    	--          corresponding analytic surface, then checking coincidence
    	--  Warning: Parameter laws are not kept, hence PCurves should be redone
	
    ConvertToPeriodic (me: in out; substitute: Boolean; preci: Real = -1)
    returns Surface from Geom;
        ---Purpose: Tries to convert the Surface to the Periodic form
    	--          Returns the resulting surface
    	--          Works only if the Surface is BSpline and is closed with 
        --          Precision::Confusion()
    	--          Else, or in case of failure, returns a Null Handle
fields

    mySurf: Surface from Geom;
    myGap : Real; -- maximal deviation of converted surface from original one

end Surface;
