-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class VertexLoop from StepShape 

inherits Loop from StepShape 

uses

	Vertex from StepShape, 
	HAsciiString from TCollection
is

	Create returns VertexLoop;
	---Purpose: Returns a VertexLoop


	Init (me : mutable;
	      aName : HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      aName : HAsciiString from TCollection;
	      aLoopVertex : Vertex from StepShape) is virtual;

	-- Specific Methods for Field Data Access --

	SetLoopVertex(me : mutable; aLoopVertex : Vertex);
	LoopVertex (me) returns Vertex;

fields

	loopVertex : Vertex from StepShape;

end VertexLoop;
