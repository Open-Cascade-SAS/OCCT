-- Created on: 1995-03-09
-- Created by: Laurent PAINNOT
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class GCurve from BRep inherits CurveRepresentation from BRep

	---Purpose: Root   class    for    the    geometric     curves
	--          representation. Contains a range.

uses

    Location from TopLoc,
    Pnt      from gp

is

    Initialize(L : Location from TopLoc; First, Last : Real);

    SetRange(me : mutable; First, Last : Real)
	---C++: inline
    is static;
    
    Range(me; First, Last : out Real)
	---C++: inline
    is static;
    
    First(me) returns Real
	---C++: inline
    is static;

    Last(me) returns Real
	---C++: inline
    is static;

    First(me : mutable; F : Real)
	---C++: inline
    is static;

    Last(me : mutable; L : Real)
	---C++: inline
    is static;


    D0(me; U : Real; P : out Pnt from gp)
	---Purpose: Computes the point at parameter U.
    is deferred;
    

    Update(me : mutable)
	---Purpose: Recomputes any derived data after a modification.
	--          This is called when the range is modified.
    is virtual;

fields
    myFirst    : Real;
    myLast     : Real;

end GCurve;
