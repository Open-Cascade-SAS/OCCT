-- Created on: 1997-02-12
-- Created by: Alexander BRIVIN
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PointLight from Vrml 

	---Purpose:defines a point  light node of VRML specifying
	--         properties of lights. 
    	--  This  node  defines  a  point  light  source   at  a  fixed  3D  location
    	--  A  point  source  illuminates equally  in  all  directions;   
    	--  that  is  omni-directional.
    	--  Color is  written  as  an  RGB  triple.
    	--  Light intensity must be in the range 0.0 to 1.0, inclusive.  

uses
 
    Color   from Quantity, 
    Vec     from gp

is
                                                    --  defaults  :
    Create returns PointLight from Vrml; 
    	    	    	    	    	    	    --  myOnOff(Standard_TRUE)
 						    --  myIntensity(1)
						    --  myColor(1 1 1)
						    --  myLocation(0 0 1)

    Create  (  aOnOff     :   Boolean from  Standard; 
    	       aIntensity :   Real    from  Standard; 
    	       aColor     :   Color   from  Quantity; 
    	       aLocation  :   Vec     from  gp ) 
    	returns PointLight from Vrml; 
     
    SetOnOff ( me : in out;  aOnOff : Boolean from  Standard );
    OnOff ( me )  returns Boolean  from  Standard;

    SetIntensity ( me : in out;  aIntensity : Real from  Standard );
    Intensity ( me )  returns Real  from  Standard;

    SetColor ( me : in out;  aColor :  Color   from  Quantity );
    Color ( me )  returns  Color   from  Quantity;

    SetLocation ( me : in out;  aLocation : Vec  from  gp );
    Location ( me )  returns Vec  from  gp;

    Print  ( me;  anOStream: in out OStream from Standard) returns OStream from Standard;
    ---C++:  return  & 

fields
 
    myOnOff     :   Boolean from  Standard; -- Whether light is on
    myIntensity :   Real    from  Standard; -- Source intensity (0 to 1)
    myColor     :   Color   from  Quantity; -- RGB source color
    myLocation  :   Vec     from  gp;       -- Illumination Location vector

end PointLight;

