-- File:        SiUnitAndLengthUnit.cdl
-- Created:     Mon Dec  4 12:02:36 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWSiUnitAndLengthUnit from RWStepBasic

	---Purpose : Read & Write Module for SiUnitAndLengthUnit

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     SiUnitAndLengthUnit from StepBasic

is

	Create returns RWSiUnitAndLengthUnit;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable SiUnitAndLengthUnit from StepBasic);

	WriteStep (me; SW : in out StepWriter; ent : SiUnitAndLengthUnit from StepBasic);

end RWSiUnitAndLengthUnit;
