-- Created on: 1999-03-24
-- Created by: data exchange team
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class AssemblyComponent from STEPSelections inherits TShared from MMgt

	---Purpose: 

uses
    
    ShapeDefinitionRepresentation from StepShape,
    HSequenceOfAssemblyLink from STEPSelections

is
    
    Create returns AssemblyComponent from STEPSelections;
    
    Create (sdr : ShapeDefinitionRepresentation from StepShape;
    	    list: HSequenceOfAssemblyLink from STEPSelections)
    returns AssemblyComponent from STEPSelections;
    
    --Methods for getting and obtaining fields
    
    GetSDR(me) returns ShapeDefinitionRepresentation from StepShape;
    	---Purpose:
	---C++: inline
    
    GetList(me) returns HSequenceOfAssemblyLink from STEPSelections;
    	---Purpose:
	---C++: inline
    
    SetSDR(me : mutable; sdr: ShapeDefinitionRepresentation from StepShape);
    	---Purpose:
	---C++: inline
    
    SetList(me : mutable; list: HSequenceOfAssemblyLink from STEPSelections);
    	---Purpose:
	---C++: inline

fields

    mySDR : ShapeDefinitionRepresentation from StepShape;
    myList: HSequenceOfAssemblyLink from STEPSelections;

end AssemblyComponent;
