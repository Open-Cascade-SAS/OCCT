-- File:        ProductDefinitionContext.cdl
-- Created:     Mon Dec  4 12:02:29 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWProductDefinitionContext from RWStepBasic

	---Purpose : Read & Write Module for ProductDefinitionContext

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     ProductDefinitionContext from StepBasic,
     EntityIterator from Interface

is

	Create returns RWProductDefinitionContext;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable ProductDefinitionContext from StepBasic);

	WriteStep (me; SW : in out StepWriter; ent : ProductDefinitionContext from StepBasic);

	Share(me; ent : ProductDefinitionContext from StepBasic; iter : in out EntityIterator);

end RWProductDefinitionContext;
