-- Created on: 1993-11-26
-- Created by: Modelistation
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class ALineToWLine from IntPatch

uses 
    WLine from IntPatch,
    ALine from IntPatch,
    Quadric from IntSurf

is 

    Create(Quad1 : Quadric from IntSurf;
    	   Quad2 : Quadric from IntSurf)
    
    	returns ALineToWLine from IntPatch;
	
    Create(Quad1       : Quadric from IntSurf;
           Quad2       : Quadric from IntSurf;
           Deflection  : Real from Standard;
    	   PasMaxUV    : Real from Standard;
           NbMaxPoints : Integer from Standard) 
    
    	returns ALineToWLine from IntPatch;
	
	
    SetTolParam(me:out; 
    	    aT:Real from Standard); 
	 
    TolParam(me) 
    	returns Real from Standard; 
	 
    SetTolOpenDomain(me:out; 
    	    aT:Real from Standard); 
	 
    TolOpenDomain(me) 
    	returns Real from Standard; 
	 
    SetTolTransition(me:out; 
    	    aT:Real from Standard); 
	 
    TolTransition(me) 
    	returns Real from Standard;  

    SetTol3D(me:out; 
    	    aT:Real from Standard); 
	 
    Tol3D(me) 
    	returns Real from Standard;  
     
    SetConstantParameter(me);
    
    SetUniformAbscissa(me);
    
    SetUniformDeflection(me);
    
    MakeWLine(me; aline: ALine from IntPatch)
    
    	returns WLine from IntPatch;
	
    MakeWLine(me; aline: ALine from IntPatch; paraminf,paramsup: Real from Standard)
    	returns WLine from IntPatch; 
    
fields
    quad1         : Quadric from IntSurf;
    quad2         : Quadric from IntSurf;
    deflectionmax : Real    from Standard;
    pasuvmax      : Real    from Standard;
    nbpointsmax   : Integer from Standard;
    type          : Integer from Standard; -- 0: Constant Parameter
                                           -- 1: Uniform Abscissa
                                           -- 2: Uniform Deflection
    myTolParam      : Real from Standard; 
    myTolOpenDomain : Real from Standard; 
    myTolTransition : Real from Standard; 
    myTol3D         : Real from Standard;        

end;
