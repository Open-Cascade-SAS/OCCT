-- Created on: 2001-04-24
-- Created by: Christian CAILLET
-- Copyright (c) 2001-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class CompoundRepresentationItem  from StepRepr
  inherits RepresentationItem  from StepRepr

    ---Purpose : Added for Dimensional Tolerances

uses
    HAsciiString from TCollection,
    HArray1OfRepresentationItem from StepRepr

is

    Create returns CompoundRepresentationItem;

    Init (me : mutable;
             aName : HAsciiString from TCollection;
	     item_element : HArray1OfRepresentationItem from StepRepr);

    ItemElement (me) returns HArray1OfRepresentationItem from StepRepr;
    NbItemElement (me) returns Integer;
    SetItemElement (me : mutable; item_element : HArray1OfRepresentationItem from StepRepr);
    ItemElementValue (me; num : Integer) returns RepresentationItem;
    SetItemElementValue (me : mutable; num : Integer;
    	anelement : RepresentationItem);

fields

    theItemElement : HArray1OfRepresentationItem from StepRepr;

end CompoundRepresentationItem;
