-- File:	IGESSolid_ToolSolidInstance.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolSolidInstance  from IGESSolid

    ---Purpose : Tool to work on a SolidInstance. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses SolidInstance from IGESSolid,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolSolidInstance;
    ---Purpose : Returns a ToolSolidInstance, ready to work


    ReadOwnParams (me; ent : mutable SolidInstance;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : SolidInstance;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : SolidInstance;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a SolidInstance <ent>, from
    --           its specific (own) parameters

    DirChecker (me; ent : SolidInstance) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : SolidInstance;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : SolidInstance; entto : mutable SolidInstance;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : SolidInstance;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolSolidInstance;
