-- Created on: 1992-10-14
-- Created by: Gilles DEBARBOUILLE
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Edge from MAT 

	---Purpose: 

inherits

    TShared from MMgt
    
uses

    Bisector from MAT,
    ListOfEdge from MAT

--raises

is

    Create returns mutable Edge from MAT;
    
    EdgeNumber(me : mutable ; anumber : Integer)

    is static;
    
    FirstBisector(me : mutable ; abisector : any Bisector from MAT)

    is static;
    
    SecondBisector(me : mutable ; abisector : any Bisector from MAT)

    is static;
    
    Distance(me : mutable ; adistance : Real)

    is static;
    
    IntersectionPoint(me : mutable ; apoint : Integer)

    is static;

    EdgeNumber(me) returns Integer

    is static;
    
    FirstBisector(me) returns any Bisector from MAT

    is static;
    
    SecondBisector(me) returns any Bisector from MAT

    is static;
    
    Distance(me) returns Real

    is static;
    
    IntersectionPoint(me) returns Integer

    is static;

    Dump(me ; ashift , alevel : Integer)
    
    is static;
    
fields

    theedgenumber        : Integer;
    thefirstbisector     : Bisector from MAT;
    thesecondbisector    : Bisector from MAT;
    thedistance          : Real;
    theintersectionpoint : Integer;

end Edge;
