-- Created on: 1992-10-22
-- Created by: Gilles DEBARBOUILLE
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Material from Materials 

	---Purpose: This  class describes  the facilities available to
	--          create and manipulate materials.

inherits

    FuzzyInstance from Materials
    
uses

    HAsciiString from TCollection,
    AsciiString from TCollection

--raises

is

    Create(amaterial : CString from Standard)
    
    ---Level: Internal 
    
    ---Purpose: Creates the material <amaterial>.
    
    returns mutable Material from Materials;
    
    Name(me) returns AsciiString from TCollection
    
    ---Level: Public 
    
    ---Purpose: Returns the name of the material.
    
    is static;
    
    Dump(me ; astream : in out OStream)
    
    ---Level: Internal 
    
    ---Purpose: Useful for debugging.
    
    is redefined;
    
fields

    thematerial      : HAsciiString from TCollection;

end Material;
