-- Created on: 1999-02-12
-- Created by: Andrey BETENEV
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class TranslateCurveBoundedSurface from StepToTopoDS 
    inherits Root from StepToTopoDS
    ---Purpose: Translate curve_bounded_surface into TopoDS_Face

uses
    TransientProcess from Transfer,
    CurveBoundedSurface from StepGeom,
    Face                from TopoDS

is
    Create returns TranslateCurveBoundedSurface;
        ---Purpose: Create empty tool

    Create (CBS: CurveBoundedSurface from StepGeom;
    	    TP: TransientProcess from Transfer)
    	returns TranslateCurveBoundedSurface;
        ---Purpose: Translate surface
	
    Init (me: in out;
          CBS: CurveBoundedSurface from StepGeom;
    	  TP: TransientProcess from Transfer)
    	returns Boolean;
        ---Purpose: Translate surface
	
    Value (me) returns Face from TopoDS;
        ---Purpose: Returns result of last translation or null wire if failed.
	---C++: return const &

fields

    myFace: Face from TopoDS;

end TranslateCurveBoundedSurface;
