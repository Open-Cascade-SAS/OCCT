-- Created on: 2010-11-15
-- Created by: Sergey SLYADNEV
-- Copyright (c) 2010-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class NMTool from StepToTopoDS

    ---Purpose: Provides data to process non-manifold topology when
    --          reading from STEP.

uses
    DataMapOfRI        from StepToTopoDS,
    DataMapOfRINames   from StepToTopoDS,
    RepresentationItem from StepRepr,
    Shape              from TopoDS,
    AsciiString        from TCollection,
    ListOfShape        from TopTools
is

    Create returns NMTool from StepToTopoDS;
 
    Create(MapOfRI      : DataMapOfRI from StepToTopoDS;
           MapOfRINames : DataMapOfRINames from StepToTopoDS)
    returns NMTool from StepToTopoDS;
    
    Init(me           : in out;
         MapOfRI      : DataMapOfRI from StepToTopoDS;
         MapOfRINames : DataMapOfRINames from StepToTopoDS);

    SetActive(me       : in out;
              isActive : Boolean);

    IsActive(me : in out)
    returns Boolean;

    CleanUp(me: in out);

    IsBound(me : in out;
    	    RI : RepresentationItem from StepRepr) 
    returns Boolean from Standard;

    IsBound(me     : in out;
    	    RIName : AsciiString from TCollection) 
    returns Boolean from Standard;
	
    Bind(me : in out;
         RI : RepresentationItem from StepRepr;
         S  : Shape from TopoDS);

    Bind(me     : in out;
         RIName : AsciiString from TCollection;
         S      : Shape from TopoDS);
	 
    Find(me : in out;
         RI : RepresentationItem from StepRepr) 
    returns Shape from TopoDS;
    ---C++: return const &

    Find(me     : in out;
         RIName : AsciiString from TCollection) 
    returns Shape from TopoDS;
    ---C++: return const &

    RegisterNMEdge(me   : in out;
                   Edge : Shape from TopoDS);

    IsSuspectedAsClosing(me             : in out;
                         BaseShell      : Shape from TopoDS;
                         SuspectedShell : Shape from TopoDS)
    returns Boolean;

    IsPureNMShell(me    : in out;
                  Shell : Shape from TopoDS)
    returns Boolean;

    SetIDEASCase(me        : in out;
                 IDEASCase : Boolean);

    IsIDEASCase(me : in out)
    returns Boolean;

    isEdgeRegisteredAsNM(me   : in out;
                         Edge : Shape from TopoDS)
    returns Boolean
    is private;

    isAdjacentShell(me     : in out;
                    ShellA : Shape from TopoDS;
                    ShellB : Shape from TopoDS)
    returns Boolean
    is private;
    
fields

    myRIMap      : DataMapOfRI from StepToTopoDS;
    
    myRINamesMap : DataMapOfRINames from StepToTopoDS;

    myNMEdges    : ListOfShape from TopTools;
  
    myIDEASCase  : Boolean;
    
    myActiveFlag : Boolean;

end NMTool;
