-- Created on: 1991-11-21
-- Created by: NW,JPB,CAL
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class PickDescriptor from Visual3d

	---Version:

	---Purpose: This class contains the pick information.
	--	    It contains a certain number of PickPaths.

	---Keywords: Pick Descriptor, Path, Structure, PickId

	---Warning:
	---References:

uses

	Structure		from Graphic3d,
	ContextPick		from Visual3d,
	PickPath		from Visual3d,
	HSequenceOfPickPath	from Visual3d

raises

	PickError		from Visual3d

is

	Create ( CTX : ContextPick from Visual3d )
		returns PickDescriptor from Visual3d;
	---Level: Public
	---Purpose: Creates a PickDescriptor <me>.

	---------------------------------------------------
	-- Category: Methods to modify the class definition
	---------------------------------------------------

	AddPickPath ( me	: in out;
		      APickPath	: PickPath from Visual3d )
		is static;
	---Level: Public
	---Purpose: Adds a PickPath to PickDescriptor <me>.
	---Category: Methods to modify the class definition

	Clear ( me : in out )
		is static;
	---Level: Public
	---Purpose: Erases all the information in <me>.
	---Category: Methods to modify the class definition

	----------------------------
	-- Category: Inquire methods
	----------------------------

	Depth ( me )
		returns Integer from Standard
		is static;
	---Level: Public
	---Purpose: Returns the pick depth, that is the
	--	    number of PickPaths available in the PickDescriptor.
	---Category: Inquire methods

	PickPath ( me )
		returns HSequenceOfPickPath from Visual3d
		is static;
	---Level: Internal
	---Purpose: Returns the group of PickPaths of <me>.
	---Category: Inquire methods

	TopStructure ( me )
		returns Structure from Graphic3d
	---Level: Public
	---Purpose: Returns the root structure.
	--	    If the pick order was of the type TOO_TOPFIRST
	--	    then it's the first structure.
	--	    If the pick order was of the type TOO_BOTTOMFIRST
	--	    Then it's the last structure.
	--	    The pick order is set by the method SetOrder
	--	    from ContextPick.
	--  Category: Inquire methods
	--  Warning: Raises PickError if Depth == 0 (no picked structure).
	raises PickError from Visual3d is static;

	TopPickId ( me )
		returns Integer from Standard
	---Level: Public
	---Purpose: Returns the root structure pickid.
	--	    If the pick order was of the type TOO_TOPFIRST
	--	    then it's the first pickid.
	--	    If the pick order was of the type TOO_BOTTOMFIRST
	--	    then it's the last pickid.
	--	    The pick order is set by the method SetOrder
	--	    from ContextPick.
	--  Category: Inquire methods
	--  Warning: Raises PickError if Depth == 0 (no picked structure).
	raises PickError from Visual3d is static;

	TopElementNumber ( me )
		returns Integer from Standard
	---Level: Public
	---Purpose: Returns the root structure element number.
	--	    If the pick order was of the type TOO_TOPFIRST
	--	    then it's the first element number.
	--	    If the pick order was of the type TOO_BOTTOMFIRST
	--	    then it's the last element number.
	--	    The pick order is set by the method SetOrder
	--	    from ContextPick.
	--  Category: Inquire methods
	--  Warning: Raises PickError if Depth == 0 (no picked structure).
	raises PickError from Visual3d is static;

--

fields

--
-- Class	:	Visual3d_PickDescriptor
--
-- Purpose	:	Declaration of variables specific to the class
--			describing a pick.
--
-- Reminders 	: 	A pick return is defined by:
--			- a sequence of (Elem_number, Pick_Id, Struct_Id)
--			- a depth

	-- pick sequence
	MyPickPathSequence	:	HSequenceOfPickPath from Visual3d;

	-- context associated to a pick
	MyContext		:	ContextPick from Visual3d;

end PickDescriptor;
