-- File:        GeometricCurveSet.cdl
-- Created:     Mon Dec  4 12:02:27 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWGeometricCurveSet from RWStepShape

	---Purpose : Read & Write Module for GeometricCurveSet

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     GeometricCurveSet from StepShape,
     EntityIterator from Interface

is

	Create returns RWGeometricCurveSet;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable GeometricCurveSet from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : GeometricCurveSet from StepShape);

	Share(me; ent : GeometricCurveSet from StepShape; iter : in out EntityIterator);

end RWGeometricCurveSet;
