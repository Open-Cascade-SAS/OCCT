-- Created on: 1999-06-24
-- Created by: Sergey ZARITCHNY
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class CopyLabel from TDF 

	---Purpose: 

uses
 
    Boolean             from Standard,
    Label               from TDF,
    Attribute           from TDF,
    DataSet             from TDF,
    RelocationTable     from TDF,
    AttributeMap        from TDF,
    LabelMap            from TDF,
    IDFilter            from TDF


is
 
    Create  returns  CopyLabel  from TDF; 
    ---Purpose: Empty  constructor  
    
    Create(aSource,  aTarget  :  Label  from  TDF) 
      returns  CopyLabel  from TDF;  
    ---Purpose: CopyTool  
    
    Load(me  :  in  out;  aSource,  aTarget  :  Label  from  TDF);  
    ---Purpose: Loads  src  and  tgt  labels 
     
    UseFilter(me  :  in  out;  aFilter : IDFilter from TDF); 
    ---Purpose:  Sets  filter

    ExternalReferences(myclass;  Lab  :  Label  from  TDF; 
    	    	    	    	 aExternals:in  out  AttributeMap  from  TDF; 
    	    	    	    	 aFilter   :  IDFilter  from  TDF) 
      returns  Boolean  from  Standard; 
    ---Purpose: Check  external  references and  if  exist  fills  the  aExternals  Map 
     
    ExternalReferences(myclass;  aRefLab, Lab  :  Label  from  TDF; 
    	    	    	   aExternals    :  in  out  AttributeMap  from  TDF; 
			   aFilter       :  IDFilter  from  TDF;
    	    	    	   aDataSet      :  in  out  DataSet  from  TDF) ;
    ---Purpose: Check  external  references and  if  exist  fills  the  aExternals  Map 
     
    Perform(me:in  out);  
    ---Purpose:  performs  algorithm  of  selfcontained  copy 
     
    IsDone(me) 
      returns  Boolean  from  Standard;  
    ---C++:  inline      
	 
    RelocationTable(me)     	 
      returns  RelocationTable  from  TDF;  
    ---Purpose: returns  relocation  table 
    ---C++: return const&
    
fields
 
    myRT        :  RelocationTable  from  TDF;
    mySL        :  Label            from  TDF; --  source  label
    myTL        :  Label            from  TDF; --  target  label 
    myFilter    :  IDFilter         from  TDF;
    myMapOfExt  :  AttributeMap     from  TDF; --  map  of  attribute  with  external  reference
    myIsDone    :  Boolean          from  Standard;

end CopyLabel;
