-- Created on: 1995-01-06
-- Created by: Christophe MARION
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class FaceIsoLiner from HLRTopoBRep

uses
    Integer from Standard,
    Real    from Standard,
    Pnt     from gp,
    Line    from Geom2d,
    Face    from TopoDS,
    Edge    from TopoDS,
    Vertex  from TopoDS,
    Data    from HLRTopoBRep

is
    Perform( myclass;
             FI     :        Integer from Standard;
             F      :        Face    from TopoDS;
    	     DS     : in out Data    from HLRTopoBRep;
	     nbIsos :        Integer from Standard);

    MakeVertex( myclass;
                E   :        Edge from TopoDS;
                P   :        Pnt  from gp;
                Par :        Real from Standard;
                Tol :        Real from Standard;
    	        DS  : in out Data from HLRTopoBRep)
    returns Vertex from TopoDS; 

    MakeIsoLine( myclass;
             F   :        Face   from TopoDS;
	     Iso :        Line   from Geom2d;	
             V1  : in out Vertex from TopoDS;
             V2  : in out Vertex from TopoDS;
             U1  :        Real   from Standard;
             U2  :        Real   from Standard;
             Tol :        Real   from Standard;
             DS  : in out Data   from HLRTopoBRep);

end FaceIsoLiner;
