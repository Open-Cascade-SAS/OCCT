-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DegeneratePcurve from StepGeom 

inherits Point from StepGeom 

uses

	Surface from StepGeom, 
	DefinitionalRepresentation from StepRepr,
	HAsciiString from TCollection
is

	Create returns DegeneratePcurve;
	---Purpose: Returns a DegeneratePcurve


	Init (me : mutable;
	      aName : HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      aName : HAsciiString from TCollection;
	      aBasisSurface : Surface from StepGeom;
	      aReferenceToCurve : DefinitionalRepresentation from StepRepr) is virtual;

	-- Specific Methods for Field Data Access --

	SetBasisSurface(me : mutable; aBasisSurface : Surface);
	BasisSurface (me) returns Surface;
	SetReferenceToCurve(me : mutable; aReferenceToCurve : DefinitionalRepresentation);
	ReferenceToCurve (me) returns DefinitionalRepresentation;

fields

	basisSurface : Surface from StepGeom;
	referenceToCurve : DefinitionalRepresentation from StepRepr;

end DegeneratePcurve;
