-- Created on: 1994-10-24
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DrawableP3D from TestTopOpeDraw inherits Marker3D from Draw

    ---Purpose: 

uses  

    Color           from Draw,
    Display         from Draw,
    Text3D          from Draw,
    MarkerShape     from Draw,
    CString         from Standard,
    Pnt             from gp,
    Pnt2d           from gp,
    Circ            from gp
    
is

    Create (P : Pnt from gp; PColor : Color from Draw;
    	    moveX : Real = 0.0; moveY : Real = 0.0)
    returns DrawableP3D from TestTopOpeDraw;

    Create (P : Pnt from gp; PColor : Color from Draw;
    	    Text : CString; TextColor : Color from Draw;
    	    moveX : Real = 0.0; moveY : Real = 0.0)
    returns DrawableP3D from TestTopOpeDraw;

    Create (P : Pnt from gp; T : MarkerShape from Draw; PColor : Color from Draw;
    	    Text : CString from Standard; TextColor : Color from Draw;
	    Size : Integer from Standard = 2;
    	    moveX : Real = 0.0; moveY : Real = 0.0)
    returns DrawableP3D from TestTopOpeDraw;

    Create (P : Pnt from gp; T : MarkerShape from Draw; 
    	    PColor : Color from Draw;
    	    Text : CString from Standard; TextColor : Color from Draw;
    	    Tol : Real from Standard;
    	    moveX : Real = 0.0; moveY : Real = 0.0)
    returns DrawableP3D from TestTopOpeDraw;

    ChangePnt(me : mutable; P : Pnt);
    
    DrawOn(me; dis : in out Display from Draw)
    is redefined;
    
fields

    myPnt    : Pnt from gp;
    myText   : CString from Standard;
    myTextColor : Color from Draw;
    myMoveX  : Real from Standard;
    myMoveY  : Real from Standard;

    myText3D : Text3D from Draw;

end DrawableP3D;
