-- Created on: 1995-02-23
-- Created by: Remi LEQUETTE
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Interpretor from Draw 

	---Purpose: Provides  an  encapsulation of the TCL interpretor
	--          to define Draw commands.

uses

        SStream         from Standard,
	PInterp         from Draw,
	CommandFunction from Draw,
	AsciiString     from TCollection,
	ExtendedString  from TCollection

is

    Create returns Interpretor from Draw;
    
    Init(me : in out);

    Add(me : in out; Command  : CString;
    	             Help     : CString;
		     Function : CommandFunction from Draw;
		     Group    : CString = "User Commands");
	---Purpose: Creates a  new command  with name <Command>,  help
	--          string <Help> in group <Group>.
	--          <Function> implement the function.

    Add(me : in out; Command  : CString;
    	             Help     : CString;
		     FileName : CString ; 
		     Function : CommandFunction from Draw;
    	    	     Group    : CString = "User Commands");
	---Purpose: Creates a  new command  with name  <Command>, help
	--          string   <Help>   in   group  <Group>.  <Function>
	--          implement the function. 
	--           <FileName> is the name of the file that contains
	--           the implementation of the command
        --

    Remove(me : in out; Command : CString)
    returns Boolean;
	---Purpose: Removes   <Command>, returns true  if success (the
	--          command existed).
	
    --
    --  The result
    --

    Result(me) returns CString;
    
    Reset(me : in out);
	---Purpose: Resets the result to empty string
	
    Append(me : in out; Result : CString) returns Interpretor from Draw; 
	---Purpose: Appends to the result
	---C++: return &
	---C++: alias operator<<
    	
    Append(me : in out; Result : AsciiString from TCollection) 
    returns Interpretor from Draw; 
	---Purpose: Appends to the result
	---C++: return &
	---C++: alias operator<<
    	
    Append(me : in out; Result : ExtendedString from TCollection) 
    returns Interpretor from Draw; 
	---Purpose: Appends to the result
	---C++: return &
	---C++: alias operator<<
    	
    Append(me : in out; Result : Integer) returns Interpretor from Draw; 
	---Purpose: Appends  to the result
	---C++: return &
	---C++: alias operator<<
    	
    Append(me : in out; Result : Real) returns Interpretor from Draw; 
	---Purpose: Appends  to the result
	---C++: return &
	---C++: alias operator<<
    	
    Append(me : in out; Result : SStream) returns Interpretor from Draw; 
	---Purpose: Appends  to the result
	---C++: return &
	---C++: alias operator<<
    	
    AppendElement(me : in out; Result : CString);
	---Purpose: Appends to the result the string as a list element



    --
    --      Interpetation
    --      
    
    Eval(me : in out; Script : CString) 
    returns Integer;
	---Purpose: Eval the script and returns OK = 0, ERROR = 1
	
    RecordAndEval(me : in out; Script : CString; Flags : Integer = 0) 
    returns Integer;
	---Purpose: Eval the script and returns OK = 0, ERROR = 1
	--          Store the script in the history record.
	
    EvalFile(me : in out; FileName : CString) 
    returns Integer;
	---Purpose: Eval the content on the file and returns status
	
    Complete(myclass; Script : CString) returns Boolean;
	---Purpose: Returns True if the script is complete, no pending
	--          closing braces. (})
    
    Destroy(me : in out);
	---C++: alias ~

    --
    --  Access to Tcl_Interp
    --  

    Create(anInterp : PInterp from Draw)
    returns Interpretor from Draw;
    
    Set(me : in out; anInterp : PInterp from Draw);
    
    Interp (me) returns PInterp from Draw;

    SetDoLog (me: in out; doLog: Boolean);
    ---Purpose: Enables or disables logging of all commands and their
    -- results
    ---Level: Advanced

    SetDoEcho (me: in out; doEcho: Boolean);
    ---Purpose: Enables or disables eachoing of all commands and their
    -- results to cout
    ---Level: Advanced

    GetDoLog (me) returns Boolean;
    ---Purpose: Returns true if logging of commands is enabled
    ---Level: Advanced

    GetDoEcho (me) returns Boolean;
    ---Purpose: Returns true if echoing of commands is enabled
    ---Level: Advanced

    Log (me: in out) returns SStream;
    ---Purpose: Returns log stream
    ---Level: Advanced
    ---C++: return &
	
 fields
 
    isAllocated : Boolean from Standard;
    myInterp    : PInterp from Draw;

    myDoLog: Boolean;
    myDoEcho: Boolean;
    myLog: SStream from Standard;

end Interpretor;
