-- Created on: 1995-08-25
-- Created by: Remi LEQUETTE
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class HSurface from GeomAdaptor inherits GHSurface from GeomAdaptor

    	---Purpose: An interface between the services provided by any
    	-- surface from the package Geom and those required
    	-- of the surface by algorithms which use it.

uses
    Surface from Geom,
    Surface from GeomAdaptor

raises
    ConstructionError from Standard

is

    Create returns mutable HSurface from GeomAdaptor;
    	---C++: inline
    
    Create( AS : Surface from GeomAdaptor) returns mutable HSurface from GeomAdaptor;
    	---C++: inline

    Create( S : Surface from Geom) returns mutable HSurface from GeomAdaptor;
    	---C++: inline
    
    Create( S : Surface from Geom; UFirst,ULast,VFirst,VLast : Real; 
    	    TolU  :  Real  =  0.0; 
            TolV  :  Real  =  0.0) 
    returns  mutable HSurface from GeomAdaptor
    raises ConstructionError from Standard;
    	---Purpose: ConstructionError is raised if UFirst>ULast or VFirst>VLast
    	---C++: inline

end HSurface;
