-- File:        OrientedClosedShell.cdl
-- Created:     Mon Dec  4 12:02:28 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWOrientedClosedShell from RWStepShape

	---Purpose : Read & Write Module for OrientedClosedShell

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     OrientedClosedShell from StepShape,
     EntityIterator from Interface

is

	Create returns RWOrientedClosedShell;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable OrientedClosedShell from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : OrientedClosedShell from StepShape);

	Share(me; ent : OrientedClosedShell from StepShape; iter : in out EntityIterator);

end RWOrientedClosedShell;
