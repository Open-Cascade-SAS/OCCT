-- Created on: 1993-01-11
-- Created by: CKY / Contract Toubro-Larsen ( Anand NATRAJAN )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PWBArtworkStackup from IGESAppli  inherits IGESEntity

        ---Purpose: defines PWBArtworkStackup, Type <406> Form <25>
        --          in package IGESAppli
        --          Used to communicate which exchange file levels are to
        --          be combined in order to create the artwork for a
        --          printed wire board (PWB). This property should be
        --          attached to the entity defining the printed wire
        --          assembly (PWA) or if no such entity exists, then the
        --          property should stand alone in the file.

uses

        HAsciiString from TCollection,
        HArray1OfInteger from TColStd

raises OutOfRange

is

        Create returns PWBArtworkStackup;

        -- Specific Methods pertaining to the class

        Init (me           : mutable;
              nbPropVal    : Integer;
              anArtIdent   : HAsciiString;
              allLevelNums : HArray1OfInteger);
        ---Purpose : This method is used to set the fields of the class
        --           PWBArtworkStackup
        --       - nbPropVal    : number of property values
        --       - anArtIdent   : Artwork Stackup Identification
        --       - allLevelNums : Level Numbers

        NbPropertyValues (me) returns Integer;
        ---Purpose : returns number of property values

        Identification (me) returns HAsciiString from TCollection;
        ---Purpose : returns Artwork Stackup Identification

        NbLevelNumbers (me) returns Integer;
        ---Purpose : returns total number of Level Numbers

        LevelNumber (me; Index : Integer) returns Integer
        raises OutOfRange;
        ---Purpose : returns Level Number
        -- raises exception if Index <= 0 or Index > NbLevelNumbers

fields

--
-- Class    : IGESAppli_PWBArtworkStackup
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class PWBArtworkStackup.
--
-- Reminder : A PWBArtworkStackup instance is defined by :
--            - number of property values
--            - Artwork Stackup Identification string
--            - Level Numbers

        theNbPropertyValues    : Integer;
        theArtworkStackupIdent : HAsciiString;
        theLevelNumbers        : HArray1OfInteger;

end PWBArtworkStackup;
