-- Created on: 1993-07-16
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Update:      Frederic MAUPAS


package PBRep 

	---Purpose: This  package    describes  a persistent  Boundary
	--          Representation  Data Structure inherited from  the
	--          abstract Topology  defined in the PTopoDS package.
	--          The  geometric data  are provided by the PGeom and
	--          PGeom2d packages.

uses
    gp,          -- Elementary geometry
    PTopLoc,     -- Local coordinate systems
    TopAbs,      -- Enumerations : Orientation, ShapeType
    PTopoDS,     -- Abstract topological data structure
    GeomAbs,     -- Enumerations : Shape
    PGeom,       -- 3D geometry : curves and surfaces
    PGeom2d,     -- 2D geometry : curves in parametric space
    PPoly,       -- Persistent Triangulations and Polygons
    PColStd      -- Persistent Standard Collection 
    
is

    deferred class CurveRepresentation;

    deferred class GCurve;

    class Curve3D;

    class CurveOnSurface;

    class CurveOnClosedSurface;

    class Polygon3D;

    class PolygonOnTriangulation;

    class PolygonOnClosedTriangulation;

    class PolygonOnSurface;

    class PolygonOnClosedSurface;

    class CurveOn2Surfaces;

    deferred class PointRepresentation;

    class PointOnCurve;

    deferred class PointsOnSurface;

    class PointOnCurveOnSurface;

    class PointOnSurface;

    class TFace;

    class TEdge;

    class TVertex;

    class TFace1;

    class TEdge1;

    class TVertex1;

end PBRep;
