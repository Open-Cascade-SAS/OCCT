-- Created on: 1994-02-22
-- Created by: Jean Louis FRENKEL
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class AnglePresentation from Prs3d inherits Root from Prs3d
    	---Purpose: A framework to define the display of angles.
uses
    Presentation from Prs3d,
    Pnt from gp,
    Drawer from Prs3d,
    ExtendedString from TCollection
    	
is  
    Draw( myclass; aPresentation: Presentation from Prs3d;
    	    	   aDrawer: Drawer from Prs3d;
		   aText: ExtendedString from TCollection;
                   AttachmentPoint1: Pnt from gp;
		   AttachmentPoint2: Pnt from gp;
                   AttachmentPoint3: Pnt from gp;
		   OffsetPoint: Pnt from gp);
	---Purpose: Defines the representation of the angle between the
    	-- line defined by the points AttachmentPoint1 and
    	-- AttachmentPoint2 and the line defined by the points
    	-- AttachmentPoint1 and AttachmentPoint3.
    	-- The text aText is displayed at the point OffsetPoint,
    	-- and the drawer aDrawer specifies the display
    	-- attributes which angles will have.
    	-- The presentation object aPresentation stores the
    	-- information defined in this framework.
        
end AnglePresentation from Prs3d;
