-- Created on: 1993-02-24
-- Created by: Laurent PAINNOT
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class ConstraintCouple from AppParCurves
	    ---Purpose: associates an index and a constraint for an object.
    	    -- This couple is used by AppDef_TheVariational when performing approximations.
uses Constraint from AppParCurves

is 

    Create returns ConstraintCouple;
    	---Purpose: returns an indefinite ConstraintCouple.

    Create(TheIndex: Integer; Cons: Constraint)
    	---Purpose: Create a couple the object <Index> will have the 
    	--          constraint <Cons>.

    returns ConstraintCouple;


    Index(me)
    	---Purpose: returns the index of the constraint object.

    returns Integer
    is static;
    

    Constraint(me) 
    	---Purpose: returns the constraint of the object.

    returns Constraint
    is static;
    

    SetIndex(me: in out; TheIndex: Integer)
    	---Purpose: Changes the index of the constraint object.
    
    is static;
    
    
    SetConstraint(me: in out; Cons: Constraint)
    	---Purpose: Changes the constraint of the object.
    
    is static;
    
    
fields

myIndex:      Integer;
myConstraint: Constraint from AppParCurves;

end ConstraintCouple;
