-- Created on: 1996-12-05
-- Created by: Philippe MANGIN
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Tensor from BlendFunc 

	---Purpose: used to store the "gradient of gradient"

uses
Array1OfReal from TColStd,
Vector from math,
Matrix from math

raises DimensionError from Standard, 
       RangeError from Standard 

is
    Create(NbRow, NbCol, NbMat : Integer) 
    returns Tensor;
 
    Init(me : in out; InitialValue: Real)
	   ---Purpose:Initialize all the elements of a Tensor to InitialValue.
    is static;
 
    Value(me; Row, Col, Mat: Integer)
    	---Purpose: accesses (in read or write mode) the value of index <Row>,
    	--          <Col> and <Mat> of a Tensor.
    	--          An exception is raised if <Row>, <Col> or <Mat> are not
    	--          in the correct range.
    	---C++: alias operator() 
    	---C++: return const & 
    	---C++: inline
    returns Real
    is static;
    
    ChangeValue(me : in out; Row, Col, Mat: Integer)
    	---Purpose: accesses (in read or write mode) the value of index <Row>,
    	--          <Col> and <Mat> of a Tensor.
    	--          An exception is raised if <Row>, <Col> or <Mat> are not
    	--          in the correct range.
    	---C++: alias operator() 
    	---C++: return & 
    	---C++: inline
    returns Real
    is static;

    Multiply(me; Right: Vector; Product:out Matrix)
    raises DimensionError
    is static;
    

fields
    Tab     : Array1OfReal;
    nbrow   : Integer;
    nbcol   : Integer;
    nbmat   : Integer;
    nbmtcl  : Integer;
end ;
