-- Created on: 1998-08-04
-- Created by: Christian CAILLET
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class RWAutoDesignDocumentReference from RWStepAP214

	---Purpose : Read & Write Module for AutoDesignDocumentReference

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     AutoDesignDocumentReference from StepAP214,
     EntityIterator from Interface

is

	Create returns RWAutoDesignDocumentReference;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable AutoDesignDocumentReference from StepAP214);

	WriteStep (me; SW : in out StepWriter; ent : AutoDesignDocumentReference from StepAP214);

	Share(me; ent : AutoDesignDocumentReference from StepAP214; iter : in out EntityIterator);

end RWAutoDesignDocumentReference;
