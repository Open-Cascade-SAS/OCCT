-- Created on: 1995-02-24
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

generic class SurfProps from Contap 
    (TheSurface     as any;
     TheSurfaceTool as any)

	---Purpose: Internal tool used  to compute the  normal and its
	--          derivatives. 

uses Pnt from gp,
     Vec from gp

is

    Normale(myclass; S: TheSurface; U,V: Real from Standard;
                     P: out Pnt from gp;
		     N: out Vec from gp);

	---Purpose: Computes  the point <P>, and  normal vector <N> on
	--          <S> at parameters U,V.



    DerivAndNorm(myclass; S: TheSurface; U,V: Real from Standard;
                          P      : out Pnt from gp;
			  d1u,d1v: out Vec from gp;
		          N      : out Vec from gp);

	---Purpose: Computes  the point <P>, and  normal vector <N> on
	--          <S> at parameters U,V.



    NormAndDn(myclass; S: TheSurface; U,V: Real from Standard;
                       P        : out Pnt from gp;
		       N,Dnu,Dnv: out Vec from gp);

	---Purpose: Computes the point <P>, normal vector <N>, and its
	--          derivatives <Dnu> and <Dnv> on <S> at parameters U,V.


end SurfProps;
