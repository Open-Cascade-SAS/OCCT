-- Created on: 1993-03-23
-- Created by: BBL,JLF
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class X11Dump from ImageUtility

uses
	X11Display 	from ImageUtility,
	X11Window  	from ImageUtility,
	X11XImage  	from ImageUtility,
	X11GC		from ImageUtility,
	Image 		from Image,
	AsciiString 	from TCollection

raises
	TypeMismatch 	from Standard

is
	Create( DisplayName : AsciiString from TCollection ;
	        aImage      : Image from Image )
		returns X11Dump from ImageUtility ;
	---Level: Internal
	---Purpose : Create a new X11 Display,Window,Colormap,GC,XImage suitable
	--		for aImage .

	Create( aX11Dump    : X11Dump from ImageUtility ;
		aImage      : Image from Image )
		returns X11Dump from ImageUtility ;
	---Level: Internal
	---Purpose : Create a new X11 XImage and share Display,Window,Colormap,
	--	     GC with a previous aX11Dump ;

	X11GC ( me ) 
		returns X11GC from ImageUtility
		is static;
	X11Window ( me ) 
		returns X11Window from ImageUtility
		is static;
	X11Display ( me ) 
		returns X11Display from ImageUtility
		is static;
	X11XImage ( me )
		returns X11XImage from ImageUtility
		is static;

	UpdateX11Colormap ( me )
		is static;
	UpdateX11XImage ( me : in out )
		is static;
	DisplayX11XImage ( me )
		is static;

fields
	myDisplay : X11Display from ImageUtility ;
	myWindow  : X11Window  from ImageUtility ;
	myXImage  : X11XImage  from ImageUtility ;
	myGC      : X11GC      from ImageUtility ;
	myImage   : Image from Image ;
end ;
