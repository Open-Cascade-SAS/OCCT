-- Created on: 1991-03-05
-- Created by: Herve Legrand, Mireille MERCIEN
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

generic class QuickSort from SortTools (Item as any;
                                        Array as Array1 from TCollection(Item);
                                        Comparator as any)

	---Purpose: This class provides the QuickSort algorithm.

is

    Sort(myclass; TheArray : in out Array; Comp : Comparator);
    ---Purpose: Sort an array using the QuickSort algorithm.
    ---Level: Public

end;

