-- Created on: 1994-11-18
-- Created by: Marie Jose MARTZ
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class GeomVector from GeomToIGES inherits GeomEntity from GeomToIGES

    ---Purpose: This class implements the transfer of the Vector from Geom
    --          to IGES . These can be :
    --          . Vector
    --              * Direction
    --              * VectorWithMagnitude
  
uses
 
    Vector               from Geom,
    VectorWithMagnitude  from Geom,
    Direction            from Geom,
    Direction            from IGESGeom,
    GeomEntity           from GeomToIGES
     
is 
    
    Create returns GeomVector from GeomToIGES;


    Create(GE : GeomEntity from GeomToIGES)  
    	 returns GeomVector from GeomToIGES;
    ---Purpose : Creates a tool GeomVector ready to run and sets its
    --         fields as GE's.

    TransferVector   (me    : in out;
                      start : Vector from Geom)
    	 returns mutable Direction from IGESGeom;
    ---Purpose :  Transfert  a  GeometryEntity which  answer True  to  the
    --            member : BRepToIGES::IsGeomVector(Geometry).  If this
    --            Entity could not be converted, this member returns a NullEntity.


    TransferVector   (me    : in out;
                      start : VectorWithMagnitude from Geom)
    	 returns mutable Direction from IGESGeom;


    TransferVector   (me    : in out;
                      start : Direction from Geom)
    	 returns mutable Direction from IGESGeom;


end GeomVector;


