-- File:	IGESDimen_ToolGeneralSymbol.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolGeneralSymbol  from IGESDimen

    ---Purpose : Tool to work on a GeneralSymbol. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses GeneralSymbol from IGESDimen,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolGeneralSymbol;
    ---Purpose : Returns a ToolGeneralSymbol, ready to work


    ReadOwnParams (me; ent : mutable GeneralSymbol;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : GeneralSymbol;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : GeneralSymbol;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a GeneralSymbol <ent>, from
    --           its specific (own) parameters

    DirChecker (me; ent : GeneralSymbol) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : GeneralSymbol;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : GeneralSymbol; entto : mutable GeneralSymbol;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : GeneralSymbol;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolGeneralSymbol;
