-- Created on: 1993-07-06
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class CurveOn2Surfaces from PBRep inherits CurveRepresentation from PBRep

	---Purpose: Defines a continuity between two surfaces.

uses
    Surface  from PGeom,
    Location from PTopLoc,
    Shape    from GeomAbs
    
raises
    NullObject from Standard
    
is

    Create(S1 , S2  : Surface  from PGeom;
	   L1 , L2  : Location from PTopLoc;
	   C        : Shape    from GeomAbs)
    returns mutable CurveOn2Surfaces from PBRep;

    Surface(me) returns any Surface from PGeom
    is static;

    Surface2(me) returns any Surface from PGeom
    is static;

    Location2(me) returns Location from PTopLoc
    is static;

    Continuity(me) returns Shape from GeomAbs
    is static;
    
    IsRegularity(me) returns Boolean
	---Purpose: Returns True.
    is redefined;
    
fields
    mySurface    : Surface  from PGeom;
    mySurface2   : Surface  from PGeom;
    myLocation2  : Location from PTopLoc;
    myContinuity : Shape    from GeomAbs;

end CurveOn2Surfaces;
