-- File:	MXCAFDoc_GraphNodeRetrievalDriver.cdl
-- Created:	Fri Sep 29 10:42:30 2000
-- Author:	Pavel TELKOV
--		<det@nordox.nnov.matra-dtv.fr>
---Copyright:	 Matra Datavision 2000


class GraphNodeRetrievalDriver from MXCAFDoc inherits ARDriver from MDF

uses

     RRelocationTable from MDF,
     Attribute        from PDF,
     Attribute        from TDF,
     MessageDriver    from CDM

is

--    Create returns mutable GraphNodeRetrievalDriver from MXCAFDoc;
    Create (theMsgDriver : MessageDriver from CDM)
    returns mutable GraphNodeRetrievalDriver from MXCAFDoc;
    
    VersionNumber(me) returns Integer from Standard;
	---Purpose: Returns the version number from which the driver
	--          is available: 0.

    SourceType(me) returns Type from Standard;

    NewEmpty (me)  returns mutable Attribute from TDF;

    Paste(me;
    	  Source     :         Attribute from PDF;
    	  Target     : mutable Attribute from TDF;
    	  RelocTable : RRelocationTable  from MDF);

end GraphNodeRetrievalDriver;
