-- File:	BRepExtrema_ExtFF.cdl
-- Created:	Wed Feb  9 13:01:29 1994
-- Author:	Laurent PAINNOT
--		<lpa@phylox>
---Copyright:	 Matra Datavision 1994


class ExtFF from BRepExtrema

uses
    Integer           from Standard,
    Real              from Standard,
    Boolean           from Standard,
    Face              from TopoDS,
    SequenceOfReal    from TColStd,
    SequenceOfPOnSurf from Extrema,
    ExtSS             from Extrema,
    Pnt               from gp,
    HSurface          from BRepAdaptor
     
raises 
    NotDone      from StdFail,
    OutOfRange   from Standard,
    TypeMismatch from Standard

is
    Create returns ExtFF from BRepExtrema;

    Create(F1 : Face   from TopoDS;
           F2 : Face   from TopoDS)
    	---Purpose: It calculates all the distances.
    returns ExtFF from BRepExtrema;

    Initialize(me: in out; F2 : Face from TopoDS)
    	---Purpose: 
    is static;
    
    Perform(me: in out; F1 : Face   from TopoDS;
     	    	    	F2 : Face   from TopoDS)
    	---Purpose: An exception is raised if the fields have not been
    	--          initialized.
    	--          Be careful: this method uses the Face F2 only for 
    	--          classify, not for the fields.
    raises TypeMismatch from Standard
    is static;
    
    IsDone(me) returns Boolean from Standard
    	---Purpose: True if the distances are found.
    is static;
    
    IsParallel (me) returns Boolean
    	---Purpose: Returns True if the surfaces are parallel.
    is static;


    NbExt(me) returns Integer from Standard
    	---Purpose: Returns the number of extremum distances.
    raises NotDone from StdFail
    is static;

    
    SquareDistance(me; N : Integer from Standard) returns Real from Standard
    	---Purpose: Returns the value of the <N>th extremum square distance.
    raises NotDone    from StdFail,
    	   OutOfRange from Standard
    is static;
    
    
    ParameterOnFace1(me; N : Integer from Standard; U, V: out Real)
    	---Purpose: Returns the parameters on the  Face F1 of the  <N>th
    	--          extremum distance.
    raises NotDone    from StdFail,
    	   OutOfRange from Standard
    is static;
    

    ParameterOnFace2(me; N : Integer from Standard; U, V: out Real) 
    	---Purpose: Returns the parameters on the  Face F2 of the  <N>th
    	--          extremum distance.
    raises NotDone    from StdFail,
    	   OutOfRange from Standard
    is static;
    
    
    PointOnFace1(me; N : Integer from Standard) returns Pnt from gp
    	---Purpose: Returns the Point of the <N>th extremum distance.
    raises NotDone    from StdFail, 
    	   OutOfRange from Standard
    is static;


    PointOnFace2(me; N : Integer from Standard) returns Pnt from gp
    	---Purpose: Returns the Point of the <N>th extremum distance.
    raises NotDone    from StdFail, 
    	   OutOfRange from Standard
    is static;
    
    
fields
    myExtrem    : ExtSS             from Extrema;
    mynbext     : Integer           from Standard;
    mySqDist    : SequenceOfReal    from TColStd;
    myPointsOnS1: SequenceOfPOnSurf from Extrema;
    myPointsOnS2: SequenceOfPOnSurf from Extrema;
    myHS        : HSurface          from BRepAdaptor;
end ExtFF;





