-- Created on: 2007-05-29
-- Created by: Vlad Romashko
-- Copyright (c) 2007-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class BooleanArrayRetrievalDriver from MDataStd inherits ARDriver from MDF

uses 

    RRelocationTable from MDF,
    Attribute        from TDF,
    Attribute        from PDF, 
    MessageDriver    from CDM

is

    Create(theMessageDriver : MessageDriver from CDM)
    returns mutable BooleanArrayRetrievalDriver from MDataStd;

    VersionNumber(me) returns Integer from Standard;

    SourceType(me) returns Type from Standard;

    NewEmpty (me) returns mutable Attribute from TDF;

    Paste(me;
    	  Source     :         Attribute from PDF;
    	  Target     : mutable Attribute from TDF;
    	  RelocTable : RRelocationTable from MDF);

end BooleanArrayRetrievalDriver;
