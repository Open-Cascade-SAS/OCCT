-- Created on: 1999-06-30
-- Created by: Sergey ZARITCHNY
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


private class Translator from TNaming

	---Purpose: 

uses
    Shape  from  TopoDS, 
    DataMapOfShapeShape from  TopTools, 
    IndexedDataMapOfTransientTransient  from TColStd

is
 
    Create  returns  Translator  from  TNaming; 
     
    Add(me  : in  out;  aShape  :  Shape  from  TopoDS); 
     
    Perform (me  :  in  out); 
     
    IsDone(me) 
    	returns  Boolean  from  Standard;
     
    Copied(me;  aShape  :  Shape  from  TopoDS)   
    returns  Shape   from  TopoDS;  
    ---Purpose: returns copied  shape
    ---C++  :  return  const 
     
    Copied(me)   
    returns  DataMapOfShapeShape   from  TopTools; 
     ---C++  :  return  const&
     ---Purpose: returns  DataMap  of  results;  (shape <-> copied  shape)
    DumpMap(me;  isWrite  :  Boolean  from  Standard  =  Standard_False); 
    
fields  

    myIsDone           : Boolean       from Standard;
    myMap              : IndexedDataMapOfTransientTransient  from TColStd;  
    myDataMapOfResults : DataMapOfShapeShape  from  TopTools;
--    myListOfShape    : ListOfShape   from  TopTools;
--    myListOfResult   : ListOfShape   from  TopTools;
    
end Translator;
