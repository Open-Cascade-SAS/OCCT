-- Created on: 2003-05-21
-- Created by: Open CASCADE Support
-- Copyright (c) 2003-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class LoaderParent from QANewBRepNaming

uses
    Shape from TopoDS,
    Builder from TNaming,
    DataMapOfShapeShape from TopTools,
    ShapeEnum from TopAbs

is

    LoadGeneratedDangleShapes (myclass; ShapeIn : Shape from TopoDS;
    	    	    	    	    	GeneratedFrom : ShapeEnum from TopAbs;
    	    	    	    	    	GenBuider : in out Builder from TNaming);

    GetDangleShapes (myclass; ShapeIn : Shape from TopoDS;
    	    	    	      GeneratedFrom : ShapeEnum from TopAbs;
    	    	    	      Dangles : in out DataMapOfShapeShape from TopTools)
    returns Boolean from Standard;

end LoaderParent from QANewBRepNaming;
