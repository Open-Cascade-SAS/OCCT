-- Created on: 1998-02-04
-- Created by: Julia GERASIMOVA
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class C0RegularityFilter from AIS inherits Filter from SelectMgr 

	---Purpose: 

uses
    EntityOwner       from SelectMgr,
    Shape             from TopoDS,
    ShapeEnum         from TopAbs,
    MapOfShape        from TopTools

is
    Create( aShape : Shape from TopoDS )
    returns C0RegularityFilter from AIS;
    
    ActsOn( me; aType : ShapeEnum from TopAbs )
    returns Boolean from Standard
    is redefined;
    
    IsOk( me; EO : EntityOwner from SelectMgr )
    returns Boolean from Standard is redefined virtual;

fields

    myMapOfEdges : MapOfShape from TopTools;

end C0RegularityFilter;
