-- Created on: 2000-01-28
-- Created by: data exchange team
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class BasicMsgRegistrator from ShapeExtend inherits TShared from MMgt

    ---Purpose: Abstract class that can be used for attaching messages
    --          to the objects (e.g. shapes).
    --          It is used by ShapeHealing algorithms to attach a message
    --          describing encountered case (e.g. removing small edge from
    --          a wire).
    --
    --          The methods of this class are empty and redefined, for instance,
    --          in the classes for Data Exchange processors for attaching
    --          messages to interface file entities or CAS.CADE shapes.

uses

    Shape   from TopoDS,
    Msg     from Message,
    Gravity from Message
     
is

    Create returns BasicMsgRegistrator from ShapeExtend;
    	---Purpose: Empty constructor.

    Send (me: mutable; object : Transient;
    	    	       message: Msg from Message;
    	    	       gravity: Gravity from Message) is virtual;
    	---Purpose: Sends a message to be attached to the object.
	--          Object can be of any type interpreted by redefined MsgRegistrator.

    Send (me: mutable; shape  : Shape from TopoDS;
    	    	       message: Msg from Message;
    	    	       gravity: Gravity from Message) is virtual;
    	---Purpose: Sends a message to be attached to the shape.

    Send (me: mutable; message: Msg from Message;
    	    	       gravity: Gravity from Message) is virtual;
    	---Purpose: Calls Send method with Null Transient.

end BasicMsgRegistrator;
