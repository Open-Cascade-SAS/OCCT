-- File:	TopOpeBRep_Hctxee2d.cdl
-- Created:	Thu Oct 29 12:39:50 1998
-- Author:	Jean Yves LEBEY
--		<jyl@langdox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1998

class Hctxee2d from TopOpeBRep inherits TShared from  MMgt

uses

    Shape from TopoDS,
    Edge from TopoDS,
    Surface from BRepAdaptor,
    Face from TopoDS,
    Curve from Geom2dAdaptor,
    CurveType from GeomAbs,
    Domain from IntRes2d
    
is

    Create returns mutable Hctxee2d from TopOpeBRep;
    SetEdges(me:mutable;E1,E2:Edge;BAS1,BAS2:Surface from BRepAdaptor);
    Edge(me;I:Integer) returns Shape;---C++ : return const &
    Curve(me;I:Integer) returns Curve from Geom2dAdaptor; ---C++ : return const &
    Domain(me;I:Integer) returns Domain from IntRes2d; ---C++ : return const &

fields

    myEdge1 : Edge from TopoDS;
    myCurve1 : Curve from Geom2dAdaptor;
    myCurveType1 : CurveType from GeomAbs;
    myDomain1 : Domain from IntRes2d;

    myEdge2 : Edge from TopoDS;
    myCurve2 : Curve from Geom2dAdaptor;
    myCurveType2 : CurveType from GeomAbs;
    myDomain2 : Domain from IntRes2d;

end Hctxee2d from TopOpeBRep;
