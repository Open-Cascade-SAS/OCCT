-- Created on: 1999-04-14
-- Created by: Roman LYGIN
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class SplitSurfaceContinuity from ShapeUpgrade inherits SplitSurface from ShapeUpgrade

    ---Purpose: Splits a Surface with a continuity criterion.
    --          At the present moment C1 criterion is used only.
    --          This tool works with tolerance. If C0 surface can be corrected
    --          at a knot with given tolerance then the surface is corrected,
    --          otherwise it is spltted at that knot.

uses

    Shape from GeomAbs

is

    Create returns mutable SplitSurfaceContinuity from ShapeUpgrade; 
        ---Purpose: Empty constructor.
	
    SetCriterion (me: mutable; Criterion: Shape from GeomAbs);
    	---Purpose: Sets criterion for splitting.
	
    SetTolerance (me: mutable; Tol: Real);
    	---Purpose: Sets tolerance.
	
    --Build (me: mutable; Segment: Boolean) is redefined;
    	--Purpose: Performs correction/splitting of the supporting surface(s).
	---         First defines splitting values, then calls inherited method.
    Compute(me: mutable; Segment: Boolean) is redefined;
    --Perform(me: mutable; Segment: Boolean);
fields

    myCriterion: Shape from GeomAbs;
    myTolerance: Real;
    myCont     : Integer;
    
end SplitSurfaceContinuity;
