-- Created on: 1993-03-18
-- Created by: Denis PASCAL
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

generic class ConnectedVerticesIterator  from GraphTools 
    	(Graph      as any;
     	 Vertex     as any;
         GIterator  as any;
	 CVIterator as any)	

--generic class ConnectedVerticesIterator from GraphTools
--            (Graph     as any;
--    	       Vertex    as any;
--	       GIterator as GraphIterator  (Graph,Vertex))
--	       CVIterator as ConnectedVerticesFromIterator

    ---Purpose: In a graph,  returns subsets of a  list of vertices in
    --          which all vertices are connected.
    
is

    Create    	
    	---Purpose: Create an empty algorithm.
    returns ConnectedVerticesIterator from GraphTools;
    
    Create (G : Graph)
	---Purpose: Create the   algorithm setting each vertex  of <G>
	--          reached by  GIterator tool, as initial conditions.
	--          Use Perform   method before visting  the result of
	--          the algorithm.
    returns ConnectedVerticesIterator from GraphTools;
    
    FromGraph (me : in out; G : Graph);	
    	---Purpose: Add each vertex of <G>  reached by GIterator  tool
	--          as   initial  conditions.   Use  Perform  method
	--          before   visiting the  result  of   the algorithm.
        ---Level: Public;
    
    FromVertex (me : in out; V : Vertex);
    	---Purpose: Add <V>  as   research condition.  This  method is
	--          cumulative.  User must used  Perform method before
	--          visting the result of the algorithm.
       ---Level: Public

    Reset (me : in out);
	---Purpose: Reset  the algorithm.  It may  be  reused with new
	--          initial conditions.  
	---Level: Public

    Perform (me : in out; G : Graph);       
    	---Purpose: Peform the  algorithm  in  <G> from initial  setted
       --          conditions.  
       ---Level: Public
    
    More(me)
	---Purpose: Returns   TRUE  if  there  are   others subset  of
	--          connected vertices.
        ---Level: Public
    returns Boolean from Standard;
    
    Next (me : in out);
	---Purpose: Set the iterator  to the next  subset of connected
	--          vertices.
        ---Level: Public
    
    NbVertices (me)
    returns Integer from Standard;
	---Purpose: Returns number of vertices  of the current  subset
	--          of connected vertices.
        ---Level: Public
    
    Value (me; index : Integer from Standard)
    returns any Vertex;
    ---Purpose: Returns a vertex  member of   the  current subset   of
    --          connected vertices.
    ---Level: Public
    ---C++: return const&         
    
fields

    myIterator : CVIterator;
    
end ConnectedVerticesIterator;







