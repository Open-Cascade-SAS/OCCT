-- Created on: 2002-12-12
-- Created by: data exchange team
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class CurveElementEndCoordinateSystem from StepFEA
inherits SelectType from StepData

    ---Purpose: Representation of STEP SELECT type CurveElementEndCoordinateSystem

uses
    FeaAxis2Placement3d from StepFEA,
    AlignedCurve3dElementCoordinateSystem from StepFEA,
    ParametricCurve3dElementCoordinateSystem from StepFEA

is
    Create returns CurveElementEndCoordinateSystem from StepFEA;
	---Purpose: Empty constructor

    CaseNum (me; ent: Transient) returns Integer;
	---Purpose: Recognizes a kind of CurveElementEndCoordinateSystem select type
	--          1 -> FeaAxis2Placement3d from StepFEA
	--          2 -> AlignedCurve3dElementCoordinateSystem from StepFEA
	--          3 -> ParametricCurve3dElementCoordinateSystem from StepFEA
	--          0 else

    FeaAxis2Placement3d (me) returns FeaAxis2Placement3d from StepFEA;
	---Purpose: Returns Value as FeaAxis2Placement3d (or Null if another type)

    AlignedCurve3dElementCoordinateSystem (me) returns AlignedCurve3dElementCoordinateSystem from StepFEA;
	---Purpose: Returns Value as AlignedCurve3dElementCoordinateSystem (or Null if another type)

    ParametricCurve3dElementCoordinateSystem (me) returns ParametricCurve3dElementCoordinateSystem from StepFEA;
	---Purpose: Returns Value as ParametricCurve3dElementCoordinateSystem (or Null if another type)

end CurveElementEndCoordinateSystem;
