-- Created on: 1995-08-25
-- Created by: Remi LEQUETTE
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class HCurve from Geom2dAdaptor inherits GHCurve from Geom2dAdaptor

	---Purpose: Provides an interface between the services provided by any
    	-- curve from the package Geom2d and those required
    	-- of the curve by algorithms, which use it.

uses
    Curve from Geom2d,
    Curve from Geom2dAdaptor

raises
    ConstructionError from Standard

is

    Create returns mutable HCurve from Geom2dAdaptor;
    
    Create( AS : Curve from Geom2dAdaptor) returns mutable HCurve from Geom2dAdaptor;

    Create( S : Curve from Geom2d) returns mutable HCurve from Geom2dAdaptor;
    
    Create( S : Curve from Geom2d; UFirst,ULast : Real) 
    returns  mutable HCurve from Geom2dAdaptor
    raises ConstructionError from Standard;
    	---Purpose: ConstructionError is raised if UFirst>ULast or VFirst>VLast

end HCurve;
