-- Created on: 1998-02-23
-- Created by: Christian CAILLET
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



deferred class Editor  from IFSelect    inherits TShared

    ---Purpose : An Editor defines a set of values and a way to edit them, on
    --           an entity or on the model (e.g. on its header)
    --           
    --           Each Value is controlled by a TypedValue, with a number (it is
    --           an Integer) and a name under two forms (complete and short)
    --           and an edit mode

uses CString, Messenger from Message,
     AsciiString from TCollection, HAsciiString from TCollection,
     Array1OfTransient from TColStd, Array1OfAsciiString from TColStd,
     Array1OfInteger from TColStd,   DictionaryOfInteger from Dico,
     HSequenceOfHAsciiString from TColStd,
     InterfaceModel from Interface,
     TypedValue from Interface, EditValue from IFSelect,
     EditForm from IFSelect, ListEditor from IFSelect

raises OutOfRange from Standard

is

    Initialize (nbval : Integer);
    ---Purpose : Prepares the list of Typed Values (gives its count)
    --           This count can be tuned later, to a LOWER value, this allows
    --           to initialize with a "maximum reservation" then cut the extra

    SetNbValues (me : mutable; nbval : Integer)
    ---Purpose : Adjusts the true count of values. It can be LOWER or equal to
    --           the initial size (which then acts as a reservation), but never
    --           greater
    	raises OutOfRange  is protected;
    --           Error if <nbval> exceeds the initial reservation

    SetValue (me : mutable; num : Integer;
    	      typval : TypedValue;
    	      shortname : CString = "";
    	      accessmode : EditValue = IFSelect_Editable);
    ---Purpose : Sets a Typed Value for a given ident and short name, with an
    --           Edit Mode

    SetList  (me : mutable; num : Integer; max : Integer = 0);
    ---Purpose : Sets a parameter to be a List
    --           max < 0 : not for a list (set when starting)
    --           max = 0 : list with no length limit (default for SetList)
    --           max > 0 : list limited to <max> items

    NbValues (me) returns Integer;
    ---Purpose : Returns the count of Typed Values

    TypedValue (me; num : Integer) returns TypedValue;
    ---Purpose : Returns a Typed Value from its ident

    IsList (me; num : Integer) returns Boolean;
    ---Purpose : Tells if a parameter is a list

    MaxList (me; num : Integer) returns Integer;
    ---Purpose : Returns max length allowed for a list
    --           = 0 means : list with no limit
    --           < 0 means : not a list

    Name  (me; num : Integer; isshort : Boolean = Standard_False) returns CString;
    ---Purpose : Returns the name of a Value (complete or short) from its ident
    --           Short Name can be empty

    EditMode (me; num : Integer) returns EditValue;
    ---Purpose : Returns the edit mode of a Value

    NameNumber   (me; name : CString) returns Integer;
    ---Purpose : Returns the number (ident) of a Value, from its name, short or
    --           complete. If not found, returns 0

    	-- Printings

    PrintNames (me; S : Messenger from Message);

    PrintDefs  (me; S : Messenger from Message; labels : Boolean = Standard_False);

    MaxNameLength (me; what : Integer) returns Integer;
    ---Purpose : Returns the MaxLength of, according to what :
    --           <what> = -1 : length of short names
    --           <what> =  0 : length of complete names
    --           <what> =  1 : length of values labels

    	-- Specific methods

    Label (me) returns AsciiString  is deferred;
    ---Purpose : Returns the specific label

    Form  (me; readonly : Boolean; undoable : Boolean = Standard_True)
    	returns EditForm  is virtual;
    ---Purpose : Builds and Returns an EditForm, empty (no data yet)
    --           Can be redefined to return a specific type of EditForm

    Recognize (me; form : EditForm) returns Boolean  is deferred;
    ---Purpose : Tells if this Editor can work on this EditForm and its content
    --           (model, entity ?)

    StringValue (me; form : EditForm;  num : Integer)
    	returns HAsciiString from TCollection  is deferred;
    ---Purpose : Returns the value of an EditForm, for a given item
    --           (if not a list. for a list, a Null String may be returned)

    ListEditor  (me; num : Integer) returns ListEditor  is virtual;
    ---Purpose : Returns a ListEditor for a parameter which is a List
    --           Default returns a basic ListEditor for a List, a Null Handle
    --           if <num> is not for a List. Can be redefined

    ListValue   (me; form : EditForm;  num : Integer)
    	returns HSequenceOfHAsciiString from TColStd  is virtual;
    ---Purpose : Returns the value of an EditForm as a List, for a given item
    --           If not a list, a Null Handle should be returned
    --           Default returns a Null Handle, because many Editors have
    --           no list to edit. To be redefined as required

    Load  (me; form : mutable EditForm; ent : Transient; model : InterfaceModel)
    	returns Boolean  is deferred;
    ---Purpose : Loads original values from some data, to an EditForm
    --           Remark: <ent> may be Null, this means all <model> is concerned
    --           Also <model> may be Null, if no context applies for <ent>
    --           And both <ent> and <model> may be Null, for a full static
    --           editor

    Update (me; form : mutable EditForm; num : Integer;
    	    newval : HAsciiString; enforce : Boolean)
    	returns Boolean  is virtual;
    ---Purpose : Updates the EditForm when a parameter is modified
    --           I.E.  default does nothing, can be redefined, as follows :
    --           Returns True when done (even if does nothing), False in case
    --           of refuse (for instance, if the new value is not suitable)
    --           <num> is the rank of the parameter for the EDITOR itself
    --           <enforce> True means that protected parameters can be touched
    --           
    --           If a parameter commands the value of other ones, when it is
    --           modified, it is necessary to touch them by Touch from EditForm

    UpdateList (me; form : mutable EditForm; num : Integer;
    	    newlist : HSequenceOfHAsciiString; enforce : Boolean)
    	returns Boolean  is virtual;
    ---Purpose : Acts as Update, but when the value is a list

    Apply (me; form : EditForm; ent : Transient; model : InterfaceModel)
    	returns Boolean  is deferred;
    ---Purpose : Applies modified values of the EditForm with some data
    --           Remark: <ent> may be Null, this means all <model> is concerned
    --           Also <model> may be Null, if no context applies for <ent>
    --           And both <ent> and <model> may be Null, for a full static
    --           editor

fields

    thenbval : Integer;
    themaxsh : Integer;
    themaxco : Integer;
    themaxla : Integer;
    thenames  : DictionaryOfInteger;
    thevalues : Array1OfTransient;
    theshorts : Array1OfAsciiString;
    themodes  : Array1OfInteger;
    thelists  : Array1OfInteger;

end Editor;
