-- File:        GeometricSet.cdl
-- Created:     Mon Dec  4 12:02:27 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWGeometricSet from RWStepShape

	---Purpose : Read & Write Module for GeometricSet

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     GeometricSet from StepShape,
     EntityIterator from Interface

is

	Create returns RWGeometricSet;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable GeometricSet from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : GeometricSet from StepShape);

	Share(me; ent : GeometricSet from StepShape; iter : in out EntityIterator);

end RWGeometricSet;
