-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Polyline from StepGeom 

inherits BoundedCurve from StepGeom 

uses

	HArray1OfCartesianPoint from StepGeom, 
	CartesianPoint from StepGeom, 
	HAsciiString from TCollection
is

	Create returns Polyline;
	---Purpose: Returns a Polyline


	Init (me : mutable;
	      aName : HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      aName : HAsciiString from TCollection;
	      aPoints : HArray1OfCartesianPoint from StepGeom) is virtual;

	-- Specific Methods for Field Data Access --

	SetPoints(me : mutable; aPoints : HArray1OfCartesianPoint);
	Points (me) returns HArray1OfCartesianPoint;
	PointsValue (me; num : Integer) returns CartesianPoint;
	NbPoints (me) returns Integer;

fields

	points : HArray1OfCartesianPoint from StepGeom;

end Polyline;
