-- Created on: 1992-08-18
-- Created by: Modelistation
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

private class Parameter from Hatch

	---Purpose: Stores an intersection on a line represented by :
	--          
	--          * A Real parameter.
	--          
	--          * A flag True when the parameter starts an interval.
	--          

uses
    Real    from Standard,
    Integer from Standard,
    Boolean from Standard

is
    Create;
    
    Create( Par1  : Real    from Standard;
            Start : Boolean from Standard;
	    Index : Integer from Standard = 0;
	    Par2  : Real    from Standard = 0)
    returns Parameter from Hatch;
    
fields
    myPar1  : Real      from Standard;
    myStart : Boolean   from Standard;
    myIndex : Integer   from Standard;
    myPar2  : Real      from Standard;
    
friends
    class Line    from Hatch,
    class Hatcher from Hatch

end Parameter;
