-- Created on: 2002-10-31
-- Created by: Michael SAZONOV
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DocumentRetrievalDriver from BinDrivers inherits DocumentRetrievalDriver from BinLDrivers

uses
    MessageDriver    from CDM,
    ADriverTable     from BinMDF, 
    Position         from Storage, 
    IStream          from Standard, 
    DocumentSection from BinLDrivers 
    
is
    -- ===== Public methods =====

    Create returns mutable DocumentRetrievalDriver from BinDrivers;
	---Purpose: Constructor

    AttributeDrivers  (me : mutable; theMsgDriver: MessageDriver from CDM)
	returns ADriverTable from BinMDF
	is redefined virtual;

    ReadShapeSection (me: mutable;
                      theSection : in out DocumentSection from BinLDrivers;
                      theIS      : in out IStream from Standard; 
    	    	      isMess     : Boolean from Standard = Standard_False) is redefined virtual;  
		       
    CheckShapeSection (me: mutable;
                      thePos : Position from Storage;
                      theIS  : in out IStream from Standard) is redefined virtual; 
		       
    PropagateDocumentVersion(me: mutable; theVersion : Integer from Standard) 
    	is redefined  virtual;		      
	
end DocumentRetrievalDriver;
