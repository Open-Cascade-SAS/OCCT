-- Created on: 2000-05-10
-- Created by: Andrey BETENEV
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1

class RepItemGroup from StepAP214
inherits Group from StepBasic

    ---Purpose: Representation of STEP entity RepItemGroup

uses
    HAsciiString from TCollection,
    RepresentationItem from StepRepr

is
    Create returns RepItemGroup from StepAP214;
	---Purpose: Empty constructor

    Init (me: mutable; aGroup_Name: HAsciiString from TCollection;
                       hasGroup_Description: Boolean;
                       aGroup_Description: HAsciiString from TCollection;
                       aRepresentationItem_Name: HAsciiString from TCollection);
	---Purpose: Initialize all fields (own and inherited)

    RepresentationItem (me) returns RepresentationItem from StepRepr;
	---Purpose: Returns data for supertype RepresentationItem
    SetRepresentationItem (me: mutable; RepresentationItem: RepresentationItem from StepRepr);
	---Purpose: Set data for supertype RepresentationItem

fields
    theRepresentationItem: RepresentationItem from StepRepr; -- supertype

end RepItemGroup;
