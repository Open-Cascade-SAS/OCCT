-- Created on: 1994-02-03
-- Created by: Gilles DEBARBOUILLE
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



generic class EnumerationParameter from Dynamic (Enum as any)

inherits

    Parameter from Dynamic     
    
    ---Purpose: This  generic class defines  a  parameter with a given
    --          enumeration.  For correct use an instanciation of this
    --          class,  the  Convert  method  must  be  defined.  This
    --          method is automaticaly called by the constructor which
    --          takes a  CString  as value for  the  enumeration.  The
    --          prototype  of the Convert method  must be described as
    --          follows :
    --          
    --          void Convert(const Standard_CString,Enum);
    --          
    --          The  prototype  and the body of  this   method, can be
    --          written  in   the  file   <mypackage.cxx>   where  the
    --          enumeration  is described.    No declaration  of   the
    --          Convert method in any .cdl file is necessary.


uses
    CString from Standard,
    OStream from Standard 

is

    Create(aparameter : CString from Standard)
    
    ---Level: Public 
    
    ---Purpose: Creates an  EnumerationParameter  of  <aparameter>  as
    --          name.

    returns mutable EnumerationParameter from Dynamic;

    Create(aparameter : CString from Standard; avalue : Enum)
    
    ---Level: Public 
    
    ---Purpose: Creates  an  EnumerationParameter  of  <aparameter> as
    --          name and <avalue> as value.

    returns mutable EnumerationParameter from Dynamic;
    
    Create(aparameter , avalue : CString from Standard) 

    ---Level: Public 
    
    ---Purpose: Creates an  EnumerationParameter  of  <aparameter>  as
    --          name  and <avalue> as value. The user has to define  a
    --          Convert method to translate  the string <avalue> in an
    --          enumeration term.

    returns mutable EnumerationParameter from Dynamic;
    
    Value(me) returns Enum
    
    ---Level: Public 
    
    ---Purpose: Returns the enumeration value <thevalue>.
    
    is static;
    
    Value (me : mutable ; avalue : Enum)
    
    ---Level: Public 
    
    ---Purpose: Sets the field <thevalue> with the enumeration value <avalue>

    is static;
    
    Dump(me ; astream : in out OStream from Standard)
    
    ---Level: Internal 
    
    ---Purpose: useful for debugging.
    
    is redefined;
    
fields

    thevalue : Enum;

end EnumerationParameter;
