-- Created on: 1991-04-24
-- Created by: Remi GILET
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

generic class Lin2d2Tan from GccIter (
    TheCurve          as any;
    TheCurveTool      as any;
    TheQualifiedCurve as any) -- as QualifiedCurve from GccEnt
    	    	      	      --                  (TheCurve)

	---Purpose: This class implements the algorithms used to 
	--          create 2d lines tangent to 2 other elements which
	--          can be circles, curves or points.
	--          More than one argument must be a curve.
	--
    	-- Note: Some constructors may check the type of the qualified argument 
    	--         and raise BadQualifier Error in case of incorrect couple (qualifier,
    	--         curv).
    	--         For example: "EnclosedCirc".

uses Pnt2d            from gp,
     Lin2d            from gp,
     QualifiedCirc    from GccEnt,
     Position         from GccEnt

raises BadQualifier from GccEnt,
       NotDone      from StdFail


private class FuncTCuCu instantiates FunctionTanCuCu from GccIter(
    	    	    	    	    	    TheCurve,TheCurveTool);

private class FuncTCuPt instantiates FunctionTanCuPnt from GccIter(
    	    	    	    	    	    TheCurve,TheCurveTool);

private class FuncTCirCu instantiates FunctionTanCirCu from GccIter(
    	    	    	    	    	    TheCurve,TheCurveTool);
is

Create (Qualified1 : TheQualifiedCurve ;
    	ThePoint   : Pnt2d             ;
        Param1     : Real              ;
    	Tolang     : Real              ) returns Lin2d2Tan from GccIter
    ---Purpose: This class implements the algorithms used to create 2d 
    --          lines passing thrue a point and tangent to a curve.
    --          Tolang is used to determine the tolerance for the 
    --          tangency points.
    --          Param2 is used for the initial guess on the curve.
raises BadQualifier from GccEnt;

Create (Qualified1 : QualifiedCirc     ;
        Qualified2 : TheQualifiedCurve ;
    	Param2     : Real              ;
    	Tolang     : Real              ) returns Lin2d2Tan from GccIter
raises BadQualifier from GccEnt;
    ---Purpose: This class implements the algorithms used to create 2d 
    --          line tangent to a circle and to a cuve.
    --          Tolang is used to determine the tolerance for the 
    --          tangency points.
    --          Param2 is used for the initial guess on the curve.
    --          Exception BadQualifier is raised in the case of 
    --          EnclosedCirc

Create (Qualified1 : TheQualifiedCurve ;
        Qualified2 : TheQualifiedCurve ;
    	Param1     : Real              ;
    	Param2     : Real              ;
    	Tolang     : Real              ) returns Lin2d2Tan from GccIter
raises BadQualifier from GccEnt;
    ---Purpose: This class implements the algorithms used to create 2d 
    --          line tangent to two curves.
    --          Tolang is used to determine the tolerance for the 
    --          tangency points.
    --          Param1 is used for the initial guess on the first curve.
    --          Param2 is used for the initial guess on the second curve.

--------------------------------------------------------------------------

IsDone (me) returns Boolean
is static;
    	---Purpose: This methode returns true when there is a solution 
    	--          and false in the other cases.

ThisSolution(me) returns Lin2d 
raises NotDone from StdFail
is static;
    ---Purpose: Returns the solution.

WhichQualifier(me                                 ; 
    	       Qualif1  : out Position from GccEnt;
    	       Qualif2  : out Position from GccEnt)
raises NotDone from StdFail
is static;
    -- It returns the informations about the qualifiers of the tangency 
    -- arguments concerning the solution number Index.
    -- It returns the real qualifiers (the qualifiers given to the 
    -- constructor method in case of enclosed, enclosing and outside 
    -- and the qualifiers computedin case of unqualified).

Tangency1(me                       ;
          ParSol,ParArg : out Real ;
          PntSol        : out Pnt2d)
raises NotDone from StdFail
is static;
    ---Purpose: Returns informations about the tangency point between the 
    --          result and the first argument.
    --          ParSol is the intrinsic parameter of the point PntSol on 
    --          the solution curv.
    --          ParArg is the intrinsic parameter of the point PntSol on 
    --          the argument curv.

Tangency2(me                       ;
          ParSol,ParArg : out Real ;
          PntSol        : out Pnt2d)
raises NotDone from StdFail
is static;
    -- Returns informations about the tangency point between the 
    -- result and the first argument.
    -- ParSol is the intrinsic parameter of the point PntSol on the solution
    -- curv.
    -- ParArg is the intrinsic parameter of the point PntSol on the argument
    -- curv.

fields

    WellDone : Boolean;
    -- True if the algorithm succeeded.

    linsol   : Lin2d;
    ---Purpose : The solutions.

    qualifier1 : Position from GccEnt;
    -- The qualifiers of the first argument.

    qualifier2 : Position from GccEnt;
    -- The qualifiers of the first argument.

    pnttg1sol   : Pnt2d;
    -- The tangency point between the solution and the first argument on 
    -- the solution.

    pnttg2sol   : Pnt2d;
    -- The tangency point between the solution and the second argument on 
    -- the solution.

    par1sol   : Real;
    -- The parameter of the tangency point between the solution and the 
    -- first argument on the solution.

    par2sol   : Real;
    -- The parameter of the tangency point between the solution and the 
    -- second argument on the solution.

    pararg1   : Real;
    -- The parameter of the tangency point between the solution and the first 
    -- argument on the first argument.

    pararg2   : Real;
    -- The parameter of the tangency point between the solution and the second 
    -- argument on the second argument.

end Lin2d2Tan;
