-- Created on: 1993-01-13
-- Created by: CKY / Contract Toubro-Larsen ( Deepak PRABHU )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class GeneralLabel from IGESDimen  inherits IGESEntity

        ---Purpose: defines GeneralLabel, Type <210> Form <0>
        --          in package IGESDimen
        --          Used for general labeling with leaders

uses

        GeneralNote          from IGESDimen,
        LeaderArrow          from IGESDimen,
        HArray1OfLeaderArrow from IGESDimen

raises OutOfRange

is

        Create returns mutable GeneralLabel;

        -- Specific Methods pertaining to the class

        Init (me          : mutable;
              aNote       : GeneralNote;
              someLeaders : HArray1OfLeaderArrow);
        ---Purpose : This method is used to set the fields of the class
        --           GeneralLabel
        --       - aNote       : General Note Entity
        --       - someLeaders : Associated Leader Entities

        Note (me) returns GeneralNote;
        ---Purpose : returns General Note Entity

        NbLeaders (me) returns Integer;
        ---Purpose : returns Number of Leaders

        Leader (me; Index : Integer) returns LeaderArrow
        raises OutOfRange;
        ---Purpose : returns Leader Entity
        -- raises exception if Index <= 0 or Index > NbLeaders()

fields

--
-- Class    : IGESDimen_GeneralLabel
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class GeneralLabel.
--
-- Reminder : A GeneralLabel instance is defined by :
--            - Note    : General Note Entity
--            - Leaders : Associated Leader Entities
-- An GeneralLabel Entity consists of a general note with one or more
-- associated leaders.

        theNote      : GeneralNote;
        theLeaders   : HArray1OfLeaderArrow;

end GeneralLabel;
