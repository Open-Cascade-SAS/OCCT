-- Created on: 1993-03-24
-- Created by: JCV
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Transformation from Geom2d inherits TShared from MMgt


        --- Purpose :
        --  The class Transformation allows to create Translation,
        --  Rotation, Symmetry, Scaling and complex transformations
        --  obtained by combination of the previous elementary
        --  transformations.        
        --  The Transformation class can also be used to
    	-- construct complex transformations by combining
    	-- these elementary transformations.
    	-- However, these transformations can never change
    	-- the type of an object. For example, the projection
    	-- transformation can change a circle into an ellipse,
    	-- and therefore change the real type of the object.
    	-- Such a transformation is forbidden in this
    	-- environment and cannot be a Geom2d_Transformation.
        --  The transformation can be represented as follow :
        --  
        --       V1   V2     T       
        --    | a11  a12    a14 |   | x |      | x'|
        --    | a21  a22    a24 |   | y |      | y'|
        --    |  0    0      1  |   | 1 |      | 1 |
        --
        --  where {V1, V2} defines the vectorial part of the
        --  transformation and T defines the translation part of 
        --  the transformation.
    	-- - Geom2d_Transformation transformations provide
    	--   the same kind of "geometric" services as
    	--   gp_Trsf2d ones but have more complex data
    	--   structures. The geometric objects provided by the
    	--   Geom2d package use gp_Trsf2d transformations
    	--   in the syntaxes Transform and Transformed.
    	-- - Geom2d_Transformation transformations are
    	--   used in a context where they can be shared by
    	--   several objects contained inside a common data structure.
        
uses Ax2d     from gp, 
     Pnt2d    from gp, 
     Trsf2d   from gp,
     TrsfForm from gp,
     Vec2d    from gp

raises ConstructionError from Standard,
       OutOfRange        from Standard

is


  Create   returns mutable Transformation;
        --- Purpose : Creates an identity transformation.


  Create (T : Trsf2d)  returns mutable Transformation;
        --- Purpose :  Creates a persistent copy of T.


  SetMirror (me : mutable; P : Pnt2d);
        --- Purpose :
        --  Makes the transformation into a symmetrical transformation
        --  with respect to a point P. 
        --  P is the center of the symmetry.


  SetMirror (me : mutable; A : Ax2d);
        --- Purpose :
        --  Makes the transformation into a symmetrical transformation
        --  with respect to an axis A. 
        --  A is the center of the axial symmetry.


  SetRotation (me : mutable; P : Pnt2d; Ang : Real);
        --- Purpose : Assigns to this transformation the geometric
    	-- properties of a rotation at angle Ang (in radians) about point P.
     
  SetScale (me : mutable; P : Pnt2d; S : Real);
        --- Purpose :
        --  Makes the transformation into a scale. P is the center of 
        --  the scale and S is the scaling value.


  SetTransformation (me : mutable; FromSystem1, ToSystem2 : Ax2d);
        --- Purpose :
        --  Makes a transformation allowing passage from the coordinate
        --  system "FromSystem1" to the coordinate system "ToSystem2".


  SetTransformation (me : mutable; ToSystem : Ax2d);
        --- Purpose :
        --  Makes the transformation allowing passage from the basic
        --  coordinate system
        --  {P(0.,0.,0.), VX (1.,0.,0.), VY (0.,1.,0.)}
        --  to the local coordinate system defined with the Ax2d ToSystem.


  SetTranslation (me : mutable; V : Vec2d);
        --- Purpose :
        --  Makes the transformation into a translation. 
        --  V is the vector of the translation.


  SetTranslation(me : mutable; P1, P2 : Pnt2d);            
        --- Purpose :
        --  Makes the transformation into a translation from the point
        --  P1 to the point P2.


  SetTrsf2d (me : mutable; T : Trsf2d);
        --- Purpose :
        --  Makes the transformation into a transformation T from 
        --  package gp.


  IsNegative (me)  returns Boolean;
        --- Purpose : Checks whether this transformation is an indirect
    	-- transformation: returns true if the determinant of the
    	-- matrix of the vectorial part of the transformation is less than 0.

  Form (me)  returns TrsfForm;
        --- Purpose :  Returns the nature of this transformation as a value
    	-- of the gp_TrsfForm enumeration.
    	--  Returns the nature of the transformation. It can be
	--  Identity, Rotation, Translation, PntMirror, Ax1Mirror,
	--  Scale, CompoundTrsf

                                                      
  ScaleFactor (me)  returns Real;
        --- Purpose :  Returns the scale value of the transformation. 


  Trsf2d (me)  returns Trsf2d;
        --- Purpose : Converts this transformation into a gp_Trsf2d transformation.
        --  Returns a non persistent copy of <me>.
    	-- -C++: return const&


  Value (me; Row, Col : Integer)   returns Real 
        --- Purpose :
        --  Returns the coefficients of the global matrix of tranformation.
        --  It is a 2 rows X 3 columns matrix.
     raises OutOfRange;
        --- Purpose :
        --  Raised if  Row < 1 or Row > 2  or  Col < 1 or Col > 2



        --- Purpose :
        --  Computes the reverse transformation. 

  Invert (me : mutable)
    	---Purpose: Computes the inverse of this transformation.
    	-- and  assigns the result to this transformatio
  raises ConstructionError;
        --- Purpose :
        --  Raised if the the transformation is singular. This means that 
        --  the ScaleFactor is lower or equal to Resolution from 
        --  package gp.


  Inverted (me)    returns mutable Transformation 
    	raises  ConstructionError;
    	---Purpose: Computes the inverse of this transformation and creates a new one.
        --  Raises ConstructionError  if the the transformation is singular. This means that 
        --  the ScaleFactor is lower or equal to Resolution from package gp.

    	
  Multiplied (me; Other : Transformation)  returns mutable Transformation;
        --- Purpose :
        --  Computes the transformation composed with Other and <me>.
        --  <me> * Other.
        --  Returns a new transformation
        ---C++: alias operator *


  Multiply (me : mutable; Other : Transformation);
        --- Purpose :
        --  Computes the transformation composed with Other and <me> .
        --  <me> = <me> * Other.
        ---C++: alias operator *=




        --- Purpose : 
        --  Computes the following composition of transformations
        --  if N > 0  <me> * <me> * .......* <me>.
        --  if N = 0  Identity
        --  if N < 0  <me>.Invert() * .........* <me>.Invert()

  Power (me : mutable; N : Integer)
     raises ConstructionError;
        --- Purpose :
        --  Raised if N < 0 and if the transformation is not inversible


  Powered (me; N : Integer) returns Transformation
     raises ConstructionError;
        --- Purpose :
        --  Raised if N < 0 and if the transformation is not inversible
 



  PreMultiply (me : mutable; Other : Transformation);
        --- Purpose :
        --  Computes the matrix of the transformation composed with 
        --  <me> and Other.     <me> = Other * <me>


  Transforms (me; X, Y : in out Real);
        --- Purpose :
        --  Applies the transformation <me> to the triplet {X, Y}.



  Copy (me)  returns mutable Transformation;
    	--- Purpose: Creates a new object, which is a copy of this transformation.
    
fields

  gpTrsf2d : Trsf2d;

end;
