-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class TextStyleWithBoxCharacteristics from StepVisual 

inherits TextStyle from StepVisual 

uses

	HArray1OfBoxCharacteristicSelect from StepVisual,
	BoxCharacteristicSelect from StepVisual,
	HAsciiString from TCollection, 
	TextStyleForDefinedFont from StepVisual
is

	Create returns mutable TextStyleWithBoxCharacteristics;
	---Purpose: Returns a TextStyleWithBoxCharacteristics


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aCharacterAppearance : mutable TextStyleForDefinedFont from StepVisual) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aCharacterAppearance : mutable TextStyleForDefinedFont from StepVisual;
	      aCharacteristics : HArray1OfBoxCharacteristicSelect) is virtual;

	-- Specific Methods for Field Data Access --

	SetCharacteristics(me : mutable; aCharacteristics :HArray1OfBoxCharacteristicSelect );
	Characteristics (me) returns HArray1OfBoxCharacteristicSelect;
	CharacteristicsValue (me; num : Integer) returns BoxCharacteristicSelect;
	NbCharacteristics (me) returns Integer;

fields

	characteristics : HArray1OfBoxCharacteristicSelect from StepVisual;

end TextStyleWithBoxCharacteristics;
