-- Created on: 1999-10-29
-- Created by: Pavel DURANDIN
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class UndefinedTypeHandler from GeomTools inherits TShared from MMgt

	---Purpose: 

uses

    Curve   from Geom,
    Surface from Geom,
    Curve   from Geom2d,
    OStream,
    IStream

is

    Create returns mutable UndefinedTypeHandler from GeomTools;
    
    -- Curve
    
    PrintCurve(me; C  : Curve from Geom;
    	      	   OS : in out OStream;
		   compact : Boolean = Standard_False) is virtual;
    
    ReadCurve(me; ctype: Integer;
    	    	  IS   : in out IStream;
    	    	  C    : in out Curve from Geom)
    returns IStream is virtual;
    ---C++: return &
    
    --PCurve
    
    PrintCurve2d(me; C  : Curve from Geom2d;
    	    	     OS : in out OStream;
		     compact : Boolean = Standard_False) is virtual;
    
    ReadCurve2d(me; ctype: Integer;
    	    	    IS   : in out IStream;
    	    	    C    : in out Curve from Geom2d)
    returns IStream is virtual;
    ---C++: return &
    
    --Surface
    
    PrintSurface(me; S  : Surface from Geom;
    	    	     OS : in out OStream;
		     compact : Boolean = Standard_False) is virtual;
    
    ReadSurface(me; ctype: Integer;
    	    	    IS   : in out IStream;
    	    	    S    : in out Surface from Geom)
    returns IStream is virtual;
    ---C++: return &
    
end UndefinedTypeHandler;
