-- Created on: 1999-04-14
-- Created by: Roman LYGIN
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class SplitCurve2dContinuity from ShapeUpgrade inherits SplitCurve2d from ShapeUpgrade

    	---Purpose: Corrects/splits a 2d curve with a continuity criterion.
    	--  Tolerance is used to correct the curve at a knot that respects
    	--  geometrically the criterion, in order to reduce the
    	--  multiplicity of the knot.

uses

    Curve from Geom2d,
    Shape from GeomAbs

is

    Create returns SplitCurve2dContinuity from ShapeUpgrade;
        ---Purpose: Empty constructor.
	
    SetCriterion (me: mutable; Criterion: Shape from GeomAbs);
    	---Purpose: Sets criterion for splitting.
	
    SetTolerance (me: mutable; Tol: Real);
    	---Purpose: Sets tolerance.
	
    
    Compute(me: mutable) is redefined;
    	---Purpose: Calculates points for correction/splitting of the curve
    


fields

    myCriterion: Shape from GeomAbs;
    myCont     : Integer;
    myTolerance: Real;
    
end SplitCurve2dContinuity;
