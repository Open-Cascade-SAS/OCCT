-- Created on: 1993-03-10
-- Created by: JCV
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Circle from Geom inherits Conic from Geom

        ---Purpose : Describes a circle in 3D space.
    	-- A circle is defined by its radius and, as with any conic
    	-- curve, is positioned in space with a right-handed
    	-- coordinate system (gp_Ax2 object) where:
    	-- - the origin is the center of the circle, and
    	-- - the origin, "X Direction" and "Y Direction" define the
    	--   plane of the circle.
    	-- This coordinate system is the local coordinate
    	-- system of the circle.
    	-- The "main Direction" of this coordinate system is the
    	-- vector normal to the plane of the circle. The axis, of
    	-- which the origin and unit vector are respectively the
    	-- origin and "main Direction" of the local coordinate
    	-- system, is termed the "Axis" or "main Axis" of the circle.
    	-- The "main Direction" of the local coordinate system
    	-- gives an explicit orientation to the circle (definition of
    	-- the trigonometric sense), determining the direction in
    	-- which the parameter increases along the circle.
    	-- The Geom_Circle circle is parameterized by an angle:
    	-- P(U) = O + R*Cos(U)*XDir + R*Sin(U)*YDir, where:
    	-- - P is the point of parameter U,
    	-- - O, XDir and YDir are respectively the origin, "X
    	-- Direction" and "Y Direction" of its local coordinate system,
    	-- - R is the radius of the circle.
    	-- The "X Axis" of the local coordinate system therefore
    	-- defines the origin of the parameter of the circle. The
    	-- parameter is the angle with this "X Direction".
    	-- A circle is a closed and periodic curve. The period is
    	-- 2.*Pi and the parameter range is [ 0, 2.*Pi [.


uses Ax2      from gp, 
     Circ     from gp,
     Pnt      from gp,
     Trsf     from gp, 
     Vec      from gp,
     Geometry from Geom


raises ConstructionError from Standard,
       RangeError        from Standard


is



  Create (C : Circ)   returns Circle;
    	---Purpose :  Constructs a circle by conversion of the gp_Circ circle C.


  Create (A2 : Ax2; Radius : Real)  returns Circle
        ---Purpose : Constructs a circle of radius Radius, where A2 locates the circle and
    	--   defines its orientation in 3D space such that:
    	--   - the center of the circle is the origin of A2,
    	--   - the origin, "X Direction" and "Y Direction" of A2
    	--    define the plane of the circle,
    	--   - A2 is the local coordinate system of the circle.
    	--  Note: It is possible to create a circle where Radius is equal to 0.0.
           raises ConstructionError;
	---Purpose : raised if Radius < 0.


  SetCirc (me : mutable; C : Circ)
        ---Purpose :
        --  Set <me> so that <me> has the same geometric properties as C.
  is static;


  SetRadius (me : mutable; R : Real)
    	---Purpose: Assigns the value R to the radius of this circle.
    	-- Note: it is possible to have a circle with a radius equal to 0.0.
    	-- Exceptions - Standard_ConstructionError if R is negative. 
     raises ConstructionError
  is static;


  Circ (me)   returns Circ
        ---Purpose :
        --  returns the non transient circle from gp with the same 
        --  geometric properties as <me>.
  is static;
  
  Radius(me) returns Real
  is static;
    	---Purpose: Returns the radius of this circle.
  
  ReversedParameter(me; U : Real) returns Real is redefined static;
    	---Purpose: Computes the parameter on the reversed circle for
    	-- the point of parameter U on this circle.
    	-- For a circle, the returned value is: 2.*Pi - U.


  Eccentricity (me)   returns Real is redefined static;
    	---Purpose : Returns the eccentricity  e = 0 for a circle.


  FirstParameter (me)   returns Real is redefined static;
        ---Purpose : Returns the value of the first parameter of this
    	-- circle. This is  0.0, which gives the start point of this circle, or
    	--  The start point and end point of a circle are coincident.


  LastParameter (me)   returns Real is redefined static;
        ---Purpose : Returns the value of the last parameter of this
    	-- circle. This is 2.*Pi, which gives the end point of this circle.
    	-- The start point and end point of a circle are coincident.


  IsClosed (me)   returns Boolean is redefined static;
        ---Purpose : returns True.


  IsPeriodic (me)  returns Boolean is redefined static;
        ---Purpose : returns True.


  D0(me; U : Real; P : out Pnt) is redefined static;
	---Purpose: Returns in P the point of parameter U.
        --  P = C + R * Cos (U) * XDir + R * Sin (U) * YDir
        --  where C is the center of the circle , XDir the XDirection and
        --  YDir the YDirection of the circle's local coordinate system.


  D1 (me; U : Real; P : out Pnt; V1 : out Vec) is redefined static;
        ---Purpose :
        --  Returns the point P of parameter U and the first derivative V1.


  D2 (me; U : Real; P : out Pnt; V1, V2 : out Vec) is redefined static;
        ---Purpose :
        --  Returns the point P of parameter U, the first and second 
        --  derivatives V1 and V2.


  D3 (me; U : Real; P : out Pnt; V1, V2, V3 : out Vec) is redefined static;
        ---Purpose :
        --  Returns the point P of parameter u, the first second and third
        --  derivatives V1 V2 and V3.
        

  DN (me; U : Real; N : Integer)   returns Vec
        ---Purpose :
        --  The returned vector gives the value of the derivative for the 
        --  order of derivation N.
    raises RangeError 
    is redefined static;
        ---Purpose : Raised if N < 1.   


  Transform (me : mutable; T : Trsf) is redefined static;
    	---Purpose: Applies the transformation T to this circle.

       
  Copy (me)  returns like me
  is redefined static;
    	---Purpose: Creates a new object which is a copy of this circle.

fields

  radius : Real;

end;

