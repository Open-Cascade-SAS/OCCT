-- File:        SizeSelect.cdl
-- Created:     Fri Dec  1 11:11:11 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993



class SizeSelect from StepBasic   inherits SelectType from StepData

	-- <SizeSelect> is an EXPRESS Select Type construct translation.
	-- it gathers : MeasureWithUnit (Entity), PositiveLengthMeasure (Real)

uses

    SelectMember from StepData

is

    Create returns SizeSelect;
    ---Purpose : Returns a SizeSelect SelectType

    CaseNum (me; ent : Transient) returns Integer;
    ---Purpose: Recognizes a TrimmingSelect Kind Entity that is :
    --        1 -> SizeMember
    --        0 else (i.e. Real)

    NewMember (me) returns SelectMember  is redefined;
    ---Purpose : Returns a SizeMember (POSITIVE_LENGTH_MEASURE) as preferred

    CaseMem (me; ent : SelectMember) returns Integer  is redefined;
    ---Purpose : Recognizes a SelectMember as Real, named as PARAMETER_VALUE
    --            1 -> PositiveLengthMeasure i.e. Real
    --            0 else (i.e. Entity)
	
    SetRealValue (me : in out; aReal : Real from Standard);
	
    RealValue (me) returns Real;
    ---Purpose : returns Value as a Real (Null if another type)
	
end SizeSelect;

