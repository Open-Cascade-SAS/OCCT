-- Created on: 1997-04-21
-- Created by: Prestataire Mary FABIEN
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Filter from TopOpeBRepDS 

---Purpose: 

uses

    Shape       from TopoDS,
    Edge        from TopoDS,
    ListOfShape from TopTools,
    IndexedMapOfShape from TopTools,
    
    Config                           from TopOpeBRepDS,    
    Interference                     from TopOpeBRepDS,
    ListOfInterference               from TopOpeBRepDS,
    ListIteratorOfListOfInterference from TopOpeBRepDS,
    ListOfShapeOn1State from TopOpeBRepDS,
    DataMapOfShapeListOfShapeOn1State from TopOpeBRepDS,
    HDataStructure from TopOpeBRepDS,
    PShapeClassifier from TopOpeBRepTool

is

    Create(HDS : HDataStructure from TopOpeBRepDS;
           pClassif: PShapeClassifier from TopOpeBRepTool = 0) returns Filter;

    ProcessInterferences(me : in out); -- oldies
    
    ProcessFaceInterferences(me : in out;
    	    	    	     MEsp : DataMapOfShapeListOfShapeOn1State from TopOpeBRepDS);
    ProcessFaceInterferences(me : in out; I : Integer;
	    		     MEsp : DataMapOfShapeListOfShapeOn1State from TopOpeBRepDS);

    ProcessEdgeInterferences(me : in out);
    ProcessEdgeInterferences(me : in out; I : Integer);

    ProcessCurveInterferences(me: in out);
    ProcessCurveInterferences(me: in out; I : Integer);


fields

    myHDS : HDataStructure from TopOpeBRepDS;
    myPShapeClassif: PShapeClassifier from TopOpeBRepTool;
    
end Filter from TopOpeBRepDS;
