-- Created on: 1999-09-24
-- Created by: Sergey ZARITCHNY
-- Copyright (c) 1999-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Box from QANewBRepNaming  inherits  TopNaming from QANewBRepNaming

    ---Purpose: To load the Box results 

uses MakeBox from BRepPrimAPI,
     Shape   from TopoDS,
     Label   from TDF,
     TypeOfPrimitive3D from QANewBRepNaming

is
 
    Create  returns  Box from QANewBRepNaming;
 
    Create  (ResultLabel :  Label from TDF) 
    returns  Box from QANewBRepNaming;

    Init(me : in out; ResultLabel : Label from TDF);


    Load (me; MakeShape : in out MakeBox from BRepPrimAPI; Type : TypeOfPrimitive3D from QANewBRepNaming);
      ---Purpose : Load  the box in  the data  framework  

    Back (me)   returns Label from TDF;
      ---Purpose : Returns the label of the back face of a box .
    
    Bottom (me) returns Label from TDF;
      ---Purpose : Returns the label of the  bottom face of a box .
    
    Front (me)  returns Label from TDF;
      ---Purpose : Returns the label of the  front face of a box .

    Left (me)   returns Label from TDF;
      ---Purpose : Returns the label of the  left face of a box .

    Right (me)  returns Label from TDF;
      ---Purpose : Returns the  label of the  right face of a box .

    Top (me)    returns Label from TDF;
      ---Purpose : Returns the  label of the  top face of a box . 
    
end Box;
