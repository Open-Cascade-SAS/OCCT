-- File:        PresentationSize.cdl
-- Created:     Mon Dec  4 12:02:29 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWPresentationSize from RWStepVisual

	---Purpose : Read & Write Module for PresentationSize

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     PresentationSize from StepVisual,
     EntityIterator from Interface

is

	Create returns RWPresentationSize;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable PresentationSize from StepVisual);

	WriteStep (me; SW : in out StepWriter; ent : PresentationSize from StepVisual);

	Share(me; ent : PresentationSize from StepVisual; iter : in out EntityIterator);

end RWPresentationSize;
