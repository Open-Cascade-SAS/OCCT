-- Created on: 1995-02-08
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



private class ParameterAndOrientation from GeomInt

	---Purpose: 

uses Orientation from TopAbs

is

    Create
    
    	returns ParameterAndOrientation from GeomInt;


    Create(P: Real from Standard; Or1,Or2: Orientation from TopAbs)
    
    	returns ParameterAndOrientation from GeomInt;


    SetOrientation1(me: in out; Or: Orientation from TopAbs)
    
    	is static;


    SetOrientation2(me: in out; Or: Orientation from TopAbs)
    
    	is static;


    Parameter(me)
    
    	returns Real from Standard
	is static;


    Orientation1(me)
    
    	returns Orientation from TopAbs
    	is static;


    Orientation2(me)
    
    	returns Orientation from TopAbs
    	is static;


fields

    prm : Real from Standard;
    or1 : Orientation from TopAbs;
    or2 : Orientation from TopAbs;

end ParameterAndOrientation;
