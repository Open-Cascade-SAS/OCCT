-- Created on: 1991-07-18
-- Created by: Arnaud BOUZY
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class GenExp from ExprIntrp inherits Generator from ExprIntrp

	---Purpose: This class permits, from a string, to create any 
	--          kind of expression of package Expr by using 
	--          built-in functions such as Sin,Cos, etc, and by 
	--          creating variables.

uses GeneralExpression from Expr,
    AsciiString from TCollection

raises NoSuchObject

is

    Create
    ---Purpose: Creates an empty generator
    ---Level: Advanced 
    returns GenExp is private;

    Create( myclass ) returns GenExp;
    
    Process(me : mutable; str : AsciiString)
    ---Purpose: Processes given string.
    ---Level: Advanced 
    is static;

    IsDone(me)
    ---Purpose: Returns false if any syntax error has occurred during 
    --          process. 
    ---Level: Advanced 
    returns Boolean
    is static;
	    
    Expression(me)
    ---Purpose: Returns expression generated. Raises an exception if 
    --          IsDone answers false.
    ---Level: Advanced 
    returns any GeneralExpression
    raises NoSuchObject
    is static;
    
fields

    done : Boolean;
    myExpression : GeneralExpression;
    
end GenExp;
