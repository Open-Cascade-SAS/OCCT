-- File:	RWStepShape_RWFaceBasedSurfaceModel.cdl
-- Created:	Fri Dec 28 16:02:01 2001 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class RWFaceBasedSurfaceModel from RWStepShape

    ---Purpose: Read & Write tool for FaceBasedSurfaceModel

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    FaceBasedSurfaceModel from StepShape

is
    Create returns RWFaceBasedSurfaceModel from RWStepShape;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : FaceBasedSurfaceModel from StepShape);
	---Purpose: Reads FaceBasedSurfaceModel

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: FaceBasedSurfaceModel from StepShape);
	---Purpose: Writes FaceBasedSurfaceModel

    Share (me; ent : FaceBasedSurfaceModel from StepShape;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWFaceBasedSurfaceModel;
