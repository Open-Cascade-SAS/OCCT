-- Created on: 1994-09-05
-- Created by: Gilles DEBARBOUILLE
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class CompositVariableInstance from Dynamic

inherits

    AbstractVariableInstance from Dynamic
	---Purpose: This  class corresponds to  the instanciation of a
	--          variable group. It allows the setting of more than
	--          one variable in  a variable instance. It is useful
	--          when a  method takes  a collection  of homogeneous
	--          objects as   argument. For   example a wire  needs
	--          edges as argument.
   
uses

    Variable     from Dynamic,
    VariableNode from Dynamic


is

    Create returns mutable CompositVariableInstance from Dynamic;
    
    ---Level: Advanced 
    
    ---Purpose: Creates  a new  empty  instance of   CompositVariable-
    --          Instance.
    
    Variable(me : mutable ; avariable : Variable from Dynamic)
    
    ---Purpose: Sets <avariable> into the collection of variable.
    
    is redefined;
    
    FirstVariableNode(me) returns VariableNode from Dynamic
    
    ---Purpose: Returns the first VariableNode  useful to explore  the
    --          list of variables addressed by <me>.
    
    is static;

fields

    thefirstvariablenode : VariableNode from Dynamic;

end CompositVariableInstance;
