-- Created on: 1998-04-17
-- Created by: Andre LIEUTIER
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class  HPG0G2Constraint  from  NLPlate  inherits  HPG0G1Constraint from  NLPlate 
---Purpose: define a PinPoint G0+G2  Constraint  used to load a Non Linear
--          Plate
uses
     XY from gp,
     XYZ from gp, 
     D1  from  Plate,
     D2  from  Plate
     
is
    Create(UV : XY; Value : XYZ; D1T : D1 from Plate; D2T : D2 from Plate) returns HPG0G2Constraint;
    -- create a G0+G2 Constraint
    -- 

    ActiveOrder(me)  returns  Integer 
    is   redefined; 
    --  returns the constraint active  order, i.e. the maximum between
    --  -- the initial constraint i.e 2 (for G2 Constraints)

 
    G2Target(me) returns D2 from Plate
    ---C++: return const &
    is  redefined; 
        

fields
     myG2Target : D2 from Plate; 
end;
