-- Created on: 1992-03-26
-- Created by: Herve LEGRAND
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package Geom2dLProp

    ---Purpose: Handles local properties of curves and surfaces from the 
    --          packages Geom and Geom2d.
    -- SeeAlso: Package LProp.


    ---Level : Public. 
    --  All methods of all  classes will be public.

uses Standard, gp, Geom2d, LProp

is
    
    class Curve2dTool;
    
    class CLProps2d from Geom2dLProp 
            instantiates CLProps from LProp(Curve         from Geom2d,
	                                    Vec2d         from gp,
					    Pnt2d         from gp,
					    Dir2d         from gp,
					    Curve2dTool   from Geom2dLProp); 
    class CurAndInf2d; 
    
    private class NumericCurInf2d instantiates NumericCurInf from LProp( 
    	    	    	    	    	       Curve         from Geom2d,
	                                       Vec2d         from gp,
					       Pnt2d         from gp,
					       Dir2d         from gp,
					       Curve2dTool   from Geom2dLProp); 
					    
end Geom2dLProp;    




