-- File:	RWStepDimTol_RWStraightnessTolerance.cdl
-- Created:	Wed Jun  4 13:34:34 2003 
-- Author:	Galina KULIKOVA
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWStraightnessTolerance from RWStepDimTol

    ---Purpose: Read & Write tool for StraightnessTolerance

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    StraightnessTolerance from StepDimTol

is
    Create returns RWStraightnessTolerance from RWStepDimTol;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : StraightnessTolerance from StepDimTol);
	---Purpose: Reads StraightnessTolerance

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: StraightnessTolerance from StepDimTol);
	---Purpose: Writes StraightnessTolerance

    Share (me; ent : StraightnessTolerance from StepDimTol;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWStraightnessTolerance;
