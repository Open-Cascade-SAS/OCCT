-- Created on: 1999-03-24
-- Created by: data exchange team
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class AssemblyExplorer from STEPSelections 

	---Purpose: 

uses
    
    Graph from Interface,
    SequenceOfAssemblyComponent        from STEPSelections,
    IndexedDataMapOfTransientTransient from TColStd,
    ProductDefinition                  from StepBasic,
    ShapeDefinitionRepresentation      from StepShape,
    AssemblyComponent                  from STEPSelections,
    NextAssemblyUsageOccurrence        from StepRepr
    
is
    
    Create (G: Graph) returns AssemblyExplorer from STEPSelections;
    
    Init(me: in out; G: Graph);
    
    Dump(me; os: in out OStream from Standard);
    
    FindSDRWithProduct(me; product: ProductDefinition from StepBasic)
    returns ShapeDefinitionRepresentation from StepShape;
    
    FillListWithGraph(me: in out; cmp: AssemblyComponent from STEPSelections);
    
    FindItemWithNAUO(me; nauo: NextAssemblyUsageOccurrence from StepRepr)
    returns Transient from Standard;
    
    --Methods for fetching the results
    
    NbAssemblies(me) returns Integer;
    	---Purpose: Returns the number of root assemblies;
	---C++: inline
    
    Root(me; rank: Integer = 1) returns AssemblyComponent from STEPSelections;
    	---Purpose: Returns root of assenbly by its rank;
	---C++: inline
    

fields

    myRoots: SequenceOfAssemblyComponent from STEPSelections;
    myGraph: Graph from Interface;
    myMap  : IndexedDataMapOfTransientTransient from TColStd;    

end AssemblyExplorer;
