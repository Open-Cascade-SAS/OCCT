-- Created on: 2003-03-05
-- Created by: Sergey KUUL
-- Copyright (c) 2003-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MaterialTool from XCAFDoc inherits Attribute from TDF

	---Purpose: Provides tools to store and retrieve attributes (materials)
	--          of TopoDS_Shape in and from TDocStd_Document
	--          A Document is intended to hold different 
	--          attributes of ONE shape and it's sub-shapes

uses
    Shape from TopoDS,
    Label from TDF,
    LabelSequence from TDF,
    Document from TDocStd,
    ShapeTool from XCAFDoc,
    RelocationTable from TDF,
    HAsciiString from TCollection

is
    Create returns MaterialTool from XCAFDoc;

    Set (myclass; L : Label from TDF) returns MaterialTool from XCAFDoc;
    	---Purpose: Creates (if not exist) MaterialTool.
    
    GetID (myclass)   
    ---C++: return const &  
    returns GUID from Standard;

    
    ---API: General structure
    
    BaseLabel(me) returns Label from TDF;
    	---Purpose: returns the label under which colors are stored
    
    ShapeTool (me: mutable) returns ShapeTool from XCAFDoc;
    	---Purpose: Returns internal XCAFDoc_ShapeTool tool
	---C++: return const &


    -- Methods for Material:

    IsMaterial (me; lab: Label from TDF) returns Boolean;
    	---Purpose: Returns True if label belongs to a material table and
        --          is a Material definition 
    
    GetMaterialLabels (me; Labels: out LabelSequence from TDF);
    	---Purpose: Returns a sequence of materials currently stored 
        --          in the material table
    
    AddMaterial (me; aName : HAsciiString from TCollection;
    	    	     aDescription : HAsciiString from TCollection;
    	    	     aDensity : Real from Standard;
    	    	     aDensName : HAsciiString from TCollection;
    	    	     aDensValType : HAsciiString from TCollection)
    returns Label from TDF;
    	---Purpose: Adds a Material definition to a table and returns its label

    SetMaterial (me; L: Label from TDF;
		     MatL: Label from TDF);
    	---Purpose: Sets a link with GUID
    
    SetMaterial (me; L: Label from TDF; aName : HAsciiString from TCollection;
    	    	     aDescription : HAsciiString from TCollection;
    	    	     aDensity : Real from Standard;
    	    	     aDensName : HAsciiString from TCollection;
    	    	     aDensValType : HAsciiString from TCollection);
    	---Purpose: Sets a link with GUID
    	--          Adds a Material as necessary
    
    GetMaterial (me; MatL: Label from TDF; aName : out HAsciiString from TCollection;
    	    	     aDescription : out HAsciiString from TCollection;
    	    	     aDensity : out Real from Standard;
    	    	     aDensName : out HAsciiString from TCollection;
    	    	     aDensValType : out HAsciiString from TCollection) returns Boolean;
        ---Purpose: Returns Material assigned to <MatL>
    	--          Returns False if no such Material is assigned
    
    GetDensityForShape (myclass; ShapeL: Label from TDF) returns Real from Standard;
        ---Purpose: Find referred material and return density from it
	--          if no material --> return 0


    ID (me)
    	---C++: return const & 
    returns GUID from Standard;

    Restore (me: mutable; with : Attribute from TDF);

    NewEmpty (me)
    returns mutable Attribute from TDF;

    Paste (me; into : mutable Attribute from TDF;
	       RT   : mutable RelocationTable from TDF);    

fields

    myShapeTool: ShapeTool from XCAFDoc;
    
end MaterialTool;

