-- Created on: 1993-11-08
-- Created by: Laurent BUCHARD
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

generic class WLine from ApproxInt ( 
    TheCurve        as any;
    TheCurveTool    as any;
    TheCurve2d      as any;
    TheCurveTool2d  as any)
    
    inherits TShared from MMgt
    
   
uses PntOn2S           from IntSurf,
     LineOn2S          from IntSurf
     
is 
     
     Create(CurveXYZ: TheCurve;
            CurveUV1: TheCurve2d;
	    CurveUV2: TheCurve2d)
	
	 returns mutable WLine from ApproxInt;

     Create(lin: LineOn2S from IntSurf;  Tang: Boolean from Standard)
     
	 returns mutable WLine from ApproxInt;
	 
     NbPnts(me) 
     
         returns Integer from Standard
	 is static;
	 
     Point(me: mutable; Index: Integer from Standard)
     
         returns PntOn2S from IntSurf
	 is static;
	 
fields 

    curvxyz  : TheCurve;
    curvuv1  : TheCurve2d;
    curvuv2  : TheCurve2d;
    pnton2s  : PntOn2S    from IntSurf;
    linon2s  : LineOn2S   from IntSurf;
end WLine;

