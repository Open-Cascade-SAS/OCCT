-- Created on: 1996-01-08
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



deferred class GeneratedShape from LocOpe inherits TShared from MMgt

	---Purpose:

uses Vertex      from TopoDS,
     Edge        from TopoDS,
     Face        from TopoDS,
     ListOfShape from TopTools

is


    GeneratingEdges(me: mutable)
    
    	returns ListOfShape from TopTools
	---C++: return const&
	is deferred;


    Generated(me: mutable; V: Vertex from TopoDS)
	---Purpose: Returns the  edge  created by  the  vertex <V>. If
	--          none, must return a null shape.
    	returns Edge from TopoDS
	is deferred;


    Generated(me: mutable; E: Edge from TopoDS)
	---Purpose: Returns the face created by the edge <E>. If none,
	--          must return a null shape.
    	returns Face from TopoDS
	is deferred;


    OrientedFaces(me: mutable)
	---Purpose: Returns  the  list of correctly oriented generated
	--          faces. 
    	returns ListOfShape from TopTools
	---C++: return const&
	is deferred;


fields

    myGEdges : ListOfShape from TopTools is protected;
    myList   : ListOfShape from TopTools is protected;

end GeneratedShape;
