-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class HalfSpaceSolid from StepShape 

inherits GeometricRepresentationItem from StepGeom

uses

	Surface from StepGeom,
	Boolean from Standard, 
	HAsciiString from TCollection
is

	Create returns mutable HalfSpaceSolid;
	---Purpose: Returns a HalfSpaceSolid


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aBaseSurface : mutable Surface from StepGeom;
	      aAgreementFlag : Boolean from Standard) is virtual;

	-- Specific Methods for Field Data Access --

	SetBaseSurface(me : mutable; aBaseSurface : mutable Surface);
	BaseSurface (me) returns mutable Surface;
	SetAgreementFlag(me : mutable; aAgreementFlag : Boolean);
	AgreementFlag (me) returns Boolean;

fields

	baseSurface : Surface from StepGeom;
	agreementFlag : Boolean from Standard;

end HalfSpaceSolid;
