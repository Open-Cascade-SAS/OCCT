-- File:        DimensionalExponents.cdl
-- Created:     Fri Dec  1 11:11:19 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class DimensionalExponents from StepBasic 

inherits TShared from MMgt

uses

	Real from Standard
is

	Create returns mutable DimensionalExponents;
	---Purpose: Returns a DimensionalExponents

	Init (me : mutable;
	      aLengthExponent : Real from Standard;
	      aMassExponent : Real from Standard;
	      aTimeExponent : Real from Standard;
	      aElectricCurrentExponent : Real from Standard;
	      aThermodynamicTemperatureExponent : Real from Standard;
	      aAmountOfSubstanceExponent : Real from Standard;
	      aLuminousIntensityExponent : Real from Standard) is virtual;

	-- Specific Methods for Field Data Access --

	SetLengthExponent(me : mutable; aLengthExponent : Real);
	LengthExponent (me) returns Real;
	SetMassExponent(me : mutable; aMassExponent : Real);
	MassExponent (me) returns Real;
	SetTimeExponent(me : mutable; aTimeExponent : Real);
	TimeExponent (me) returns Real;
	SetElectricCurrentExponent(me : mutable; aElectricCurrentExponent : Real);
	ElectricCurrentExponent (me) returns Real;
	SetThermodynamicTemperatureExponent(me : mutable; aThermodynamicTemperatureExponent : Real);
	ThermodynamicTemperatureExponent (me) returns Real;
	SetAmountOfSubstanceExponent(me : mutable; aAmountOfSubstanceExponent : Real);
	AmountOfSubstanceExponent (me) returns Real;
	SetLuminousIntensityExponent(me : mutable; aLuminousIntensityExponent : Real);
	LuminousIntensityExponent (me) returns Real;

fields

	lengthExponent : Real from Standard;
	massExponent : Real from Standard;
	timeExponent : Real from Standard;
	electricCurrentExponent : Real from Standard;
	thermodynamicTemperatureExponent : Real from Standard;
	amountOfSubstanceExponent : Real from Standard;
	luminousIntensityExponent : Real from Standard;

end DimensionalExponents;
