-- Created on: 1993-08-24
-- Created by: GG
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class FontMap from Xw inherits Transient 

	---Version: 0.0

	---Purpose: This class defines a FontMap object.

	---Keywords:
	---Warning:
	---References:

uses

	FontMap			from Aspect,
	FontMapEntry		from Aspect

raises

	FontMapDefinitionError	from Aspect,
	BadAccess from Aspect

is

	Create
	returns mutable FontMap from Xw
	is protected;
	---Level: Internal

	Create (Connexion : CString from Standard) 
	returns mutable FontMap from Xw 
	---Level: Public
	---Purpose: Creates a FontMap with an unallocated FontMapEntry.
	raises FontMapDefinitionError from Aspect;
	---Error if FontMap creation failed according
	--       to the supported hardware

	SetEntry (me : mutable; 
		  Entry : FontMapEntry from Aspect)
	---Level: Public
	---Purpose: Modifies an entry already defined or adds <Entry>
	--	    in the font map <me> if it don't exist.
	raises BadAccess from Aspect is virtual;
	---Purpose:  Warning if FontMap size is exceeded.
	--	   or FontMap is not defined properly
	--	   or FontMapEntry Index is out of range according
	--	   to the supported hardware

	SetEntries (me : mutable;
	          Fontmap : FontMap from Aspect)
	---Level: Public
	---Purpose: Modifies all entries of <me> from the new Fontmap.
	raises BadAccess from Aspect is virtual;
	---Purpose:  Warning if FontMap size is exceeded.
	--         or FontMap is not defined properly
	--         or One of new FontMapEntry Index is out of range according
	--         to the supported hardware

	Destroy (me : mutable) is virtual;
	---Level: Public
	---Purpose: Destroies the Fontmap
	---C++: alias ~

	----------------------------
	-- Category: Inquire methods
	----------------------------

	FreeFonts (me)
	returns Integer from Standard 
	---Level: Public
	---Purpose: Returns the number of Free Fonts in the Fontmap
	--	    depending of the HardWare
	raises BadAccess from Aspect is static;
	---Error If FontMap is not defined properly

	ExtendedFontMap (me)
	returns Address from Standard
	is static protected;
	---Level: Public
	---Purpose: Returns extended data fontmap structure pointer.
	---Category: Inquire methods


fields

	MyExtendedDisplay 	: Address from Standard;
	MyExtendedFontMap 	: Address from Standard;

friends

	class GraphicDevice from Xw

end FontMap;
