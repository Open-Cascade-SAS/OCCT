-- Created on: 1997-02-05
-- Created by: Alexander BRIVIN
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Instancing from Vrml 

	---Purpose: defines  "instancing" - using  the  same  instance  of  a  node   
	--          multiple  times.
	--  It  is  accomplished  by  using  the  "DEF"  and  "USE"  keywords.      
    	--  The  DEF  keyword  both  defines  a  named  node,  and  creates  a  single 
	--  instance  of  it.   
    	--  The  USE  keyword  indicates  that  the  most  recently  defined  instance 
    	--  should  be  used  again.   
    	--  If  several  nades  were  given  the  same  name,  then  the  last  DEF 
	--  encountered  during  parsing  "wins". 
	--  DEF/USE  is  limited  to  a  single  file.
uses

     AsciiString from TCollection

is
 
    Create ( aString        : AsciiString from TCollection ) 
        returns Instancing from Vrml;
 
        ---Purpose: Adds "DEF  <myName>" in  anOStream  (VRML  file).
    DEF ( me;  anOStream: in out OStream from Standard) returns OStream from Standard;
    ---C++:  return  & 

        ---Purpose: Adds "USE  <myName>" in  anOStream (VRML  file).
    USE ( me;  anOStream: in out OStream from Standard) returns OStream from Standard;
    ---C++:  return  & 

fields
 
    myName  : AsciiString from TCollection;  --  Name  using  DEF/USE  for a  node

end Instancing;

