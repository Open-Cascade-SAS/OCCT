-- File:	StepData_HeaderTool.cdl
-- Created:	Fri Jul 23 10:35:17 1993
-- Author:	Christian CAILLET
--		<cky@meteox>
---Copyright:	 Matra Datavision 1993


class HeaderTool  from StepData

    ---Purpose : HeaderTool exploits data from Header to build a Protocol :
    --           it uses the Header Entity FileSchema to do this.
    --           It builds a Protocol from the Global List of Protocols
    --           stored in the Library ReaderLib

uses OStream, AsciiString from TCollection, SequenceOfAsciiString from TColStd,
     StepReaderData, Protocol from StepData, FileProtocol

is

    Create (data : StepReaderData) returns HeaderTool;
    ---Purpose : Creates a HeaderTool from data read from a File. Computes the
    --           list of Schema Names. The Protocol will be computed later
    --           (because there are several options)

    Create (names : SequenceOfAsciiString from TColStd) returns HeaderTool;
    ---Purpose : Creates a HeaderTool directly from a list of Schema Names

    NbSchemaNames (me) returns Integer;
    ---Purpose : Returns the count of SchemaNames

    SchemaName (me; num : Integer) returns AsciiString from TCollection;
    ---Purpose : Returns a SchemaName, given its rank
    ---C++ : return const &

    NamedProtocol (me; name : AsciiString from TCollection)
    	returns Protocol from StepData;
    ---Purpose : Returns the Protocol which corresponds to a Schema Name
    --           Returns a Null Handle if this Schema Name is attached to no
    --           Protocol recorded in the Global List of ReaderLib

    	--  Building a Protocol  --

    Build (me : in out; protocol : mutable FileProtocol);
    ---Purpose : Fills a FileProtocol with the list of Protocols attached to
    --           the list of Schema Names. It can remain empty ...

    Protocol (me : in out) returns Protocol from StepData;
    ---Purpose : Returns a Protocol computed from the list of Schema Names :
    --           - a Null Handle if no SchemaName has been recognized (or list
    --             empty)
    --           - a single Protocol if only one SchemaName has been recognized
    --           - a FileProtocol with its componants if several SchemaNames
    --             have been recognized
    ---See also : method Ignored, to see if some SchemaNames were not
    --            recognized, then they remain Ignored

    IsDone (me) returns Boolean;
    ---Purpose : Returns True if either Build or Protocol has been called
    --           If it is False, Ignored and NbIgnored should not be called

    NbIgnoreds (me) returns Integer;
    ---Purpose : Returns the count of ignored SchemaNames (0 if all were OK)

    Ignored (me; num : Integer) returns AsciiString from TCollection;
    ---Purpose : Returns an ignored SchemaName, given its rank in the list of
    --           Ignored SchemaNames (not in the total list)
    ---C++ : return const &

    Print (me; S : in out OStream);
    ---Purpose : Sends the state of the HeaderTool in a comprehensive way,
    --           to an output stream

fields

    thenames   : SequenceOfAsciiString from TColStd;
    thedone    : Boolean;
    theignored : SequenceOfAsciiString from TColStd;

end HeaderTool;
