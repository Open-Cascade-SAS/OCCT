-- Created on: 1995-12-04
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.





class RWNamedUnit from RWStepBasic

	---Purpose : Read & Write Module for NamedUnit

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     NamedUnit from StepBasic,
     EntityIterator from Interface

is

	Create returns RWNamedUnit;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable NamedUnit from StepBasic);

	WriteStep (me; SW : in out StepWriter; ent : NamedUnit from StepBasic);

	Share(me; ent : NamedUnit from StepBasic; iter : in out EntityIterator);

end RWNamedUnit;
