-- Created on: 2008-04-10
-- Created by: Peter KURNEV <pkv@irinox>
-- Copyright (c) 2008-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class DiscretRoot from BRepMesh

inherits Transient from Standard

    ---Purpose:
    -- This is a common interface for meshing algorithms
    -- instantiated by Mesh Factory and implemented by plugins.

uses
    Shape from TopoDS

--raises

is
    Initialize
        returns DiscretRoot from BRepMesh;

    SetDeflection (           me : mutable;
                   theDeflection : Real from Standard);
    ---Purpose:
    -- Setup linear deflection.

    ---C++: alias "Standard_EXPORT virtual ~BRepMesh_DiscretRoot();"

    Deflection (me)
        returns Real from Standard;
    ---Purpose:
    -- Returns linear deflection.

    SetAngle (      me : mutable;
              theAngle : Real from Standard);
    ---Purpose:
    -- Setup angular deflection.

    Angle (me)
        returns Real from Standard;
    ---Purpose:
    -- Returns angular deflection.

    SetShape (      me : mutable;
              theShape : Shape from TopoDS);
    ---Purpose:
    -- Set the shape to triangulate.

    Shape (me)
        returns Shape from TopoDS;
    ---C++: return const &

    Perform (me : mutable)
        is deferred;
    ---Purpose:
    -- Compute triangulation for set shape.

    IsDone (me)
        returns Boolean from Standard;
    ---Purpose:
    -- Returns true if triangualtion was performed and has success.

    --
    --  Protected methods
    --
    SetDone (me : mutable)
        is protected;

    SetNotDone (me : mutable)
        is protected;

    Init (me : mutable)
        is virtual protected;

fields
    myDeflection : Real from Standard is protected;
    myAngle      : Real from Standard is protected;
    myShape      : Shape from TopoDS  is protected;
    myIsDone     : Boolean from Standard is protected;

end DiscretRoot;
