-- Created on: 1992-08-26
-- Created by: Remi GILET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class MakeElips from gce inherits Root from gce

    	---Purpose :This class implements the following algorithms used to 
    	--          create an ellipse from gp.
    	--          
    	--          * Create an ellipse from its center, and two points:
    	--            one on the ciconference giving the major radius, the 
    	--            other giving the value of the small radius.

uses Pnt   from gp,
     Ax2   from gp,
     Elips from gp

raises NotDone from StdFail

is

Create (A2 :                       Ax2  from gp;
        MajorRadius, MinorRadius : Real from Standard) 
    returns MakeElips;
    	--- Purpose :The major radius of the ellipse is on the "XAxis" and the
    	--           minor radius is on the "YAxis" of the ellipse. The "XAxis"
    	--           is defined with the "XDirection" of A2 and the "YAxis" is
    	--           defined with the "YDirection" of A2.
    	-- Warnings :
    	--           It is not forbidden to create an ellipse with 
    	--           MajorRadius = MinorRadius.

Create(S1,S2  : Pnt from gp;
       Center : Pnt from gp) returns MakeElips;
	---Purpose: Make an ellipse with its center and two points.
	-- Warning
    	-- The MakeElips class does not prevent the
    	-- construction of an ellipse where the MajorRadius is
    	-- equal to the MinorRadius.
    	-- If an error occurs (that is, when IsDone returns
    	-- false), the Status function returns:
    	-- -   gce_InvertRadius if MajorRadius is less than MinorRadius;
    	-- -   gce_NegativeRadius if MinorRadius is less than 0.0;
    	-- -   gce_NullAxis if the points S1 and Center are coincident; or
    	-- -   gce_InvertAxis if:
    	--   -   the major radius computed with Center and S1
    	--    is less than the minor radius computed with Center, S1 and S2, or
    	--   -   Center, S1 and S2 are collinear.         
		
Value(me) returns Elips from gp
    raises NotDone
    is static;
      	---C++: return const&
    	---Purpose: Returns the constructed ellipse.
    	-- Exceptions StdFail_NotDone if no ellipse is constructed.   
    
Operator(me) returns Elips from gp
    is static;
    	---C++: return const&
    	---C++: alias "Standard_EXPORT operator gp_Elips() const;"

fields

    TheElips : Elips from gp;
    --The solution from gp.
    
end MakeElips;




