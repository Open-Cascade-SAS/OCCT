-- Created on: 1995-12-07
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class GeometricRepresentationContextAndGlobalUnitAssignedContext from StepGeom 

inherits RepresentationContext from StepRepr


	--- This classe is an implementation of EXPRESS
	--  ANDOR Subtype Declaration.
uses

	GeometricRepresentationContext from StepGeom, 
	GlobalUnitAssignedContext from StepRepr, 
	HAsciiString from TCollection, 
	Integer from Standard, 
	HArray1OfNamedUnit from StepBasic,
	NamedUnit from StepBasic
is

	Create returns mutable GeometricRepresentationContextAndGlobalUnitAssignedContext;
	---Purpose: Returns a GeometricRepresentationContextAndGlobalUnitAssignedContext


	Init (me : mutable;
	      aContextIdentifier : mutable HAsciiString from TCollection;
	      aContextType : mutable HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      aContextIdentifier : mutable HAsciiString from TCollection;
	      aContextType : mutable HAsciiString from TCollection;
	      aGeometricRepresentationContext : mutable GeometricRepresentationContext from StepGeom;
	      aGlobalUnitAssignedContext : mutable GlobalUnitAssignedContext from StepRepr) is virtual;

	Init (me : mutable;
	      aContextIdentifier : mutable HAsciiString from TCollection;
	      aContextType : mutable HAsciiString from TCollection;
	      aCoordinateSpaceDimension : Integer from Standard;
	      aUnits : mutable HArray1OfNamedUnit from StepBasic) is virtual;

	-- Specific Methods for Field Data Access --

	SetGeometricRepresentationContext(me : mutable; aGeometricRepresentationContext : mutable GeometricRepresentationContext);
	GeometricRepresentationContext (me) returns mutable GeometricRepresentationContext;
	SetGlobalUnitAssignedContext(me : mutable; aGlobalUnitAssignedContext : mutable GlobalUnitAssignedContext);
	GlobalUnitAssignedContext (me) returns mutable GlobalUnitAssignedContext;

	-- Specific Methods for ANDOR Field Data Access --

	SetCoordinateSpaceDimension(me : mutable; aCoordinateSpaceDimension : Integer);
	CoordinateSpaceDimension (me) returns Integer;

	-- Specific Methods for ANDOR Field Data Access --

	SetUnits(me : mutable; aUnits : mutable HArray1OfNamedUnit);
	Units (me) returns mutable HArray1OfNamedUnit;
	UnitsValue (me; num : Integer) returns mutable NamedUnit;
	NbUnits (me) returns Integer;

fields

	geometricRepresentationContext : GeometricRepresentationContext from StepGeom;
	globalUnitAssignedContext : GlobalUnitAssignedContext from StepRepr;

end GeometricRepresentationContextAndGlobalUnitAssignedContext;
