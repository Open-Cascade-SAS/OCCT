-- Created on: 1993-12-06
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class BlendTool from BRepBlend

	---Purpose: 

uses 
     Pnt2d     from gp,
     State     from TopAbs,
     HCurve2d from Adaptor2d,
     HSurface from Adaptor3d,
     HVertex from Adaptor3d

is

    Project(myclass; P: Pnt2d from gp;
                     S: HSurface from Adaptor3d ;
                     C: HCurve2d from Adaptor2d ;
                     Paramproj: out Real from Standard;
                     Dist: out Real from Standard)

	---Purpose: Projects the point P on the arc C.
	--          If the methods returns Standard_True, the projection is
	--          successful, and Paramproj is the parameter on the arc
	--          of the projected point, Dist is the distance between
	--          P and the curve..
	--          If the method returns Standard_False, Param proj and Dist
	--          are not significant.
	--          

	returns Boolean from Standard;

    Inters (myclass; P1,P2: Pnt2d from gp;
                     S: HSurface from Adaptor3d ;
                     C: HCurve2d from Adaptor2d ;
                     Param: out Real from Standard;
                     Dist: out Real from Standard)
	returns Boolean from Standard;

    Parameter(myclass; V: HVertex from Adaptor3d; A: HCurve2d from Adaptor2d )
    
	---Purpose: Returns the parameter of the vertex V on the edge A.
    
	---C++: inline
    	returns Real from Standard;


    Tolerance(myclass; V: HVertex from Adaptor3d; A: HCurve2d from Adaptor2d )

	---Purpose: Returns the parametric tolerance on the arc A
	--          used to consider that the vertex and another point meet,
	--          i-e if Abs(Parameter(Vertex)-Parameter(OtherPnt))<=
	--          Tolerance, the points are "merged".

	---C++: inline
    	returns Real from Standard;


-- Methodes pour Rayon constant, en plus des 2 precedentes


    SingularOnUMin(myclass; S:HSurface from Adaptor3d )
    	returns Boolean from Standard;
    	---C++: inline

    SingularOnUMax(myclass; S:HSurface from Adaptor3d ) 
    	returns Boolean from Standard;
    	---C++: inline

    SingularOnVMin(myclass; S:HSurface from Adaptor3d )
    	returns Boolean from Standard;
    	---C++: inline

    SingularOnVMax(myclass; S:HSurface from Adaptor3d )
    	returns Boolean from Standard;
    	---C++: inline

    NbSamplesU(myclass; S: HSurface from Adaptor3d ;
                        u1,u2: Real from Standard)
        returns Integer from Standard;

    NbSamplesV(myclass; S: HSurface from Adaptor3d ;
                        v1,v2: Real from Standard)
        returns Integer from Standard;


    Bounds(myclass; C: HCurve2d from Adaptor2d ; 
                    Ufirst,Ulast: out Real from Standard);

	---Purpose: Returns the parametric limits on the arc C.
	--          These limits must be finite : they are either
	--          the real limits of the arc, for a finite arc,
	--          or a bounding box for an infinite arc.


    CurveOnSurf(myclass; C: HCurve2d from Adaptor2d ; S: HSurface from Adaptor3d )
	---C++: inline
    	returns HCurve2d from Adaptor2d ;


end BlendTool;
