-- Created on: 1998-07-22
-- Created by: data exchange team
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class ShapeTolerance from ShapeFix 

	---Purpose: Modifies tolerances of sub-shapes (vertices, edges, faces)

uses

    Shape     from TopoDS,
    ShapeEnum from TopAbs

is
    
    Create returns ShapeTolerance from ShapeFix;

    LimitTolerance (me; shape: Shape from TopoDS;
    	    	        tmin  : Real;
    	    	        tmax  : Real = 0.0;
    	    	        styp : ShapeEnum from TopAbs = TopAbs_SHAPE)
    returns Boolean;
    	---Purpose: Limits tolerances in a shape as follows :
    	--          tmin = tmax -> as SetTolerance (forces)
    	--          tmin = 0   -> maximum tolerance will be <tmax>
    	--          tmax = 0 or not given (more generally, tmax < tmin) ->
    	--             <tmax> ignored, minimum will be <tmin>
    	--          else, maximum will be <max> and minimum will be <min>
    	--          styp = VERTEX : only vertices are set
    	--          styp = EDGE   : only edges are set
    	--          styp = FACE   : only faces are set
    	--          styp = WIRE   : to have edges and their vertices set
    	--          styp = other value : all (vertices,edges,faces) are set
    	--          Returns True if at least one tolerance of the sub-shape has
    	--          been modified

    SetTolerance (me; shape: Shape from TopoDS;
    	    	      preci: Real;
    	    	      styp : ShapeEnum from TopAbs = TopAbs_SHAPE);
    	---Purpose: Sets (enforces) tolerances in a shape to the given value
    	--          styp = VERTEX : only vertices are set
    	--          styp = EDGE   : only edges are set
    	--          styp = FACE   : only faces are set
    	--          styp = WIRE   : to have edges and their vertices set
    	--          styp = other value : all (vertices,edges,faces) are set

end ShapeTolerance;
