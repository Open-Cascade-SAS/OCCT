-- Created on: 1992-05-22
-- Created by: Jean Claude VAUTHIER
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class BSplineCurve2d


from DrawTrSurf


inherits Curve2d from DrawTrSurf


uses BSplineCurve from Geom2d,
     Color from Draw,
     MarkerShape from Draw,
     Display from Draw,
     Drawable3D from Draw


is


  Create (C : BSplineCurve from Geom2d)
        --- Purpose :
        --  creates a drawable BSpline curve from a BSpline curve of 
        --  package Geom2d.
     returns BSplineCurve2d from DrawTrSurf;


  Create (C : BSplineCurve from Geom2d;
          CurvColor, PolesColor, KnotsColor : Color from Draw;
          KnotsShape : MarkerShape from Draw; KnotsSize : Integer;
          ShowPoles, ShowKnots : Boolean; Discret : Integer)
     returns BSplineCurve2d from DrawTrSurf;


  DrawOn (me; dis : in out Display from Draw)
     is redefined static;

  ShowPoles (me : mutable)
     is static;

  ShowKnots (me : mutable)
     is static;
     
  ClearPoles (me : mutable)
     is static;
  
  ClearKnots (me : mutable)
     is static;

  FindPole(me; X,Y : Real; D : Display from Draw; Prec : Real; 
           Index : in out Integer)
    ---Purpose: Returns in <Index> the index of the first pole  of the
    --          curve projected by the Display <D> at a distance lower
    --          than <Prec> from <X,Y>. If no pole  is found  index is
    --          set to 0, else index is always  greater than the input
    --          value of index.
  is static;

  FindKnot(me; X,Y : Real; D : Display from Draw; Prec : Real; 
           Index : in out Integer)
  is static;

  SetPolesColor (me : mutable; aColor : Color from Draw)
        ---C++: inline
     is static;

  SetKnotsColor (me : mutable; aColor : Color from Draw)
        ---C++: inline
     is static;

  SetKnotsShape (me : mutable; Shape : MarkerShape from Draw)
        ---C++: inline
     is static;

  KnotsShape (me)  returns MarkerShape from Draw
        ---C++: inline
     is static;
  
  KnotsColor (me)  returns Color from Draw
        ---C++: inline
     is static;
  
  PolesColor (me)  returns Color from Draw
        ---C++: inline
     is static;
    
  Copy(me) returns Drawable3D from Draw
	---Purpose: For variable copy.
  is redefined;
  
      
fields

  drawPoles  : Boolean;
  drawKnots  : Boolean;
  knotsForm  : MarkerShape from Draw;
  knotsLook  : Color from Draw;
  knotsDim   : Integer;
  polesLook  : Color from Draw;

end BSplineCurve2d;
