-- File:	StepFEA_FreedomsList.cdl
-- Created:	Sat Dec 14 11:02:05 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class FreedomsList from StepFEA
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity FreedomsList

uses
    HArray1OfDegreeOfFreedom from StepFEA

is
    Create returns FreedomsList from StepFEA;
	---Purpose: Empty constructor

    Init (me: mutable; aFreedoms: HArray1OfDegreeOfFreedom from StepFEA);
	---Purpose: Initialize all fields (own and inherited)

    Freedoms (me) returns HArray1OfDegreeOfFreedom from StepFEA;
	---Purpose: Returns field Freedoms
    SetFreedoms (me: mutable; Freedoms: HArray1OfDegreeOfFreedom from StepFEA);
	---Purpose: Set field Freedoms

fields
    theFreedoms: HArray1OfDegreeOfFreedom from StepFEA;

end FreedomsList;
