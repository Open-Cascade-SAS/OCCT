-- Created on: 1997-03-19
-- Created by: Prestataire Mary FABIEN
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Mesure from TestTopOpeTools

uses

    AsciiString from TCollection,
    Array1OfPnt from TColgp,
    HArray1OfPnt from TColgp,
    Pnt from gp

is

    Create returns Mesure from TestTopOpeTools;

    Create(name : AsciiString from TCollection)
    returns Mesure from TestTopOpeTools;

    Create(Pnts : HArray1OfPnt from TColgp)
    returns Mesure from TestTopOpeTools;

    Add(me :in out; n : in Integer from Standard; t : in Real from Standard);

    SetName(me : in out; Name : AsciiString from TCollection);

    Name(me) returns AsciiString from TCollection;
    ---C++: return const&

    Pnts(me) returns Array1OfPnt from TColgp;
    ---C++: return const&

    Pnt(me; I : in Integer) returns Pnt from gp;
    ---C++: return const&

    NPnts(me) returns Integer from Standard;

    Clear(me : in out);

fields

    myName  : AsciiString from TCollection;
    myPnts  : HArray1OfPnt from TColgp;
    myNPnts : Integer from Standard;

end Mesure from TestTopOpeTools;
