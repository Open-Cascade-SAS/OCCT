-- Created on: 1991-03-22
-- Created by: Philippe DAUTRY
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



package GccInt

	---Purpose: This package implements the services needed by the 
	--          toolkit Gcc to use curves other than lines or circles.
	--          This package is also used for intersections and 
	--          bisecting curves.

uses gp,
     MMgt,
     Standard

is

enumeration IType is Lin, Cir, Ell, Par, Hpr, Pnt;

deferred class Bisec;

class BCirc;

class BElips;

class BLine;

class BParab;

class BPoint;

class BHyper;

end GccInt;
