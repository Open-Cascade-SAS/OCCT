-- Created on: 1994-04-21
-- Created by: Christian CAILLET
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class SelectSignature  from IFSelect    inherits SelectExtract

    ---Purpose : A SelectSignature sorts the Entities on a Signature Matching.
    --           The signature to match is given at creation time. Also, the
    --           required match is given at creation time : exact (IsEqual) or
    --           contains (the Type's Name must contain the criterium Text)
    --           
    --           Remark that no more interpretation is done, it is an
    --           alpha-numeric signature : for instance, DynamicType is matched
    --           as such, super-types are not considered
    --           
    --           Also, numeric (integer) comparisons are supported : an item
    --           can be <val ou <=val or >val or >=val , val being an Integer
    --           
    --           A SelectSignature may also be created from a SignCounter,
    --           which then just gives its LastValue as SignatureValue

uses CString, AsciiString from TCollection, Transient,
     SequenceOfAsciiString from TColStd,    SequenceOfInteger     from TColStd,
     InterfaceModel, Graph, Signature, SignCounter

is

    Create (matcher : Signature;
    	signtext : CString;
    	exact : Boolean = Standard_True)
    	returns mutable SelectSignature;
    ---Purpose : Creates a SelectSignature with its Signature and its Text to
    --           Match.
    --           <exact> if True requires exact match,
    --           if False requires <signtext> to be contained in the Signature
    --           of the entity (default is "exact")

    Create (matcher : Signature;
    	    signtext : AsciiString from TCollection;
    	    exact : Boolean = Standard_True)
    	returns mutable SelectSignature;
    ---Purpose : As above with an AsciiString

    Create (matcher : SignCounter;
    	signtext : CString;
    	exact : Boolean = Standard_True)
    	returns mutable SelectSignature;
    ---Purpose : Creates a SelectSignature with a Counter, more precisely a
    --           SelectSignature. Which is used here to just give a Signature
    --           Value (by SignOnly Mode)
    --           Matching is the default provided by the class Signature

    Signature (me) returns mutable Signature;
    ---Purpose : Returns the used Signature, then it is possible to access it,
    --           modify it as required. Can be null, hence see Counter

    Counter   (me) returns mutable SignCounter;
    ---Purpose : Returns the used SignCounter. Can be used as alternative for
    --           Signature

    SortInGraph (me; rank : Integer; ent : Transient; G : Graph)
    	returns Boolean  is redefined;
    ---Purpose : Returns True for an Entity (model->Value(num)) of which the
    --           signature matches the text given as creation time
    --           May also work with a Counter from the Graph

    Sort (me; rank : Integer; ent : Transient; model : InterfaceModel)
    	returns Boolean;
    ---Purpose : Not called, defined only to remove a deferred method here

    SignatureText (me) returns AsciiString from TCollection;
    ---Purpose : Returns Text used to Sort Entity on its Signature or SignCounter
    ---C++ : return const &

    IsExact (me) returns Boolean;
    ---Purpose : Returns True if match must be exact

    ExtractLabel (me) returns AsciiString from TCollection;
    ---Purpose : Returns a text defining the criterium.
    --           (it refers to the text and exact flag to be matched, and is
    --           qualified by the Name provided by the Signature)

fields

    thematcher  : Signature;
    thecounter  : SignCounter;
    thesigntext : AsciiString from TCollection;
    theexact    : Integer;
    thesignlist : SequenceOfAsciiString from TColStd;
    thesignmode : SequenceOfInteger     from TColStd;

end SelectSignature;
