-- Created on: 1996-02-21
-- Created by: Laurent PAINNOT
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PolygonOnTriangulation from Poly inherits TShared from MMgt

    	---Purpose: This class provides a polygon in 3D space, based on the triangulation
    	-- of a surface. It may be the approximate representation of a
    	-- curve on the surface, or more generally the shape.
    	-- A PolygonOnTriangulation is defined by a table of
    	-- nodes. Each node is an index in the table of nodes specific
    	-- to a triangulation, and represents a point on the surface. If
    	-- the polygon is closed, the index of the point of closure is
    	-- repeated at the end of the table of nodes.
    	-- If the polygon is an approximate representation of a curve
    	-- on a surface, you can associate with each of its nodes the
    	-- value of the parameter of the corresponding point on the
    	-- curve.represents a 3d Polygon 


uses Array1OfInteger  from TColStd,
     Array1OfReal     from TColStd,
     HArray1OfReal    from TColStd,
     Triangulation    from Poly

raises NullObject from Standard

is

    Create(Nodes: Array1OfInteger from TColStd)
    returns mutable PolygonOnTriangulation from Poly;
    	---Purpose: Constructs a 3D polygon on the triangulation of a shape,
    	-- defined by the table of nodes, <Nodes>.
    
    Create(Nodes     : Array1OfInteger from TColStd;
           Parameters: Array1OfReal    from TColStd) 
    returns mutable PolygonOnTriangulation from Poly;
    	---Purpose:
    	-- Constructs a 3D polygon on the triangulation of a shape, defined by:
    	--  -   the table of nodes, Nodes, and the table of parameters, <Parameters>.  
    	-- where:
    	-- -   a node value is an index in the table of nodes specific
    	--   to an existing triangulation of a shape
    	-- -   and a parameter value is the value of the parameter of
    	--   the corresponding point on the curve approximated by
    	--   the constructed polygon.
    	-- Warning
    	-- The tables Nodes and Parameters must be the same size.
    	-- This property is not checked at construction time.
    
    Deflection(me) returns Real;
    	---Purpose: Returns the deflection of this polygon    
    Deflection(me : mutable; D : Real);
    	---Purpose: Sets the deflection of this polygon to D.
 	-- See more on deflection in Poly_Polygones2D.

    NbNodes(me) returns Integer;
	---Purpose:
    	-- Returns the number of nodes for this polygon.
    	-- Note: If the polygon is closed, the point of closure is
    	-- repeated at the end of its table of nodes. Thus, on a closed
    	-- triangle, the function NbNodes returns 4.
    	---C++: inline

    Nodes(me) returns Array1OfInteger from TColStd
	---Purpose: Returns the table of nodes for this polygon. A node value
    	-- is an index in the table of nodes specific to an existing
    	-- triangulation of a shape.
 	---C++: return const &
   raises NullObject from Standard;
    	
    
    HasParameters(me) returns Boolean from Standard;
    	---Purpose:
    	-- Returns true if parameters are associated with the nodes in this polygon.   
    Parameters(me) returns HArray1OfReal from TColStd
    	---	Purpose: Returns the table of the parameters associated with each node in this polygon.
    	-- Warning
    	-- Use the function HasParameters to check if parameters
    	-- are associated with the nodes in this polygon.
	--          
    raises NullObject from Standard;
    
    
fields

    myDeflection    : Real            from Standard;
    myNodes         : Array1OfInteger from TColStd;
    myParameters    : HArray1OfReal   from TColStd;
    
end PolygonOnTriangulation;
