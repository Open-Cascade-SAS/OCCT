-- File:        AutoDesignDateAndPersonAssignment.cdl
-- Created:     Fri Dec  1 11:11:13 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class AutoDesignDateAndPersonAssignment from StepAP214 

inherits PersonAndOrganizationAssignment from StepBasic

uses

	HArray1OfAutoDesignDateAndPersonItem from StepAP214, 
	AutoDesignDateAndPersonItem from StepAP214, 
	PersonAndOrganization from StepBasic,
	PersonAndOrganizationRole from StepBasic
is

	Create returns mutable AutoDesignDateAndPersonAssignment;
	---Purpose: Returns a AutoDesignDateAndPersonAssignment


	Init (me : mutable;
	      aAssignedPersonAndOrganization : mutable PersonAndOrganization from StepBasic;
	      aRole : mutable PersonAndOrganizationRole from StepBasic) is redefined;

	Init (me : mutable;
	      aAssignedPersonAndOrganization : mutable PersonAndOrganization from StepBasic;
	      aRole : mutable PersonAndOrganizationRole from StepBasic;
	      aItems : mutable HArray1OfAutoDesignDateAndPersonItem from StepAP214) is virtual;

	-- Specific Methods for Field Data Access --

	SetItems(me : mutable; aItems : mutable HArray1OfAutoDesignDateAndPersonItem);
	Items (me) returns mutable HArray1OfAutoDesignDateAndPersonItem;
	ItemsValue (me; num : Integer) returns AutoDesignDateAndPersonItem;
	NbItems (me) returns Integer;

fields

	items : HArray1OfAutoDesignDateAndPersonItem from StepAP214; -- a SelectType

end AutoDesignDateAndPersonAssignment;
