-- Created on: 1991-06-24
-- Created by: Didier PIFFAULT
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class Interference from Intf

	---Purpose: Describes the   Interference  computation    result
	--          between polygon2d or polygon3d or polyhedron.

uses    SectionPoint      from Intf,
    	SeqOfSectionPoint from Intf,
    	SectionLine       from Intf,
    	SeqOfSectionLine  from Intf,
    	TangentZone       from Intf,
    	SeqOfTangentZone  from Intf


raises  OutOfRange from Standard


is  Initialize(Self : Boolean from Standard);

    SelfInterference(me   : in out;
    	    	     Self : Boolean from Standard) is protected;
    ---Purpose: Only one argument for the intersection.

    NbSectionPoints(me)
    	    	    returns Integer is static;
    ---Purpose: Gives the number   of  points of  intersection  in the
    --          interference.
    ---C++: inline

    PntValue       (me;
    	    	    Index      : in Integer)
		    returns SectionPoint from Intf
    	    	    raises OutOfRange from Standard
    	    	    is static;
    ---Purpose: Gives the point of  intersection of address  Index in
    --          the interference.
    --
    ---C++: return const &
    ---C++: inline

    NbSectionLines (me)
    	    	    returns Integer is static;
    ---Purpose: Gives the number  of polylines of  intersection in the
    --          interference.
    ---C++: inline

    LineValue      (me;
    	    	    Index      : in Integer)
    	    	    returns SectionLine from Intf
    	    	    raises OutOfRange from Standard
    	    	    is static;
    ---Purpose: Gives the polyline of intersection at address <Index> in
    --          the interference.
    --
    ---C++: return const &
    ---C++: inline

    NbTangentZones  (me)
    	    	    returns Integer is static;
    ---Purpose: Gives the number of zones of tangence in the interference.
    ---C++: inline

    ZoneValue      (me;
    	    	    Index      : in Integer)
    	    	    returns TangentZone from Intf
    	    	    raises OutOfRange from Standard
    	    	    is static;
    ---Purpose: Gives  the zone of  tangence at address   Index in the
    --          interference.
    --
    ---C++: return const &
    ---C++: inline

    GetTolerance   (me)
    	    	    returns Real
    	    	    is static;
    ---Purpose: Gives the tolerance used for the calculation.
    ---C++: inline

-- Implementation functions :

    Contains       (me;
     	    	    ThePnt : in SectionPoint from Intf)
		    returns Boolean
    	    	    is static;
    ---Purpose: Tests if the polylines of  intersection or the zones of
    --          tangence contain the point of intersection <ThePnt>.


    Insert         (me         : in out;
     	    	    TheZone    : in TangentZone from Intf)
		    returns Boolean
    	    	    is static;
    ---Purpose: Inserts a new zone of tangence in  the current list of
    --          tangent zones of  the interference  and  returns  True
    --          when done.


    Insert         (me         : in out;
     	    	    pdeb       : in SectionPoint from Intf;
     	    	    pfin       : in SectionPoint from Intf)
    	    	    is static;
    ---Purpose: Insert a new segment of intersection in the current  list of
    --          polylines of intersection of the interference.


    Dump           (me) is static;


fields    mySPoins  : SeqOfSectionPoint from Intf is protected;
    	  mySLines  : SeqOfSectionLine  from Intf is protected;
    	  myTZones  : SeqOfTangentZone  from Intf is protected;
    	  SelfIntf  : Boolean from Standard is protected;
          Tolerance : Real from Standard is protected;

end Interference;
