-- Created on: 1993-01-11
-- Created by: CKY / Contract Toubro-Larsen (TCD)
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package IGESGraph

        ---Purpose : This package contains the group of classes necessary
        --           to define Graphic data among Structure Entities.
        --           (e.g., Fonts, Colors, Screen management ...)

uses

        Standard,
        TCollection,
        gp,
	TColgp,
	TColStd,
	Message,
        Interface,
        IGESData,
        IGESBasic

is

        class LineFontDefTemplate;

        class LineFontDefPattern;

        class TextFontDef;

        class TextDisplayTemplate;

        class Color;

        class DefinitionLevel;

        class NominalSize;

        class DrawingSize;

        class DrawingUnits;

        class IntercharacterSpacing;

        class LineFontPredefined;

        class HighLight;

        class Pick;

        class UniformRectGrid;

    	--    Tools for Entities    --

        class ToolLineFontDefTemplate;
        class ToolLineFontDefPattern;
        class ToolTextFontDef;
        class ToolTextDisplayTemplate;
        class ToolColor;
        class ToolDefinitionLevel;
        class ToolNominalSize;
        class ToolDrawingSize;
        class ToolDrawingUnits;
        class ToolIntercharacterSpacing;
        class ToolLineFontPredefined;
        class ToolHighLight;
        class ToolPick;
        class ToolUniformRectGrid;

    -- Definition and Exploitation of Entities defined in this Package

    class Protocol;
    class ReadWriteModule;
    class GeneralModule;
    class SpecificModule;

    -- The class instantiations :

    class  Array1OfColor  instantiates   Array1 from TCollection (Color);
    class  Array1OfTextDisplayTemplate instantiates
    	  Array1 from TCollection (TextDisplayTemplate);
    class  Array1OfTextFontDef         instantiates
    	  Array1 from TCollection (TextFontDef);

    class HArray1OfColor  instantiates  HArray1 from TCollection
    	     (Color,Array1OfColor);
    class HArray1OfTextDisplayTemplate instantiates HArray1 from TCollection
    	     (TextDisplayTemplate,Array1OfTextDisplayTemplate);
    class HArray1OfTextFontDef         instantiates HArray1 from TCollection
    	     (TextFontDef,Array1OfTextFontDef);

    -- Package Methods

    Init;
    ---Purpose : Prepares dynamic data (Protocol, Modules) for this package

    Protocol  returns Protocol from IGESGraph;
    ---Purpose : Returns the Protocol for this Package

end IGESGraph;
