-- Created on: 1993-08-11
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PointOnCurve from PBRep inherits PointRepresentation from PBRep
  ---Purpose: Representation by a parameter on a 3D curve.
uses
    Curve    from PGeom,
    Location from PTopLoc

is
    Create(P : Real;
    	   C : Curve    from PGeom;
	   L : Location from PTopLoc)
    returns PointOnCurve from PBRep;
    	---Level: Internal 
    

    Curve(me) returns any Curve from PGeom
    is static;
    	---Level: Internal 

    IsPointOnCurve(me) returns Boolean from Standard
    	---Purpose: Returns True;
    is redefined;
    
fields

    myCurve : Curve from PGeom;

end PointOnCurve;
