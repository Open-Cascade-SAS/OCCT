-- Created on: 1996-11-25
-- Created by: Philippe MANGIN
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class AppFunc from BRepBlend inherits AppFuncRoot from BRepBlend

	---Purpose: Function to approximate by AppSurface
	--          for Surface/Surface contact.
	---Level: Advanced

uses
 Line        from BRepBlend,
 Point       from Blend,
 AppFunction from Blend,
 Function    from Blend,
 Vector      from math
 
raises OutOfRange

is
   Create(Line : in out Line from BRepBlend;
    	  Func : in out Function from Blend;
          Tol3d: Real;
          Tol2d: Real)
   ---Warning: The Object Func cannot be killed before me. 
   returns AppFunc; 

   Point(me;
    	 Func  : AppFunction from Blend; 
	 Param : Real;
	 Sol   : Vector from math;
	 Pnt   : in out Point from Blend);
	
   Vec(me;
       Sol : in out Vector from math;
       Pnt : Point from Blend);
	
end AppFunc;
