-- Created on: 1996-01-26
-- Created by: Christian CAILLET
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class SignValidity  from IFSelect  inherits Signature

    ---Purpose : This Signature returns the Validity Status of an entity, as
    --           deducted from data in the model : it can be
    --           "OK" "Unknown" "Unloaded" "Syntactic Fail"(but loaded)
    --           "Syntactic Warning" "Semantic Fail" "Semantic Warning"


uses CString, Transient, InterfaceModel

is

    Create returns mutable SignValidity;
    ---Purpose : Returns a SignValidity

    CVal  (myclass; ent : any Transient; model : InterfaceModel) returns CString;
    ---Purpose : Returns the Signature for a Transient object, as a validity
    --           deducted from data (reports) stored in the model.
    --           Class method, can be called by any one

    Value (me; ent : any Transient; model : InterfaceModel) returns CString;
    ---Purpose : Returns the Signature for a Transient object, as a validity
    --           deducted from data (reports) stored in the model
    --           Calls the class method CVal

end SignValidity;
