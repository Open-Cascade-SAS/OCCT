-- Created on: 2004-05-11
-- Created by: Sergey ZARITCHNY <szy@opencascade.com>
-- Copyright (c) 2004-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



package BinTools 

	---Purpose: Tool to keep shapes in binary format

uses 
    Geom2d, 
    Geom,
    TColStd,
    TopoDS, 
    TopAbs, 
    TopLoc,
    BRep,
    BRepTools, 
    TopTools
is
    
    class  ShapeSet; 

    class  Curve2dSet; 

    class  CurveSet;  

    class  SurfaceSet; 
     
    class  LocationSet;
    
    pointer LocationSetPtr to LocationSet from BinTools;


    PutReal (OS : out OStream from Standard; theValue : Real from Standard) returns OStream; 
    ---C++: return & 
    
    PutInteger (OS : out OStream from Standard; theValue : Integer from Standard) returns OStream;
    ---C++: return &  

    PutBool (OS : out OStream from Standard; theValue : Boolean from Standard) returns OStream;
    ---C++: return &  

    PutExtChar (OS : out OStream from Standard; theValue : ExtCharacter from Standard) returns OStream;
    ---C++: return &

    GetReal (IS : out IStream from Standard; theValue : out Real from Standard) returns IStream; 
    ---C++: return & 

    GetInteger (IS : out IStream from Standard; theValue : out Integer from Standard) returns IStream; 
    ---C++: return &  
     
    GetBool (IS : out IStream from Standard; theValue : out Boolean from Standard) returns IStream; 
    ---C++: return & 
     
    GetExtChar (IS : out IStream from Standard; theValue : out ExtCharacter from Standard) returns IStream; 
    ---C++: return &

end BinTools;

