-- File:        AreaOrView.cdl
-- Created:     Fri Dec  1 11:11:10 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993



class AreaOrView from StepVisual inherits SelectType from StepData

	-- <AreaOrView> is an EXPRESS Select Type construct translation.
	-- it gathers : PresentationArea, PresentationView

uses

	PresentationArea,
	PresentationView
is

	Create returns AreaOrView;
	---Purpose : Returns a AreaOrView SelectType

	CaseNum (me; ent : Transient) returns Integer;
	---Purpose: Recognizes a AreaOrView Kind Entity that is :
	--        1 -> PresentationArea
	--        2 -> PresentationView
	--        0 else

	PresentationArea (me) returns any PresentationArea;
	---Purpose : returns Value as a PresentationArea (Null if another type)

	PresentationView (me) returns any PresentationView;
	---Purpose : returns Value as a PresentationView (Null if another type)


end AreaOrView;

