-- Created on: 2007-05-29
-- Created by: Vlad Romashko
-- Copyright (c) 2007-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class BooleanList from TDataStd inherits Attribute from TDF

    ---Purpose: Contains a list of bolleans.

uses 

    Attribute from TDF,
    GUID from Standard,
    Label from TDF,
    RelocationTable from TDF,
    ListOfByte from TDataStd

is 

    ---Purpose: Static methods
    --          ==============

    GetID (myclass)   
    ---C++: return const & 
    ---Purpose: Returns the ID of the list of booleans attribute.
    returns GUID from Standard;

    Set (myclass; label : Label from TDF)
    ---Purpose: Finds or creates a list of boolean values attribute.
    returns BooleanList from TDataStd;

    
    ---Category: BooleanList methods
    --           ===================

    Create
    returns BooleanList from TDataStd; 

    IsEmpty (me)
    returns Boolean from Standard;
    
    Extent (me)
    returns Integer from Standard;
    
    Prepend (me : mutable;
    	     value : Boolean from Standard);

    Append (me : mutable;
    	    value : Boolean from Standard);
    
    Clear (me : mutable);
    
    First (me)
    returns Boolean from Standard;
    
    Last (me)
    returns Boolean from Standard;

    List (me)
    ---C++: return const &
    ---Purpose: 1 - means TRUE,
    --          0 - means FALSE.
    returns ListOfByte from TDataStd;
    
    
    ---Category: Methodes of TDF_Attribute
    --           =========================
    
    ID (me)
    ---C++: return const & 
    returns GUID from Standard;

    Restore (me: mutable; With : Attribute from TDF);

    NewEmpty (me)
    returns Attribute from TDF;

    Paste (me; Into : Attribute from TDF;
	       RT   : RelocationTable from TDF);    
    
    Dump(me; anOS : in out OStream from Standard)
    returns OStream from Standard
    is redefined;
    ---C++: return &


fields

    myList : ListOfByte from TDataStd;


end BooleanList;
