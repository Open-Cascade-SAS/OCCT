-- Created on: 1997-06-06
-- Created by: Alexander BRIVIN
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Projector from VrmlConverter inherits TShared from MMgt

	---Purpose: 
    	--     defines projector  and calculates properties of cameras and lights from Vrml
	--     ( OrthograpicCamera, PerspectiveCamera, DirectionalLight, PointLight, SpotLight  
    	--     and  MatrixTransform  )  to display all scene  shapes  with  arbitrary locations 
	--     for requested the Projection Vector,  High Point Direction and the Focus
	--     and adds them ( method Add ) to anOSream.

uses
 
    Projector from HLRAlgo,
    Array1OfShape  from  TopTools, 
    Length    from Quantity,
    PerspectiveCamera  from Vrml, 
    OrthographicCamera  from Vrml, 
    DirectionalLight  from  Vrml, 
    PointLight  from Vrml,
    SpotLight  from Vrml,
    TypeOfCamera from VrmlConverter, 
    TypeOfLight from VrmlConverter,
    MatrixTransform  from Vrml

is

    Create ( Shapes:  Array1OfShape from TopTools; 
    	     Focus: Length from Quantity;        
	     DX, DY, DZ: Length from Quantity;                             -- Projection Vector
	     XUp, YUp, ZUp: Length from Quantity;                          -- High Point Direction
	     Camera:  TypeOfCamera from VrmlConverter  = VrmlConverter_NoCamera;
   	     Light:   TypeOfLight from VrmlConverter   = VrmlConverter_NoLight ) 
    returns mutable Projector from VrmlConverter; 
    

    SetCamera ( me: mutable; aCamera : TypeOfCamera from VrmlConverter );
    Camera ( me )  returns  TypeOfCamera from VrmlConverter;
    
    SetLight ( me: mutable; aLight : TypeOfLight from VrmlConverter );
    Light ( me )  returns  TypeOfLight from VrmlConverter;


    Add(me;   anOStream: in out OStream from Standard);
    	---Purpose:  
        --    Adds  into anOStream  if  they  are  defined in  Create.
    	--      PerspectiveCamera,
    	--      OrthographicCamera, 
    	--      DirectionLight,
    	--      PointLight,
    	--      SpotLight 
        --   with  MatrixTransform  from VrmlConverter;
 
      
    Projector(me) returns Projector from HLRAlgo
    is static;
				       
fields
 
    myProjector:           Projector          from HLRAlgo;
    myPerspectiveCamera:   PerspectiveCamera  from Vrml; 
    myOrthographicCamera:  OrthographicCamera from Vrml; 
    myDirectionalLight:    DirectionalLight   from Vrml; 
    myPointLight:          PointLight         from Vrml;
    mySpotLight:           SpotLight          from Vrml;
    myTypeOfCamera:    	   TypeOfCamera       from VrmlConverter;
    myTypeOfLight:    	   TypeOfLight        from VrmlConverter;
    myMatrixTransform:     MatrixTransform    from Vrml;

end Projector;


