-- File:	StepData_EnumTool.cdl
-- Created:	Wed Oct 25 10:49:31 1995
-- Author:	Christian CAILLET
--		<cky@anion>
---Copyright:	 Matra Datavision 1995


class EnumTool  from StepData

    ---Purpose : This class gives a way of conversion between the value of an
    --           enumeration and its representation in STEP
    --           An enumeration corresponds to an integer with reserved values,
    --           which begin to 0
    --           In STEP, it is represented by a name in capital letter and
    --           limited by two dots, e.g. .UNKNOWN.
    --           
    --           EnumTool works with integers, it is just required to cast
    --           between an integer and an enumeration of required type.
    --           
    --           Its definition is intended to allow static creation in once,
    --           without having to recreate once for each use.
    --           
    --           It is possible to define subclasses on it, which directly give
    --           the good list of definition texts, and accepts a enumeration
    --           of the good type instead of an integer

uses CString, AsciiString, SequenceOfAsciiString

is

    Create (e0,e1,e2,e3,e4,e5,e6,e7,e8,e9,e10,e11,e12,e13,e14,e15,e16,e17,e18,e19,e20,e21,e22,e23,e24,e25,e26,e27,e28,e29,e30,e31,e32,e33,e34,e35,e36,e37,e38,e39 : CString = "")
    	returns EnumTool;
    ---Purpose : Creates an EnumTool with definitions given by e0 .. e<max>
    --           Each definition string can bring one term, or several
    --           separated by blanks. Each term corresponds to one value of the
    --           enumeration, if dots are not presents they are added
    --           
    --           Such a static constructor allows to build a static description
    --            as : static StepData_EnumTool myenumtool("e0","e1"...);
    --            then use it without having to initialise it
    --           
    --           A null definition can be input by given "$" :the corresponding
    --           position is attached to "null/undefined" value (as one
    --           particular item of the enumeration list)

    AddDefinition (me : in out; term : CString);
    ---Purpose : Processes a definition, splits it according blanks if any
    --           empty definitions are ignored
    --           A null definition can be input by given "$" :the corresponding
    --           position is attached to "null/undefined" value (as one
    --           particular item of the enumeration list)
    --           See also IsSet

    IsSet (me) returns Boolean;
    ---Purpose : Returns True if at least one definition has been entered after
    --           creation time (i.e. by AddDefinition only)
    --           
    --           This allows to build a static description by a first pass :
    --           static StepData_EnumTool myenumtool("e0" ...);
    --           ...
    --           if (!myenumtool.IsSet()) {             for further inits
    --             myenumtool.AddDefinition("e21");
    --             ...
    --           }

    MaxValue (me) returns Integer;
    ---Purpose : Returns the maximum integer for a suitable value
    --           Remark : while values begin at zero, MaxValue is the count of
    --           recorded values minus one

    Optional (me : in out; mode : Boolean);
    ---Purpose : Sets or Unsets the EnumTool to accept undefined value (for
    --           optional field). Ignored if no null value is defined (by "$")
    --           Can be changed during execution (to read each field),
    --           Default is True (if a null value is defined)

    NullValue (me) returns Integer;
    ---Purpose : Returns the value attached to "null/undefined value"
    --           If none is specified or if Optional has been set to False,
    --             returns -1
    --           Null Value has been specified by definition "$"

    Text (me; num : Integer) returns AsciiString;
    ---Purpose : Returns the text which corresponds to a given numeric value
    --           It is limited by dots
    --           If num is out of range, returns an empty string
    ---C++ : return const &

    Value (me; txt : CString) returns Integer;
    ---Purpose : Returns the numeric value found for a text
    --           The text must be in capitals and limited by dots
    --           A non-suitable text gives a negative value to be returned

    Value (me; txt : AsciiString) returns Integer;
    ---Purpose : Same as above but works on an AsciiString

fields

    thetexts : SequenceOfAsciiString;
    theinit  : Integer;
    theopt   : Boolean;

end EnumTool;
