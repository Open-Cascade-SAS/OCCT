-- Created on: 2002-12-12
-- Created by: data exchange team
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class FeaParametricPoint from StepFEA
inherits Point from StepGeom

    ---Purpose: Representation of STEP entity FeaParametricPoint

uses
    HAsciiString from TCollection,
    HArray1OfReal from TColStd

is
    Create returns FeaParametricPoint from StepFEA;
	---Purpose: Empty constructor

    Init (me: mutable; aRepresentationItem_Name: HAsciiString from TCollection;
                       aCoordinates: HArray1OfReal from TColStd);
	---Purpose: Initialize all fields (own and inherited)

    Coordinates (me) returns HArray1OfReal from TColStd;
	---Purpose: Returns field Coordinates
    SetCoordinates (me: mutable; Coordinates: HArray1OfReal from TColStd);
	---Purpose: Set field Coordinates

fields
    theCoordinates: HArray1OfReal from TColStd;

end FeaParametricPoint;
