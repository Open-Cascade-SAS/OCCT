-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class LoopAndPath from StepShape 

inherits TopologicalRepresentationItem from StepShape 


	--- This classe is an implementation of EXPRESS
	--  ANDOR Subtype Declaration.
uses

	Loop from StepShape, 
	Path from StepShape, 
	HAsciiString from TCollection, 
	HArray1OfOrientedEdge from StepShape, 
	OrientedEdge from StepShape
is

	Create returns LoopAndPath;
	---Purpose: Returns a LoopAndPath


	Init (me : mutable;
	      aName : HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      aName : HAsciiString from TCollection;
	      aLoop : Loop from StepShape;
	      aPath : Path from StepShape) is virtual;

	Init (me : mutable;
	      aName : HAsciiString from TCollection;
	      aEdgeList : HArray1OfOrientedEdge from StepShape) is virtual;

	-- Specific Methods for Field Data Access --

	SetLoop(me : mutable; aLoop : Loop);
	Loop (me) returns Loop;
	SetPath(me : mutable; aPath : Path);
	Path (me) returns Path;

	-- Specific Methods for ANDOR Field Data Access --


	-- Specific Methods for ANDOR Field Data Access --

	SetEdgeList(me : mutable; aEdgeList : HArray1OfOrientedEdge);
	EdgeList (me) returns HArray1OfOrientedEdge;
	EdgeListValue (me; num : Integer) returns OrientedEdge;
	NbEdgeList (me) returns Integer;

fields

	loop : Loop from StepShape;
	path : Path from StepShape;

end LoopAndPath;
