-- Created on: 1993-11-03
-- Created by: Christian CAILLET
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SelectSharing  from IFSelect  inherits SelectDeduct

    ---Purpose : A SelectSharing selects Entities which directly Share (Level
    --           One) the Entities of the Input list
    --           Remark : if an Entity of the Input List directly shares
    --           another one, it is of course present in the Result List

uses AsciiString from TCollection, EntityIterator, Graph

is

    Create returns SelectSharing;
    ---Purpose : Creates a SelectSharing;

    RootResult (me; G : Graph) returns EntityIterator;
    ---Purpose : Returns the list of selected entities (list of entities
    --           which share (level one) those of input list)

    Label (me) returns AsciiString from TCollection;
    ---Purpose : Returns a text defining the criterium : "Sharing (one level)"

end SelectSharing;
