-- Created on: 1997-02-10
-- Created by: Robert COUBLANC
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

--   GG  :  GER61351 17/11/1999 Change SetColor() with a compatible Quantity_Color instead
--                                     the restricted NameOfColor.

class GraphicTool from AIS 

	---Purpose: 

uses
    Drawer          from Prs3d,
    TypeOfAttribute from AIS,
    NameOfColor     from Quantity,
    Color     	    from Quantity,
    TypeOfLine      from Aspect,
    MaterialAspect  from Graphic3d


is

    GetLineColor(myclass; aDrawer : Drawer from Prs3d; TheTypeOfAttributes :  TypeOfAttribute  from  AIS) 
    returns NameOfColor from Quantity; 
    
    GetLineColor(myclass; aDrawer : Drawer from Prs3d; 
		TheTypeOfAttributes :  TypeOfAttribute  from  AIS;
		TheLineColor: out Color from Quantity);
    
    GetLineWidth(myclass; aDrawer : Drawer from Prs3d; TheTypeOfAttributes :  TypeOfAttribute  from  AIS)
    returns Real from Standard;
    
    
    GetLineType (myclass; aDrawer : Drawer from Prs3d; TheTypeOfAttributes :  TypeOfAttribute  from  AIS)  
    returns TypeOfLine from Aspect;
    
    
    GetLineAtt(myclass;
    	       aDrawer : Drawer from Prs3d;
    	       TheTypeOfAttributes :  TypeOfAttribute  from  AIS; 
    	       aCol   : in out NameOfColor from Quantity;
	       aWidth : in out Real from Standard;
	       aTyp   : in out TypeOfLine from Aspect);
	       
	       
    GetInteriorColor(myclass;
    	    	    aDrawer : Drawer from Prs3d) 
    returns NameOfColor from  Quantity;

    GetInteriorColor(myclass;
    	    	    aDrawer : Drawer from Prs3d;
		    aColor: out Color from Quantity);

    GetMaterial(myclass; aDrawer:Drawer from Prs3d)
    returns MaterialAspect from Graphic3d;
	       
end GraphicTool;

