-- File:	PGeom2d_Curve.cdl
-- Created:	Tue Apr  6 17:20:21 1993
-- Author:	Philippe DAUTRY
--		<fid@mastox>
-- Copyright:	 Matra Datavision 1993


deferred class Curve from PGeom2d inherits Geometry from PGeom2d

         --- Purpose :
         --  Defines the general abstract class curve in the 3D space.
         --  
	 ---See Also : Curve from Geom2d.

is

end;
