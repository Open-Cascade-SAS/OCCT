-- Created on: 1993-01-11
-- Created by: CKY / Contract Toubro-Larsen ( Anand NATRAJAN )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class PWBDrilledHole from IGESAppli  inherits IGESEntity

        ---Purpose: defines PWBDrilledHole, Type <406> Form <26>
        --          in package IGESAppli
        --          Used to identify an entity that locates a drilled hole
        --          and to specify the characteristics of the drilled hole

uses  Integer, Real  -- no one specific type

is

        Create returns mutable PWBDrilledHole;

        -- Specific Methods pertaining to the class

        Init (me         : mutable;
              nbPropVal  : Integer;
              aDrillDia  : Real;
              aFinishDia : Real;
              aCode      : Integer);
        ---Purpose : This method is used to set the fields of the class
        --           PWBDrilledHole
        --       - nbPropVal  : number of property values, always = 3
        --       - aDrillDia  : Drill diameter size
        --       - aFinishDia : Finish diameter size
        --       - aCode      : Function code for drilled hole

        NbPropertyValues (me) returns Integer;
        ---Purpose : returns number of property values, always = 3

        DrillDiameterSize (me) returns Real;
        ---Purpose : returns Drill diameter size

        FinishDiameterSize (me) returns Real;
        ---Purpose : returns Finish diameter size

        FunctionCode (me) returns Integer;
        ---Purpose : returns Function code for drilled hole
        -- is 0, 1, 2, 3, 4, 5 or 5001-9999

fields

--
-- Class    : IGESAppli_PWBDrilledHole
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class PWBDrilledHole.
--
-- Reminder : A PWBDrilledHole instance is defined by :
--            - number of property values, always = 3
--            - Drill diameter size
--            - Finish diameter size
--            - Function code for drilled hole

        theNbPropertyValues : Integer;
        theDrillDiameter    : Real;
        theFinishDiameter   : Real;
        theFunctionCode     : Integer;

end PWBDrilledHole;
