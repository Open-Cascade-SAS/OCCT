-- Created on: 1996-12-24
-- Created by: Alexander BRIVIN
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Cone from Vrml 

	---Purpose: defines a Cone node of VRML specifying geometry shapes.
    	-- This  node  represents  a  simple  cone,  whose  central  axis  is  aligned 
	-- with  the  y-axis.  By  default ,  the  cone  is  centred  at  (0,0,0) 
	-- and  has  size  of  -1  to  +1  in  the  all  three  directions. 
	-- the  cone  has  a  radius  of  1  at  the  bottom  and  height  of  2, 
	-- with  its  apex  at  1  and  its  bottom  at  -1.  The  cone  has  two  parts: 
	-- the  sides  and  the  bottom
uses
     
    ConeParts from Vrml
is

    Create ( aParts        : ConeParts from Vrml = Vrml_ConeALL; 
    	     aBottomRadius : Real      from Standard = 1; 
             aHeight       : Real      from Standard = 2 )  
        returns Cone from Vrml;
    
    SetParts ( me : in out; aParts : ConeParts from Vrml );
    Parts ( me )  returns  ConeParts from Vrml;

    SetBottomRadius ( me : in out; aBottomRadius : Real from Standard );
    BottomRadius ( me )  returns Real  from  Standard;

    SetHeight ( me : in out; aHeight : Real from Standard );
    Height ( me )  returns Real  from  Standard;

    Print  ( me;  anOStream: in out OStream from Standard) returns OStream from Standard;
    ---C++:  return  & 

fields

    myParts        : ConeParts from Vrml;      -- Visible parts of cone
    myBottomRadius : Real      from Standard;  -- Radius of bottom circular face
    myHeight       : Real      from Standard;  -- Size in y dimension
   
end Cone;
