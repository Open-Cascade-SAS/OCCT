-- Created on: 2000-08-11
-- Created by: Andrey BETENEV
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class AISObject from XCAFPrs inherits Shape from AIS

    ---Purpose: Implements AIS_InteractiveObject functionality
    --          for shape in DECAF document

uses
    Shape from TopoDS,
    PresentationManager3d from PrsMgr,
    Presentation from Prs3d,
    Label from TDF,
    Color from Quantity,
    NameOfMaterial from Graphic3d,
    MaterialAspect from Graphic3d,
    Style from XCAFPrs
    
is

    Create (lab: Label from TDF);
    	---Purpose: Creates an object to visualise the shape label

    SetColor(me:mutable;aColor:Color from Quantity) is redefined virtual;

    UnsetColor(me:mutable) is redefined virtual;
        
    SetMaterial(me:mutable;aName:NameOfMaterial from Graphic3d) is redefined virtual;

    SetMaterial(me:mutable;aName:MaterialAspect from Graphic3d) is redefined virtual;
        
    UnsetMaterial(me:mutable) is redefined virtual;
        
    SetTransparency(me:mutable;aValue : Real from Standard=0.6) is redefined virtual;  
    
    UnsetTransparency(me:mutable) is redefined virtual;
 
    AddStyledItem (me: mutable; style: Style from XCAFPrs;
                   shape: Shape from TopoDS;
                   aPresentationManager : PresentationManager3d from PrsMgr;
                   aPresentation        : mutable Presentation from Prs3d;
    	           aMode                : Integer from Standard = 0) 
    is private;

    Compute (me                   : mutable;
             aPresentationManager : PresentationManager3d from PrsMgr;
             aPresentation        : mutable Presentation from Prs3d;
    	     aMode                : Integer from Standard = 0) 
    is redefined virtual protected;
    	---Purpose: Redefined method to compute presentation

    DefaultStyle (me;
                  aStyle: out Style from XCAFPrs)
    is virtual protected;
    ---Purpose: Fills out a default style object which is used when styles are
    --          not explicitly defined in the document.
    --          By default, the style uses white color for curves and surfaces.

fields
    myLabel : Label from TDF;

end AISObject;
