-- Created on: 2007-05-29
-- Created by: Vlad Romashko
-- Copyright (c) 2007-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class IntegerList from TDataStd inherits Attribute from TDF

    ---Purpose: Contains a list of integers.

uses 

    Attribute from TDF,
    GUID from Standard,
    Label from TDF,
    RelocationTable from TDF,
    ListOfInteger from TColStd

is 

    ---Purpose: Static methods
    --          ==============

    GetID (myclass)   
    ---C++: return const & 
    ---Purpose: Returns the ID of the list of integer attribute.
    returns GUID from Standard;

    Set (myclass; label : Label from TDF)
    ---Purpose: Finds or creates a list of integer values attribute.
    returns IntegerList from TDataStd;

    
    ---Category: IntegerList methods
    --           ===================

    Create
    returns mutable IntegerList from TDataStd; 

    IsEmpty (me)
    returns Boolean from Standard;
    
    Extent (me)
    returns Integer from Standard;
    
    Prepend (me : mutable;
    	     value : Integer from Standard);
	     
    Append (me : mutable;
    	    value : Integer from Standard);
	    
    InsertBefore (me : mutable;
    	    	  value : Integer from Standard;
		  before_value : Integer from Standard)
    ---Purpose: Inserts the <value> before the first meet of <before_value>.
    returns Boolean from Standard;

    InsertAfter (me : mutable;
    	    	 value : Integer from Standard;
		 after_value : Integer from Standard)
    ---Purpose: Inserts the <value> after the first meet of <after_value>.
    returns Boolean from Standard;

    Remove (me : mutable;
    	    value : Integer from Standard)
    ---Purpose: Removes the first meet of the <value>.
    returns Boolean from Standard;
    
    Clear (me : mutable);
    
    First (me)
    returns Integer from Standard;
    
    Last (me)
    returns Integer from Standard;

    List (me)
    ---C++: return const &
    returns ListOfInteger from TColStd;
    
    ---Category: Methodes of TDF_Attribute
    --           =========================
    
    ID (me)
    ---C++: return const & 
    returns GUID from Standard;

    Restore (me: mutable; With : Attribute from TDF);

    NewEmpty (me)
    returns mutable Attribute from TDF;

    Paste (me; Into : mutable Attribute from TDF;
	       RT   : mutable RelocationTable from TDF);    
    
    Dump(me; anOS : in out OStream from Standard)
    returns OStream from Standard
    is redefined;
    ---C++: return &


fields

    myList : ListOfInteger from TColStd;


end IntegerList;
