-- File:	RWStepDimTol_RWRoundnessTolerance.cdl
-- Created:	Wed Jun  4 13:34:34 2003 
-- Author:	Galina KULIKOVA
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWRoundnessTolerance from RWStepDimTol

    ---Purpose: Read & Write tool for RoundnessTolerance

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    RoundnessTolerance from StepDimTol

is
    Create returns RWRoundnessTolerance from RWStepDimTol;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : RoundnessTolerance from StepDimTol);
	---Purpose: Reads RoundnessTolerance

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: RoundnessTolerance from StepDimTol);
	---Purpose: Writes RoundnessTolerance

    Share (me; ent : RoundnessTolerance from StepDimTol;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWRoundnessTolerance;
