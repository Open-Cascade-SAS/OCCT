-- Created on: 1997-03-26
-- Created by: Christian CAILLET
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class AutoDesignPresentedItemSelect from StepAP214 inherits SelectType from StepData

	-- <AutoDesignPresentedItemSelect> is an EXPRESS Select Type construct translation.
	-- it gathers : ProductDefinition, ProductDefinitionShape, RepresentationRelationship, ShapeAspect

uses
     ProductDefinition from StepBasic,
     ProductDefinitionRelationship from StepBasic,
     ProductDefinitionShape from StepRepr,
     RepresentationRelationship from StepRepr,
     ShapeAspect from StepRepr,
     DocumentRelationship from StepBasic

is

	Create returns AutoDesignPresentedItemSelect;
	---Purpose : Returns a AutoDesignPresentedItemSelect SelectType

	CaseNum (me; ent : Transient) returns Integer;
	---Purpose: Recognizes a AutoDesignPresentedItemSelect Kind Entity that is :
	--  1 -> ProductDefinition,
	--  2 -> ProductDefinitionRelationship,
	--  3 -> ProductDefinitionShape
	--  4 -> RepresentationRelationship
	--  5 -> ShapeAspect
	--  6 -> DocumentRelationship,
	--        0 else

    ProductDefinitionRelationship (me) returns any ProductDefinitionRelationship;
    ---Purpose : returns Value as a ProductDefinitionRelationship (Null if another type)

    ProductDefinition (me) returns any ProductDefinition;
    ---Purpose : returns Value as a ProductDefinition (Null if another type)

    ProductDefinitionShape (me) returns any ProductDefinitionShape;
    ---Purpose : returns Value as a ProductDefinitionShape (Null if another type)

    RepresentationRelationship (me) returns any RepresentationRelationship;
    ---Purpose : returns Value as a RepresentationRelationship (Null if another type)

    ShapeAspect (me) returns any ShapeAspect;
    ---Purpose : returns Value as a ShapeAspect (Null if another type)

    DocumentRelationship (me) returns any DocumentRelationship;
    ---Purpose : returns Value as a DocumentRelationship (Null if another type)

end AutoDesignPresentedItemSelect;
