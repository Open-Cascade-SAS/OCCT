-- Created on: 1995-11-28
-- Created by: Jean-Pierre COMBE
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class PerpenPresentation from DsgPrs

        ---Purpose: A framework to define display of perpendicular
    	-- constraints between shapes.
uses
    Presentation from Prs3d,
    Pnt from gp,
    Dir from gp,
    Drawer from Prs3d,
    ExtendedString from TCollection
    	
is  
    Add( myclass; aPresentation: Presentation from Prs3d;
    	    	  aDrawer: Drawer from Prs3d;
    	    	  pAx1:          Pnt from gp;
		  pAx2:          Pnt from gp;
                  pnt1:          Pnt from gp;
		  pnt2:          Pnt from gp;
		  OffsetPoint:   Pnt from gp;
    	    	  intOut1:       Boolean from Standard;
    	    	  intOut2:       Boolean from Standard);
	---Purpose: Defines the display of elements showing
    	-- perpendicular constraints between shapes.
    	-- These include the two axis points pAx1 and pAx2,
    	-- the two points pnt1 and pnt2, the offset point
    	-- OffsetPoint and the two Booleans intOut1} and intOut2{.
    	-- These arguments are added to the presentation
    	-- object aPresentation. Their display attributes are
    	-- defined by the attribute manager aDrawer.


end PerpenPresentation;
