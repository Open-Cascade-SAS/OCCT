-- Created on: 1991-02-21
-- Created by: Isabelle GRIGNON
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class   POnSurf from Extrema
    	---Purpose: Definition of a point on surface.

uses    Pnt from gp

is
    Create returns POnSurf;
    	---Purpose: Creation of an indefinite point on surface.
    	---C++: inline

    Create (U,V: Real; P: Pnt) returns POnSurf;
    	---Purpose: Creation of a point on surface with parameter 
    	--          values on the surface and a Pnt from gp.
    	---C++: inline

    Value (me) returns Pnt
    	---Purpose: Returns the 3d point.
    	---C++: return const&
    	---C++: inline
    	is static;

    Parameter (me; U,V: out Real) 
    	---Purpose: Returns the parameter values on the surface.
    	---C++: inline
    	is static;          
    
fields
    myU: Real;
    myV: Real;
    myP: Pnt from gp;

end POnSurf;
