-- Created on: 1991-09-06
-- Created by: Denis PASCAL
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

generic class RelationGraph from GraphDS 
             (GraphDS_Item      as any;
              GraphDS_Attribute as any)
		     
    ---Purpose: This  generic class describe  a  network (or graph) of
    --          Relations between Entities.  an Item can be associated
    --          to the  Entity and respectively  an  Attribute  to the
    --          Relation.   This  class can     be compared   to   the
    --          DirectedGraph of this package.   But here the Relation
    --          (compared to the Edge) can describe links between more
    --          than two  Entities.   Each  link can  be described  as
    --          oriented or  not.  Nested  classes permit to  edit and
    --          visit that structure.  Interface of visiting tools are
    --          done as iterators.


uses  TShared        from MMgt,
      MapOfTransient from TColStd,
      EntityRole     from GraphDS

raises NoSuchObject from Standard, 
       NoMoreObject from Standard,
       DomainError  from Standard

    class Entity from GraphDS inherits TShared from MMgt
    
    uses RelationRole   from GraphDS,
         MapOfTransient from TColStd
    
    is
    
    	Create (value : GraphDS_Item) 
    	returns mutable Entity from GraphDS;

       	GetItem (me)            
    	---Level: Internal
	---C++ : return const& 
    	returns any GraphDS_Item;

	Contains (me; R : Relation from GraphDS)  
    	---Level: Internal
        returns Boolean from Standard;

    	HasRelation (me)  
    	---Level: Internal 
    	returns Boolean from Standard;
	
    	GetRole (me; R : Relation from GraphDS)  
    	---Level: Internal
	returns RelationRole from GraphDS;
	
        IsFront (me; R : Relation from GraphDS)  
    	---Level: Internal 
    	returns Boolean from Standard;
  
        IsBack (me; R : Relation from GraphDS)  
    	---Level: Internal 
    	returns Boolean from Standard;

    	Add (me : mutable; R : Relation from GraphDS)
	is private;

    	Remove (me : mutable; R : Relation from GraphDS)
        is private;
	
    	GetRelations (me)
	---C++: return const&
	returns MapOfTransient from TColStd
	is private;

    fields

    	myItem      : GraphDS_Item;  
    	myRelations : MapOfTransient from TColStd;

    friends

        class RelationGraph from GraphDS,
    	class EntitiesIterator          from GraphDS,
	class IncidentEntitiesIterator  from GraphDS,
    	class RelationsIterator         from GraphDS,	
	class IncidentRelationsIterator from GraphDS

    end Entity from GraphDS;

		
    class Relation inherits TShared from MMgt

    uses EntityRole    from GraphDS,
         EntityRoleMap from GraphDS
    
    is

    	Create (value : GraphDS_Attribute) 
    	returns mutable Relation;

       	GetAttribute (me)             
    	---Level: Internal
	---C++: return const&
    	returns any GraphDS_Attribute;

	Contains (me; E : Entity from GraphDS)   
    	---Level: Internal
    	returns Boolean from Standard;

    	IsEmpty (me) 
    	---Level: Internal
    	returns Boolean from Standard;
	
	GetRole (me; E : Entity from GraphDS)  
    	---Level: Internal
	returns EntityRole from GraphDS;

        IsInput (me; E : Entity from GraphDS) 
    	 ---Level: Internal
	returns Boolean from Standard;
	
        IsOutput (me; E : Entity from GraphDS)
    	---Level: Internal
	returns Boolean from Standard;
	
	Remove   (me : mutable; E : Entity from GraphDS)
	is private;
	
        Add      (me : mutable; E : Entity from GraphDS; 
                                R : EntityRole from GraphDS)
	is private;			
	
	SetRole  (me : mutable; E : Entity from GraphDS;
	                        R : EntityRole from GraphDS)
	is private;			
	
    	GetEntities (me) 
	---C++: return const&
    	returns EntityRoleMap from GraphDS
	is private;
	
    fields

    	myAttribute : GraphDS_Attribute;  
	myEntities  : EntityRoleMap from GraphDS;

    friends	

    	class RelationGraph             from GraphDS,
    	class EntitiesIterator          from GraphDS,
	class IncidentEntitiesIterator  from GraphDS,
	class RelationsIterator         from GraphDS,	
	class IncidentRelationsIterator from GraphDS
	
    end Relation;


    class EntitiesIterator from GraphDS 

    	---Purpose: Public nested class which  defines an  iterator to
    	--          visit each Entity member of a given RelationGraph.

    uses MapOfTransient from TColStd,
         MapIteratorOfMapOfTransient from TColStd
    
    raises NoMoreObject from Standard,
           NoSuchObject from Standard
    is

    	Create 
    	returns EntitiesIterator from GraphDS;
	
	Create (G : RelationGraph from GraphDS)
    	returns EntitiesIterator from GraphDS;
	
	Create (G : RelationGraph from GraphDS;
	        E : Entity        from GraphDS)
    	returns EntitiesIterator from GraphDS;
	
	Create (G : RelationGraph from GraphDS;
	        E : Relation      from GraphDS)
    	returns EntitiesIterator from GraphDS;
	
    	Initialize (me : in out; G : RelationGraph from GraphDS);
            ---Level: Public

    	Initialize (me : in out; G : RelationGraph from GraphDS;
	                         E : Entity        from GraphDS);
            ---Level: Public
	
    	Initialize (me : in out; G : RelationGraph from GraphDS; 
 	                         R : Relation      from GraphDS);
            ---Level: Public

    	More (me)   
    	---Level: Public
    	returns Boolean from Standard;

    	Next (me : in out)   
    	---Level: Public 
    	raises NoMoreObject from Standard;

    	Value (me) 
    	---C++: return const&
    	---Level: Public 
    	returns Entity from GraphDS
    	raises NoSuchObject from Standard;

    fields

    	myMap      : MapOfTransient from TColStd;
    	myEntities : MapIteratorOfMapOfTransient from TColStd;

    end EntitiesIterator;


    class RelationsIterator from GraphDS 

    	---Purpose: Public nested  class which defines  an iterator to
    	--          visit   each  Relation    member   of  a     given
    	--          RelationGraph.

    uses MapOfTransient from TColStd,
         MapIteratorOfMapOfTransient from TColStd

    raises NoMoreObject from Standard,
           NoSuchObject from Standard
    is 
    
    	Create
        returns RelationsIterator from GraphDS;
	
	Create (G : RelationGraph from GraphDS)
        returns RelationsIterator from GraphDS;
	
	Create (G : RelationGraph from GraphDS;
	        R : Relation      from GraphDS)
        returns RelationsIterator from GraphDS;
	
	Create (G : RelationGraph from GraphDS;
	        E : Entity        from GraphDS)
        returns RelationsIterator from GraphDS;	
	
	Initialize (me : in out; G : RelationGraph from GraphDS);
            ---Level: Public

    	Initialize (me : in out; G : RelationGraph from GraphDS; 
                                 R : Relation      from GraphDS);
            ---Level: Public
	
    	Initialize (me : in out; G : RelationGraph from GraphDS; 
                                 E : Entity        from GraphDS);
            ---Level: Public
	
    	More (me) 
    	returns Boolean from Standard;
            ---Level: Public
	
    	Next (me : in out) 
    	raises NoMoreObject from Standard;
            ---Level: Public
	
    	Value (me) 
    	---C++: return const&
    	returns Relation from GraphDS
        raises NoSuchObject from Standard;
            ---Level: Public
	
    fields
    
     	myMap       : MapOfTransient from TColStd;
        myRelations : MapIteratorOfMapOfTransient from TColStd;
	
    end RelationsIterator;


    class IncidentEntitiesIterator from GraphDS
    
    uses MapOfTransient from TColStd,
         MapIteratorOfMapOfTransient from TColStd
    
    raises NoMoreObject from Standard,
           NoSuchObject from Standard

    is 

    	Create 
        returns IncidentEntitiesIterator from GraphDS;
	
	Create (G : RelationGraph from GraphDS; 
    	        E : Entity        from GraphDS) 
        returns IncidentEntitiesIterator from GraphDS;

    	Initialize (me : in out; G : RelationGraph from GraphDS; 
    	                         E : Entity        from GraphDS); 
        ---Level: Public
	
	More (me)  
    	---Level: Public
    	returns Boolean from Standard;
	
    	Next (me : in out)
    	---Level: Public 
    	raises NoMoreObject from Standard;
	
    	Value (me) 
    	---C++: return const&  
    	---Level: Public
    	returns Entity from GraphDS 
        raises NoSuchObject from Standard;
	
    fields
    
    	myMap      : MapOfTransient from TColStd;
    	myEntities : MapIteratorOfMapOfTransient from TColStd;
	
    end IncidentEntitiesIterator;    


    class IncidentRelationsIterator  from GraphDS
    
    uses MapOfTransient from TColStd,
         MapIteratorOfMapOfTransient from TColStd
    
    raises NoMoreObject from Standard,
           NoSuchObject from Standard
    is
    	Create 
        returns IncidentRelationsIterator from GraphDS;
	
	Create (G : RelationGraph from GraphDS; 
    	        R : Relation      from GraphDS) 
        returns IncidentRelationsIterator from GraphDS;
	
    	Initialize (me : in out; G : RelationGraph from GraphDS; 
                                 R : Relation      from GraphDS); 
            ---Level: Public
	
    	More (me)  
    	---Level: Public 
    	returns Boolean from Standard;
	
    	Next (me : in out) 
    	---Level: Public 
    	raises NoMoreObject from Standard;
	
    	Value (me) 
    	---C++: return const&
    	---Level: Public 
    	returns Relation from GraphDS
    	raises NoSuchObject from Standard;
	
    fields

        myMap       : MapOfTransient from TColStd;
    	myRelations : MapIteratorOfMapOfTransient from TColStd;    
	
    end IncidentRelationsIterator;

is

    Create 
    returns RelationGraph from GraphDS;
    	---Purpose: Creates an empty relation graph.

    Create (other : RelationGraph from GraphDS)
    returns RelationGraph from GraphDS;

    IsEmpty (me) 
    	---Purpose: tests if <me> contains any Entity.
        ---Level: Public
    returns Boolean from Standard;
    
    Clear (me : in out);
	---Purpose: Removes all the  Entities and all  the relations of
	--          <me>.
        ---Level: Public
    
    Contains (me; E : Entity from GraphDS) 
    	---Purpose: tests if <me> contains <E>.
        ---Level: Public    
    returns Boolean from Standard;
    
    Contains (me; R : Relation from GraphDS) 
	---Purpose: tests if <me> contains <rel>.
        ---Level: Public    
    returns Boolean from Standard;

    NbEntities (me) 
    	---Purpose: returns the number of Entity of me.
        ---Level: Public
    returns Integer from Standard;
    
    NbRelations (me) 
	---Purpose: returns the number of Relations of <me>.
        ---Level: Public
    returns Integer from Standard;

    IsInRelation (me; E : Entity from GraphDS) 
	---Purpose: To  Know if <E> is  in relation (as input,output
	--          or both as well) with others Entities of <me>.
        ---Level: Public    
    returns Boolean from Standard
    raises NoSuchObject from Standard;

    IsInput (me; E : Entity from GraphDS) 
    returns Boolean from Standard
	---Purpose: returns True if <E>
        ---Level: Public
    raises NoSuchObject from Standard;

    IsOutput (me; E : Entity from GraphDS) 
    returns Boolean from Standard
    	---Purpose: returns True if <E> is  at least output  of one of
    	--          its relation.
        ---Level: Public
    raises NoSuchObject from Standard;

    IsDependent (me; E : Entity from GraphDS) 
    returns Boolean from Standard
	---Purpose: returns True if <E> is  not input of  one of its
	--          relation.
        ---Level: Public
    raises NoSuchObject from Standard;

    AddEntity (me : in out; value : GraphDS_Item)	
    ---Purpose: Creates an adds a new Entity (which contains item)
    --          to <me>.
    ---Level: Public
    returns Entity from GraphDS;
    
    RemoveEntity (me : in out; E : Entity from GraphDS)
    	---Purpose: Removes a Entity <E> of <me>.  Be carefull than an
    	--          exception is raised if <E> is  still member of any
    	--          relation of <me>.
        ---Level: Public
    raises NoSuchObject from Standard,
           DomainError  from Standard;

    AddRelation (me : in out; value : GraphDS_Attribute)
    	---Purpose: Creates  an adds a  new  Relation  (which contains
    	--          attribute)   to <me>. 
        ---Level: Public
    returns Relation from GraphDS;

    RemoveRelation (me : in out; R : Relation from GraphDS)
    	---Purpose: Removes a relation  <R> of <me>. 
        ---Level: Public
    raises NoSuchObject from Standard;

    ---Purpose: relation editing function

    IsEmpty (me; R : Relation)
	---Purpose: returns TRUE if noone entity is member of <R>.
        ---Level: Public
    returns Boolean from Standard
    raises NoSuchObject from Standard;    
    
    Add (me : in out; R : Relation; E : Entity)
    	---Purpose: add an InputAndOutput entity <E> to <R>
        ---Level: Public
    raises NoSuchObject from Standard;
 
    AddInput  (me : in out; R : Relation; E : Entity)
    	---Purpose: add OnlyInput entity <E> to <R>.
        ---Level: Public
    raises NoSuchObject from Standard;

    AddOutput (me : in out; R : Relation; E : Entity)
    	---Purpose: add an OnlyOutput entity <E> to <R>.
        ---Level: Public
    raises NoSuchObject from Standard;
    
    Add (me : in out; R    : Relation; 
                      E    : Entity;
		      role : EntityRole from GraphDS)
    	---Purpose: add an entity <E> to <R> with role <role>.
        ---Level: Public
    raises NoSuchObject from Standard;
    
    SetRole (me : in out; R    : Relation; 
                          E    : Entity;
		          role : EntityRole from GraphDS)
    	---Purpose: set a new role <role> for the entity <E> member of <R>.
        ---Level: Public
    raises NoSuchObject from Standard;
    
    Remove (me : in out; R : Relation; E : Entity)
    	---Purpose: remove the entity <E> member of <R>.
        ---Level: Public
    raises NoSuchObject from Standard;

fields

    myEntities   : MapOfTransient from TColStd;
    myRelations  : MapOfTransient from TColStd;
    
friends

    class EntitiesIterator from GraphDS,
    class RelationsIterator from GraphDS

end RelationGraph;








