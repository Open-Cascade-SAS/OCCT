-- File:	ShapeProcess_UOperator.cdl
-- Created:	Tue Aug 22 12:06:13 2000
-- Author:	Andrey BETENEV
--		<abv@nnov.matra-dtv.fr>
---Copyright:	 Matra Datavision 2000


class UOperator from ShapeProcess inherits Operator from ShapeProcess

    ---Purpose: Defines operator as container for static function
    --          OperFunc. This allows user to create new operators 
    --          without creation of new classes

uses

    OperFunc from ShapeProcess,
    Context from ShapeProcess

is

    Create (func: OperFunc from ShapeProcess);
    	---Purpose: Creates operator with implementation defined as
	--          OperFunc (static function)

    Perform (me: mutable; context: Context from ShapeProcess) 
    returns Boolean is redefined;
    	---Purpose: Performs operation and records changes in the context

fields

    myFunc: OperFunc from ShapeProcess;

end UOperator;
