-- Created on: 1996-02-13
-- Created by: Yves FRICAUD
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Modified by skv - Tue Mar 15 16:17:37 2005
-- Add methods for supporting history.

class MakeOffsetShape from BRepOffsetAPI inherits MakeShape from BRepBuilderAPI

	---Purpose: Describes functions to build a shell out of a shape. The
    	-- result is an unlooped shape parallel to the source shape.
    	-- A MakeOffsetShape object provides a framework for:
    	-- - defining the construction of a shell
    	-- - implementing the construction algorithm
    	-- - consulting the result.

uses
    MakeOffset  from BRepOffset,
    Mode        from BRepOffset,
    Shape       from TopoDS,
    Face        from TopoDS,
    Edge        from TopoDS,
    Vertex      from TopoDS, 
    ListOfShape from TopTools,		    	    
    JoinType    from GeomAbs
    
is

    Create returns MakeOffsetShape from BRepOffsetAPI;
    
    Create ( S            : Shape    from TopoDS;
             Offset       : Real     from Standard;
	     Tol          : Real     from Standard;
	     Mode         : Mode     from BRepOffset = BRepOffset_Skin;
    	     Intersection : Boolean  from Standard   = Standard_False;
	     SelfInter    : Boolean  from Standard   = Standard_False;
             Join         : JoinType from GeomAbs    = GeomAbs_Arc)
    	---Purpose: Constructs a shape parallel to the shape S, where
    	-- - S may be a face, a shell, a solid or a compound of these shape kinds;
    	-- - Offset is the offset value. The offset shape is constructed:
    	-- - outside S, if Offset is positive,
    	-- - inside S, if Offset is negative;
    	-- - Tol defines the coincidence tolerance criterion for generated shapes;
    	-- - Mode defines the construction type of parallels
    	--   applied to the free edges of shape S; currently, only one
    	--   construction type is implemented, namely the one where the free
    	-- edges do not generate parallels; this corresponds to the default
    	--   value BRepOffset_Skin;
    	-- - Intersection specifies how the algorithm must work in
    	--   order to limit the parallels to two adjacent shapes:
    	-- - if Intersection is false (default value), the intersection
    	-- is calculated with the parallels to the two adjacent shapes,
    	-- - if Intersection is true, the intersection is calculated by
    	-- taking all generated parallels into account; this computation method is
    	-- more general as it avoids some self-intersections generated in the
    	-- offset shape from features of small dimensions on shape S, however this
    	-- method has not been completely implemented and therefore is not
    	-- recommended for use;
    	-- - SelfInter tells the algorithm whether a computation
    	--   to eliminate self-intersections must be applied to the resulting
    	-- shape; however, as this functionality is not yet
    	-- implemented, it is recommended to use the default value (false);
    	-- - Join defines how to fill the holes that may appear between
    	--   parallels to the two adjacent faces. It may take values
    	--   GeomAbs_Arc or GeomAbs_Intersection:
    	-- - if Join is equal to GeomAbs_Arc, then pipes are generated
    	-- between two free edges of two adjacent parallels,
    	-- and spheres are generated on "images" of vertices;
    	--           it is the default value,
    	-- - if Join is equal to GeomAbs_Intersection, then the parallels to the
    	-- two adjacent faces are enlarged and intersected,
    	-- so that there are no free edges on parallels to faces.
    	--   Warnings
    	-- 1. All the faces of the shape S should be based on the surfaces
    	-- with continuity at least C1.
    	-- 2. The offset value should be sufficiently small to avoid
    	-- self-intersections in resulting shape. Otherwise these
    	-- self-intersections may appear inside an offset face if its
    	-- initial surface is not plane or sphere or cylinder, also some
    	-- non-adjacent offset faces may intersect each other. Also, some
    	-- offset surfaces may "turn inside out".
    	--   3. The algorithm may fail if the shape S contains vertices where
    	-- more than 3 edges converge.
    	-- 4. Since 3d-offset algorithm involves intersection of surfaces,
    	-- it is under limitations of surface intersection algorithm.
    	-- 5. A result cannot be generated if the underlying geometry of S is
    	-- BSpline with continuity C0. 
    	-- Exceptions
    	-- Geom_UndefinedDerivative if the underlying
    	-- geometry of S is BSpline with continuity C0.
    returns MakeOffsetShape from BRepOffsetAPI;
    
    MakeOffset (me) returns MakeOffset from BRepOffset
    	---C++: return const &
	---Level: Advanced
    is virtual;
    
    Build (me : in out)
	---Purpose: Builds the resulting shape (redefined from MakeShape).
	---Level: Public     
    is redefined;
    
    
    Generated (me: in out; S : Shape from TopoDS)
    	---Purpose: Returns the  list   of shapes generated   from the
    	--          shape <S>. 
        ---C++: return const & 
        ---Level: Public
    returns ListOfShape from TopTools
    is redefined virtual;


-- Modified by skv - Tue Mar 15 16:17:37 2005 Begin
-- Add methods for supporting history.

    GeneratedEdge  (me: in out; S : Shape from TopoDS)
    	---Purpose: Returns the list of edges generated from the shape <S>. 
        ---C++: return const & 
        ---Level: Public
    returns ListOfShape from TopTools;


-- Query offset join type.

    GetJoinType(me) 
    	---Purpose: Returns offset join type.
    returns JoinType from GeomAbs 
    is static;
 
 
-- Modified by skv - Tue Mar 15 16:17:37 2005 End

fields

    myOffsetShape     : MakeOffset  from BRepOffset is protected;

end MakeOffsetShape;
