-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class CompositeCurveSegment from StepGeom 

inherits TShared from MMgt

uses

	TransitionCode from StepGeom, 
	Boolean from Standard, 
	Curve from StepGeom
is

	Create returns mutable CompositeCurveSegment;
	---Purpose: Returns a CompositeCurveSegment

	Init (me : mutable;
	      aTransition : TransitionCode from StepGeom;
	      aSameSense : Boolean from Standard;
	      aParentCurve : mutable Curve from StepGeom) is virtual;

	-- Specific Methods for Field Data Access --

	SetTransition(me : mutable; aTransition : TransitionCode);
	Transition (me) returns TransitionCode;
	SetSameSense(me : mutable; aSameSense : Boolean);
	SameSense (me) returns Boolean;
	SetParentCurve(me : mutable; aParentCurve : mutable Curve);
	ParentCurve (me) returns mutable Curve;

fields

	transition : TransitionCode from StepGeom; -- an Enumeration
	sameSense : Boolean from Standard;
	parentCurve : Curve from StepGeom;

end CompositeCurveSegment;
