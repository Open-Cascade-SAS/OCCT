-- Created on: 1991-01-14
-- Created by: Arnaud BOUZY
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


deferred class SingleRelation from Expr

inherits GeneralRelation from Expr

uses GeneralExpression from Expr,
    NamedUnknown from Expr,
    AsciiString from TCollection

raises OutOfRange

is

    SetFirstMember(me :mutable; exp : GeneralExpression)
    ---Purpose: Defines the first member of the relation
    ---Level : Internal
    is static;
    
    SetSecondMember(me :mutable; exp : GeneralExpression)
    ---Purpose: Defines the second member of the relation
    ---Level : Internal
    is static;
    
    FirstMember(me)
    ---Purpose: Returns the first member of the relation
    ---Level : Internal
    returns GeneralExpression
    is static;

    SecondMember(me)
    ---Purpose: Returns the second member of the relation
    ---Level : Internal
    returns GeneralExpression
    is static;

    IsLinear(me)
    ---Purpose: Tests if <me> is linear between its NamedUnknowns.
    returns Boolean
    is static;

    NbOfSubRelations(me)
    ---Purpose: Returns the number of relations contained in <me>.
    returns Integer
    is static;
    
    NbOfSingleRelations(me)
    ---Purpose: Returns the number of SingleRelations contained in 
    --          <me> (Always 1).
    returns Integer
    is static;

    SubRelation(me; index : Integer)
    ---Purpose: Returns the relation denoted by <index> in <me>.
    --          An exception is raised if index is out of range.
    returns any GeneralRelation
    raises OutOfRange
    is static;

    Contains(me; exp : GeneralExpression)
    ---Purpose: Tests if <me> contains <exp>.
    returns Boolean;
    
    Replace(me : mutable ; var : NamedUnknown ; with : GeneralExpression);
    ---Purpose: Replaces all occurences of <var> with <with> in <me>.
    
fields

    myFirstMember : GeneralExpression;
    mySecondMember : GeneralExpression;

end SingleRelation;
