-- Created on: 1991-08-02
-- Created by: Laurent BUCHARD
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

generic class PolygonTool from IntCurveSurface(
                  ThePoint       as any;
                  ThePolygon     as any;
                  TheBoundingBox as any)

	---Purpose: 

raises  OutOfRange from Standard


is  


    Bounding       (myclass; thePolygon : ThePolygon)
    	    	    returns TheBoundingBox;
    ---Purpose: Give the bounding box of the polygon.
    ---C++: inline 
    ---C++: return const &

    DeflectionOverEstimation
    	    	   (myclass; thePolygon : ThePolygon)
    		   ---C++: inline
		   returns Real from Standard;

    Closed         (myclass; thePolygon : ThePolygon)
    	            ---C++: inline
    	    	    returns Boolean from Standard;

    NbSegments     (myclass; thePolygon : ThePolygon)
                    ---C++: inline
		   returns Integer from Standard;

    BeginOfSeg     (myclass; thePolygon : ThePolygon;
    	    	    Index : in Integer)
		    ---C++: inline
    	    	    returns ThePoint
    	    	    raises OutOfRange from Standard;
                    ---C++: return const &
    ---Purpose: Give the point of range Index in the Polygon. 

    EndOfSeg       (myclass; thePolygon : ThePolygon;
    	    	    Index : in Integer)
		    ---C++: inline
    	    	    returns ThePoint
    	    	    raises OutOfRange from Standard;
		    ---C++: return const &
    ---Purpose: Give the point of range Index in the Polygon. 


    Dump           (myclass; thePolygon : ThePolygon);
		 
end PolygonTool;








