-- Created on: 1994-04-18
-- Created by: Modelistation
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.





class Text2D from Draw inherits Drawable2D from Draw

	---Purpose: 

uses Pnt2d from gp,
    Color from Draw,
    Display from Draw,
    AsciiString from TCollection

is

    Create(p : Pnt2d; T : CString; col : Color)
    returns mutable Text2D from Draw;
    
    Create(p : Pnt2d; T : CString; col : Color;
    	   moveX : Integer; moveY : Integer)
    returns mutable Text2D from Draw;
    
    SetPnt2d(me : mutable; p : Pnt2d);

    DrawOn(me; dis : in out Display);

fields

    myPoint : Pnt2d        from gp;
    myColor : Color        from Draw;
    myText  : AsciiString  from TCollection;
    mymoveX : Integer      from Standard;
    mymoveY : Integer      from Standard;
    
end Text2D;
