-- Created on: 1992-08-27
-- Created by: Christophe MARION
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DrawableEdgeTool from HLRTest inherits Drawable3D from Draw

	---Purpose: 

uses
    Boolean  from Standard,
    Integer  from Standard,
    Display  from Draw,
    Algo     from HLRBRep,
    Data     from HLRBRep,
    EdgeData from HLRBRep

is
    Create(Alg     : Algo    from HLRBRep;
           Visible : Boolean from Standard;
           IsoLine : Boolean from Standard;
           Rg1Line : Boolean from Standard;
           RgNLine : Boolean from Standard;
           ViewId  : Integer from Standard)
    returns DrawableEdgeTool from HLRTest;
    
    DrawOn(me; D : in out Display from Draw);
    
    InternalDraw(me; D   :in out Display from Draw;
                     typ :       Integer from Standard)
    is static private;
    
    DrawFace(me; D      : in out Display from Draw;
                 typ    :        Integer from Standard;
                 nCB    :        Integer from Standard;
                 iface  :        Integer from Standard;
		 e2,iCB : in out Integer from Standard;
                 DS     : in out Data    from HLRBRep)
    is static private;
    
    DrawEdge(me; D      : in out Display  from Draw;
                 inFace :        Boolean  from Standard;
                 typ    :        Integer  from Standard;
                 nCB    :        Integer  from Standard;
                 ie     :        Integer  from Standard;
		 e2,iCB : in out Integer  from Standard;
                 ed     : in out EdgeData from HLRBRep)
    is static private;
    
fields
    myAlgo    : Algo    from HLRBRep;
    myVisible : Boolean from Standard;
    myIsoLine : Boolean from Standard;
    myRg1Line : Boolean from Standard;
    myRgNLine : Boolean from Standard;
    myViewId  : Integer from Standard;

end DrawableEdgeTool;
