-- Created on: 1992-10-22
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

generic class PathPoint from IntStart
    (TheVertex as any;
     TheArc    as any)

	---Purpose: This class describes a point on an arc which
	--          solution intersection between 2 surfaces.

uses Pnt          from gp,
     Vec          from gp,
     Dir2d        from gp

raises DomainError from Standard

is

    Create
    
	returns PathPoint from IntStart;


    Create(P: Pnt from gp; Tol: Real from Standard;
           V: TheVertex; A: TheArc; Parameter: Real from Standard)

    	returns PathPoint from IntStart;
	

    Create(P: Pnt from gp; Tol: Real from Standard;
           A: TheArc; Parameter: Real from Standard)
	
	returns PathPoint from IntStart;


    SetValue(me: in out; P: Pnt from gp; Tol: Real from Standard;
                         V: TheVertex; A: TheArc;
                         Parameter: Real from Standard)

	---C++: inline
    
    	is static;


    SetValue(me: in out; P: Pnt from gp; Tol: Real from Standard;
                         A: TheArc; Parameter: Real from Standard)
	
	---C++: inline
    
	is static;


    Value(me)
    
    	returns Pnt from gp
	---C++: return const&
	---C++: inline
    
	is static;


    Tolerance(me)
    
    	returns Real from Standard
	---C++: inline
    
	is static;


    IsNew(me)
    
    	returns Boolean from Standard
	---C++: inline
    
	is static;
    

    Vertex(me)
    
    	returns any TheVertex
	---C++: return const&
	---C++: inline
    
	raises DomainError from Standard
	is static;


    Arc(me)
    
    	returns any TheArc
	---C++: return const&
	---C++: inline
    
	is static;


    Parameter(me)
    
    	returns Real        from Standard
	---C++: inline
    
	raises  DomainError from Standard
	is static;

fields

    point : Pnt          from gp;
    tol   : Real         from Standard;
    isnew : Boolean      from Standard;
    vtx   : TheVertex;
    arc   : TheArc;
    param : Real         from Standard;

end PathPoint;
