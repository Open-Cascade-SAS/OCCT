-- Created on: 1998-03-12
-- Created by: Pierre BARRAS
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SplitCurve2d from ShapeUpgrade inherits SplitCurve from ShapeUpgrade

    	---Purpose: Splits a 2d curve with a criterion.
    
uses     
    Curve          from Geom2d,
    HArray1OfCurve from TColGeom2d
   
is 
 
    Create returns SplitCurve2d from ShapeUpgrade;
    	---Purpose: Empty constructor.

    Init (me: mutable; C: Curve from  Geom2d);
       	---Purpose: Initializes with pcurve with its first and last parameters.
	
    Init (me: mutable; C          : Curve from  Geom2d;
    	    	       First, Last: Real);
       	---Purpose: Initializes with pcurve with its parameters.
	
    Build (me: mutable; Segment: Boolean) is redefined;
       ---Purpose: If Segment is True, the result is composed with
       --  segments of the curve bounded by the SplitValues.  If
       --  Segment is False, the result is composed with trimmed
       --  Curves all based on the same complete curve.
       --  
    GetCurves(me) returns HArray1OfCurve from TColGeom2d;
       ---C++: return const &
       
fields 
 
    myCurve          : Curve from Geom2d is protected;
    myResultingCurves: HArray1OfCurve from TColGeom2d is protected;
    
end;
    
