-- Created on: 1992-08-18
-- Created by: Modelistation
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




private class Line from Hatch

	---Purpose: Stores a Line in the Hatcher. Represented by :
	--          
	--          * A Lin2d from gp, the geometry of the line.
	--          
	--          * Bounding parameters for the line.
	--          
	--          * A sorted List  of Parameters, the  intersections
	--          on the line.

uses
    Real                from Standard,
    Integer             from Standard,
    Boolean             from Standard,
    Lin2d               from gp,
    LineForm            from Hatch,
    SequenceOfParameter from Hatch

is

    Create;
    
    Create(L : Lin2d from gp; T : LineForm from Hatch)
    returns Line from Hatch;
    
    AddIntersection(me       : in out; 
                    Par1     : Real    from Standard;
		    Start    : Boolean from Standard;
                    Index    : Integer from Standard;
                    Par2     : Real    from Standard;
    	    	    theToler : Real    from Standard)
	---Purpose: Insert a new intersection in the sorted list.
    is static;
    
fields

    myLin    : Lin2d               from gp;
    myForm   : LineForm            from Hatch;
    myInters : SequenceOfParameter from Hatch;

friends
    class Hatcher from Hatch

end Line;
