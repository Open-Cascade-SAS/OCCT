-- Created on: 1998-03-26
-- Created by: # Andre LIEUTIER
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class GlobalTranslationConstraint from Plate
---Purpose: force a set of UV points to translate without deformation
--          
--          
uses 
 XY from gp, 
 SequenceOfXY from  TColgp,
 LinearXYZConstraint from Plate

is
    Create(SOfXY  :  SequenceOfXY) returns GlobalTranslationConstraint;
    --  SofXY is  a set of UV parametres  for which The Plate function
    --  will give the same value 
    --  
    --  The Sequence length have to be at least 2.

      
    --      
    -- Accessors :
    LXYZC(me) returns LinearXYZConstraint;
    ---C++: inline 
    ---C++: return const &


fields
    myLXYZC : LinearXYZConstraint;
    
end;


