-- File:        ShellBasedSurfaceModel.cdl
-- Created:     Mon Dec  4 12:02:31 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWShellBasedSurfaceModel from RWStepShape

	---Purpose : Read & Write Module for ShellBasedSurfaceModel

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     ShellBasedSurfaceModel from StepShape,
     EntityIterator from Interface

is

	Create returns RWShellBasedSurfaceModel;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable ShellBasedSurfaceModel from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : ShellBasedSurfaceModel from StepShape);

	Share(me; ent : ShellBasedSurfaceModel from StepShape; iter : in out EntityIterator);

end RWShellBasedSurfaceModel;
