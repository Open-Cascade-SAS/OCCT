-- Created on: 1997-11-03
-- Created by: Jean-Louis Frenkel
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class StorageDriver from PCDM inherits Writer from PCDM

    ---Purpose: persistent implemention of storage.
    --
    --          The  application  must redefine one the two Make()
    --           methods.  The first one, if  the application wants to
    --          put only one document in the storage file.
    --          
    --            The  second  method  should  be   redefined  to  put
    --            additional document  that   could  be  used by   the
    --          retrieval instead of the principal document, depending
    --          on the schema used during the retrieval.  For example,
    --          a    second     document   could   be     a   standard
    --             CDMShape_Document.    This  means   that a   client
    --          application will already be able to extract a CDMShape_Document
    --          of the file, if the Shape Schema remains unchanged.
    --          
    ---Category: persistent implemention of storage.

uses
    Document from CDM,
    Document from PCDM,
    Data from Storage,
    ExtendedString from TCollection,
    Schema from Storage,
    SequenceOfExtendedString from TColStd,
    SequenceOfDocument from PCDM,
    StoreStatus from PCDM

raises NoSuchObject from Standard,DriverError from PCDM
is


    Make(me: mutable; aDocument: Document from CDM)
    returns Document from PCDM 
    is virtual;
    ---Purpose: raises NotImplemented.

    Make(me: mutable; aDocument: Document from CDM; Documents: out SequenceOfDocument from PCDM)
    is virtual;
    ---Purpose:By default, puts  in the Sequence the  document returns
    --            by the previous Make method.
    --            

    --          
    SchemaName(me) returns ExtendedString from TCollection
    is deferred;
    
    LoadExtensions(me: mutable; aSchema: Schema from Storage; Extensions: SequenceOfExtendedString from TColStd)
    is virtual;
    
    Write(me: mutable; aDocument: Document from CDM; aFileName: ExtendedString from TCollection)
    raises DriverError
    ---Purpose:  Warning! raises DriverError if an error occurs during inside the
    --          Make method.
    is redefined virtual;
    ---Purpose: stores the content of the Document into a new file.
    --          
    --          by  default  Write will  use Make   method to build a persistent
    --          document and the Schema method to write the persistent document.
    --          

    SetFormat (me : mutable; aformat : ExtendedString from TCollection);

    GetFormat (me)
    returns ExtendedString from TCollection;
    
    IsError   (me) returns Boolean from Standard;
    SetIsError(me : mutable; theIsError : Boolean);
    
    GetStoreStatus   (me) returns StoreStatus from PCDM;
    SetStoreStatus(me : mutable; theStoreStatus : StoreStatus from PCDM);
 
fields 

    myFormat : ExtendedString from TCollection;
    myIsError: Boolean        from Standard;
    myStoreStatus: StoreStatus from PCDM;

end StorageDriver from PCDM;
