-- Created on: 1995-01-13
-- Created by: GG
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MarkMap from Aspect inherits TShared from MMgt

	---Version: 0.0

	---Purpose: This class defines a MarkMap object.
	---Keywords:
	---Warning:
	---References:
uses
	MarkerStyle		from Aspect,
	MarkMapEntry 		from Aspect,
	SequenceOfMarkMapEntry 	from Aspect

raises
	BadAccess 	from Aspect

is
	Create returns MarkMap from Aspect;

        AddEntry (me : mutable; AnEntry : MarkMapEntry from Aspect)
	---Level: Public
        ---Purpose: Adds an entry in the mark map <me>.
        --  Warning: Raises BadAccess if MarkMap size is exceeded.
        raises BadAccess from Aspect;

        AddEntry (me : mutable; aStyle : MarkerStyle from Aspect)
                                        returns Integer from Standard;
        ---Level: Public
        ---Purpose: Search an identical marker style entry in the mark map <me>
        -- and returns the MarkMapEntry Index if exist.
        -- Or add a new entry and returns the computed MarkMapEntry index used.
 
        Size( me ) returns Integer from Standard is static;
        ---Level: Public
        ---Purpose: Returns the Allocated markmap Size
 
        Index( me ; aMarkmapIndex : Integer ) returns Integer from Standard
        ---Level: Public
        ---Purpose: Returns the MarkMapEntry.Index of the MarkMap
        --          at rank <aMarkmapIndex> .
        raises BadAccess from Aspect is static;
        ---Trigger: Raises BadAccess if the index less than 1 or
        --          greater than Size.
 
	Dump( me ) ;

	Entry ( me ;
		AnIndex : Integer from Standard )
	returns MarkMapEntry from Aspect
	---Level: Public
	---Purpose: Returns the Mark map entry with the index <AnIndex>.
	--  Warning: Raises BadAccess if the index less than 1 or
	--	    greater than Size.
	raises BadAccess from Aspect is static;

fields

	mydata	    : 	SequenceOfMarkMapEntry from Aspect is protected;

end MarkMap ;
