-- File:        CompositeCurve.cdl
-- Created:     Mon Dec  4 12:02:24 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWCompositeCurve from RWStepGeom

	---Purpose : Read & Write Module for CompositeCurve

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     CompositeCurve from StepGeom,
     EntityIterator from Interface

is

	Create returns RWCompositeCurve;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable CompositeCurve from StepGeom);

	WriteStep (me; SW : in out StepWriter; ent : CompositeCurve from StepGeom);

	Share(me; ent : CompositeCurve from StepGeom; iter : in out EntityIterator);

end RWCompositeCurve;
