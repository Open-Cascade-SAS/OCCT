-- Created on: 2000-08-21
-- Created by: Andrey BETENEV
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



package ShapeProcess 

    	---Purpose: Shape Processing module
	-- allows to define and apply general Shape Processing as a
	-- customizable sequence of Shape Healing operators. The
	-- customization is implemented via user-editable resource
	-- file which defines sequence of operators to be executed
	-- and their parameters.

uses

    Dico,
    Resource,
    TCollection,
    TColStd,
    GeomAbs,
    TopAbs,
    TopoDS,
    TopTools,
    BRepTools,
    Message,
    ShapeExtend,
    ShapeBuild

is

    class Context; 
    	---Purpose: Provides general context for processing (resource file)
    	class ShapeContext;
	    ---Purpose: Extends context to support processing of the shape

    deferred class Operator;
    	---Purpose: Defines interface to Operator which do the job
	primitive OperFunc;
	class UOperator;
	    ---Purpose: Customizable operator-container loaded by OperFunc

    class OperLibrary;
    	---Purpose: Provides standard set of operators

    class DictionaryOfOperator instantiates 
    	  Dictionary from Dico (Operator from ShapeProcess);

    RegisterOperator (name: CString; op: Operator from ShapeProcess)
    returns Boolean;
    	---Purpose: Registers operator to make it visible for Performer

    FindOperator (name: CString; op: out Operator from ShapeProcess)
    returns Boolean;
    	---Purpose: Finds operator by its name

    Perform (context: Context from ShapeProcess; seq: CString) 
    returns Boolean;
    	---Purpose: Performs a specified sequence of operators on Context
	--          Resource file and other data should be already loaded
	--          to Context (including description of sequence seq)

end ShapeProcess;
