-- Created on: 2000-05-10
-- Created by: Andrey BETENEV
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1

class RoleSelect from StepBasic
inherits SelectType from StepData

    ---Purpose: Representation of STEP SELECT type RoleSelect

uses
    ActionAssignment from StepBasic,
    ActionRequestAssignment from StepBasic,
    ApprovalAssignment from StepBasic,
    ApprovalDateTime from StepBasic,
    CertificationAssignment from StepBasic,
    ContractAssignment from StepBasic,
    DocumentReference from StepBasic,
    EffectivityAssignment from StepBasic,
    GroupAssignment from StepBasic,
    NameAssignment from StepBasic,
    SecurityClassificationAssignment from StepBasic

is
    Create returns RoleSelect from StepBasic;
	---Purpose: Empty constructor

    CaseNum (me; ent: Transient) returns Integer;
	---Purpose: Recognizes a kind of RoleSelect select type
	--          1 -> ActionAssignment from StepBasic
	--          2 -> ActionRequestAssignment from StepBasic
	--          3 -> ApprovalAssignment from StepBasic
	--          4 -> ApprovalDateTime from StepBasic
	--          5 -> CertificationAssignment from StepBasic
	--          6 -> ContractAssignment from StepBasic
	--          7 -> DocumentReference from StepBasic
	--          8 -> EffectivityAssignment from StepBasic
	--          9 -> GroupAssignment from StepBasic
	--          10 -> NameAssignment from StepBasic
	--          11 -> SecurityClassificationAssignment from StepBasic
	--          0 else

    ActionAssignment (me) returns ActionAssignment from StepBasic;
	---Purpose: Returns Value as ActionAssignment (or Null if another type)

    ActionRequestAssignment (me) returns ActionRequestAssignment from StepBasic;
	---Purpose: Returns Value as ActionRequestAssignment (or Null if another type)

    ApprovalAssignment (me) returns ApprovalAssignment from StepBasic;
	---Purpose: Returns Value as ApprovalAssignment (or Null if another type)

    ApprovalDateTime (me) returns ApprovalDateTime from StepBasic;
	---Purpose: Returns Value as ApprovalDateTime (or Null if another type)

    CertificationAssignment (me) returns CertificationAssignment from StepBasic;
	---Purpose: Returns Value as CertificationAssignment (or Null if another type)

    ContractAssignment (me) returns ContractAssignment from StepBasic;
	---Purpose: Returns Value as ContractAssignment (or Null if another type)

    DocumentReference (me) returns DocumentReference from StepBasic;
	---Purpose: Returns Value as DocumentReference (or Null if another type)

    EffectivityAssignment (me) returns EffectivityAssignment from StepBasic;
	---Purpose: Returns Value as EffectivityAssignment (or Null if another type)

    GroupAssignment (me) returns GroupAssignment from StepBasic;
	---Purpose: Returns Value as GroupAssignment (or Null if another type)

    NameAssignment (me) returns NameAssignment from StepBasic;
	---Purpose: Returns Value as NameAssignment (or Null if another type)

    SecurityClassificationAssignment (me) returns SecurityClassificationAssignment from StepBasic;
	---Purpose: Returns Value as SecurityClassificationAssignment (or Null if another type)

end RoleSelect;
