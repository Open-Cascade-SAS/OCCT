-- Created on: 1993-05-04
-- Created by: Modelistation
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ShapeToHLR from HLRBRep

	---Purpose: compute  the   OutLinedShape  of  a Shape with  an
	--          OutLiner,    a  Projector  and   create  the  Data
	--          Structure of a Shape.

uses
    Shape             from TopoDS,
    Face              from TopoDS,
    IndexedMapOfShape from TopTools,
    OutLiner          from HLRTopoBRep,
    Projector         from HLRAlgo,
    Data              from HLRBRep,
    MapOfShapeTool    from BRepTopAdaptor

is
    Load(myclass; S     :        OutLiner  from HLRTopoBRep;
                  P     :        Projector from HLRAlgo;
		  MST   : in out MapOfShapeTool from BRepTopAdaptor;
                  nbIso :        Integer   from Standard = 0)
    returns Data from HLRBRep;
	---Purpose: Creates  a DataStructure   containing the OutLiner
	--          <S> depending on the projector <P> and nbIso.
		   
    ExploreFace(myclass;
                S      :         OutLiner          from HLRTopoBRep;
                DS     : mutable Data              from HLRBRep;
	        FM     :         IndexedMapOfShape from TopTools;
	        EM     :         IndexedMapOfShape from TopTools;
		i      : in out  Integer           from Standard;
                F      :         Face              from TopoDS;
                closed :         Boolean           from Standard)
    is private;

    ExploreShape(myclass;
                 S    :         OutLiner          from HLRTopoBRep;
                 DS   : mutable Data              from HLRBRep;
		 FM   :         IndexedMapOfShape from TopTools; 
		 EM   :         IndexedMapOfShape from TopTools) 
    is private;

end ShapeToHLR;
