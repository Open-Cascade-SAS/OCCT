-- Created on: 1991-02-06
-- Created by: Arnaud BOUZY
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class RUIterator from Expr

	---Purpose: Iterates on NamedUnknowns in a GeneralRelation. 
    	---Level : Internal

uses GeneralRelation from Expr,
    NamedUnknown from Expr,
    MapOfNamedUnknown from Expr
    
raises NoMoreObject from Standard,
    NoSuchObject from Standard

is

    Create(rel : GeneralRelation)
    ---Purpose: Creates an iterator on every NamedUnknown contained in 
    --          <rel>.
    returns RUIterator;
    
    More(me)
    ---Purpose: Returns False if on other unknown remains.
    returns Boolean
    is static;
    
    Next(me : in out)
    raises NoMoreObject
    is static;
    
    Value(me)
    ---Purpose: Returns current NamedUnknown.
    --          Raises exception if no more unknowns remain.
    returns NamedUnknown
    raises NoSuchObject
    is static;

fields

    myMap : MapOfNamedUnknown;
    myCurrent : Integer;

end RUIterator;
