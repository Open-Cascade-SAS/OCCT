-- Created on: 1993-06-23
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class ShapeData from TopOpeBRepDS

uses 
    
    ListOfInterference from TopOpeBRepDS,
    ListOfShape from TopTools,
    Config from TopOpeBRepDS,
    Orientation from TopAbs
    
is  
    
    Create returns ShapeData;
    Interferences(me) returns ListOfInterference;
    ---C++:return const & 
    ChangeInterferences(me:in out) returns ListOfInterference;
    ---C++:return &
    
    Keep(me) returns Boolean from Standard
    is static;
    ChangeKeep(me : in out; B : Boolean from Standard)
    is static;

fields

    myInterferences : ListOfInterference from TopOpeBRepDS;
    mySameDomain    : ListOfShape from TopTools;
    mySameDomainRef : Integer from Standard;
    mySameDomainOri : Config from TopOpeBRepDS;
    mySameDomainInd : Integer;
    myOrientation : Orientation from TopAbs;
    myOrientationDef : Boolean;
    myAncestorRank : Integer; -- 1 or 2
    myKeep      : Boolean from Standard;

friends 
    
    class DataStructure from TopOpeBRepDS

end ShapeData from TopOpeBRepDS;
