-- Created on: 1993-07-22
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class MakeRevolution from BRepPrimAPI inherits MakeOneAxis from BRepPrimAPI

	---Purpose: Describes functions to build revolved shapes.
    	-- A MakeRevolution object provides a framework for:
    	-- -   defining the construction of a revolved shape,
    	-- -   implementing the construction algorithm, and
    	-- -   consulting the result.

uses
    Ax2        from gp,
    Curve      from Geom,
    OneAxis    from BRepPrim,
    Revolution from BRepPrim

raises
    DomainError from Standard

is
    Create(Meridian  : Curve from Geom)
    returns MakeRevolution from BRepPrimAPI
	---Purpose: Make a revolution body by rotating a curve around Z.
	---Level: Public
    raises
    	DomainError from Standard; -- if M is not in a plane containing Z.

    Create(Meridian  : Curve from Geom; angle : Real)
    returns MakeRevolution from BRepPrimAPI
	---Purpose: Make a revolution body by rotating a curve around Z.
	---Level: Public
    raises
    	DomainError from Standard; -- if M is not in a plane containing Z.

    Create(Meridian  : Curve from Geom; VMin, VMax : Real)
    returns MakeRevolution from BRepPrimAPI
	---Purpose: Make a revolution body by rotating a curve around Z.
	---Level: Public
    raises
    	DomainError from Standard; -- if M is not in a plane containing Z.

    Create(Meridian  : Curve from Geom; VMin, VMax, angle : Real)
    returns MakeRevolution from BRepPrimAPI
	---Purpose: Make a revolution body by rotating a curve around Z.
	---Level: Public
    raises
    	DomainError from Standard; -- if M is not in a plane containing Z.

    Create(Axes : Ax2 from gp; Meridian  : Curve from Geom)
    returns MakeRevolution from BRepPrimAPI
	---Purpose: Make a revolution body by rotating a curve around Z.
	---Level: Public
    raises
    	DomainError from Standard; -- if M is not in a plane containing Z.

    Create(Axes : Ax2 from gp; Meridian  : Curve from Geom; angle : Real)
    returns MakeRevolution from BRepPrimAPI
	---Purpose: Make a revolution body by rotating a curve around Z.
	---Level: Public
    raises
    	DomainError from Standard; -- if M is not in a plane containing Z.

    Create(Axes : Ax2 from gp; Meridian  : Curve from Geom; VMin, VMax : Real)
    returns MakeRevolution from BRepPrimAPI
	---Purpose: Make a revolution body by rotating a curve around Z.
	---Level: Public
    raises
    	DomainError from Standard; -- if M is not in a plane containing Z.

    Create(Axes : Ax2 from gp; Meridian  : Curve from Geom; VMin, VMax, angle : Real)
    returns MakeRevolution from BRepPrimAPI
	---Purpose: Make a revolution body by rotating a curve around Z.
	---Level: Public
    raises
    	DomainError from Standard; -- if M is not in a plane containing Z.
    	---Purpose: For all algorithms the resulting shape is composed of
    	-- -   a lateral revolved face,
    	-- -   two planar faces in planes parallel to the plane z =
    	--   0, and passing by the extremities of the revolved
    	--   portion of Meridian, if these points are not on the Z
    	--   axis (in case of a complete revolved shape, these faces are circles),
    	-- -   and in the case of a portion of a revolved shape, two
    	--   planar faces to close the shape (in the planes u = 0 and u = angle).

    OneAxis(me : in out) returns Address;
	---Purpose: Returns the algorithm.
	---Level: Advanced

    Revolution(me : in out) returns Revolution from BRepPrim
	---Purpose: Returns the algorithm.
	--          
	---C++: return &
	---Level: Public
    is static;

fields 

    myRevolution : Revolution from BRepPrim;

end MakeRevolution;
