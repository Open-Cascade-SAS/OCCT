-- Created on: 1993-01-09
-- Created by: CKY / Contract Toubro-Larsen ( Arun MENON )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Name from IGESBasic  inherits NameEntity

        ---Purpose: defines Name, Type <406> Form <15>
        --          in package IGESBasic
        --          Used to specify a user defined name

uses

        HAsciiString from TCollection

is

        Create returns mutable Name;

        -- Specific Methods pertaining to the class

        Init (me :  mutable; nbPropVal : Integer; aName : HAsciiString);
        ---Purpose : This method is used to set the fields of the class Name
        --       - nbPropVal  : Number of property values, always = 1
        --       - aName      : Stores the Name

        NbPropertyValues (me) returns Integer ;
        ---Purpose : returns the number of property values, which should be 1

        Value (me) returns HAsciiString from TCollection;
        ---Purpose : returns the user defined Name

fields

--
-- Class    : IGESBasic_Name
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class Name.
--
-- Reminder : A Name instance is defined by :
--            - the number of property values (equal to 1)
--            - the name

        theNbPropertyValues : Integer;
        theName             : HAsciiString from TCollection;

end Name;
