-- Created on: 1994-08-31
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




package Draft

uses BRepTools,
     TopoDS,
     TopTools,
     TopLoc,
     TopAbs,

     GeomAbs,
     Geom,
     Geom2d,
     gp,
     
     TColStd,
     StdFail,
     TCollection
     
     
is

    class Modification; --- inherits Modification from BRepTools


    class FaceInfo;
    
    class EdgeInfo;
    
    class VertexInfo;
    
    enumeration ErrorStatus is
    	NoError,
	FaceRecomputation,
	EdgeRecomputation,
	VertexRecomputation
    end ErrorStatus;
    
    
    class DataMapOfFaceFaceInfo instantiates
    	DataMap from TCollection(Face           from TopoDS,
	                         FaceInfo       from Draft,
				 ShapeMapHasher from TopTools);


    class DataMapOfEdgeEdgeInfo instantiates
    	DataMap from TCollection(Edge           from TopoDS,
	                         EdgeInfo       from Draft,
				 ShapeMapHasher from TopTools);


    class DataMapOfVertexVertexInfo instantiates
    	DataMap from TCollection(Vertex         from TopoDS,
	                         VertexInfo     from Draft,
				 ShapeMapHasher from TopTools);




    Angle(F: Face from TopoDS;  Direction: Dir from gp)
    
    	returns Real from Standard
	raises DomainError from Standard;
	
	---Purpose: Returns the draft angle of the  face <F> using the
	--          direction <Direction>.  The  method is valid for :
	--          - Plane  faces,
	--          - Cylindrical or conical faces, when the direction
	--          of the axis of the surface is colinear with the
	--          direction.
	--          Otherwise, the exception DomainError is raised.


end Draft;

