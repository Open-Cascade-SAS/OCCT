-- Created by: Peter KURNEV
-- Copyright (c) 2010-2012 OPEN CASCADE SAS
-- Copyright (c) 2007-2010 CEA/DEN, EDF R&D, OPEN CASCADE
-- Copyright (c) 2003-2007 OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN, CEDRAT,
--                         EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class IteratorSI from BOPDS  
    inherits Iterator from BOPDS

---Purpose:  
    -- The class BOPDS_IteratorSI is  
    --  1.to compute self-intersections between BRep sub-shapes  
    --    of each argument of an operation (see the class BOPDS_DS)
    --    in terms of theirs bounding boxes           
    --  2.provides interface to iterare the pairs of  
    --    intersected sub-shapes of given type 

uses  
    BaseAllocator from BOPCol 

is 
    Create   
    returns IteratorSI from BOPDS;
    ---C++: alias "Standard_EXPORT virtual ~BOPDS_IteratorSI();"   
    ---Purpose:  
    --- Empty contructor  
    ---   
 
    Create (theAllocator: BaseAllocator from BOPCol)  
    returns IteratorSI from BOPDS;
     ---Purpose:  
    ---  Contructor    
    ---  theAllocator - the allocator to manage the memory     
    --- 
    Intersect(me:out) 
    is redefined protected;  
 
end IteratorSI;
