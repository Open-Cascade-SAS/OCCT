-- Created on: 1993-01-29
-- Created by: Isabelle GRIGNON
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class PolyLine from IntPatch

inherits Polygo from IntPatch

uses Pnt2d from gp,
     Box2d from Bnd,
     IType from IntPatch,
     WLine from IntPatch,
     RLine from IntPatch

is

    Create
    returns PolyLine from IntPatch;

    Create (InitDefle: Real from Standard)
   	returns PolyLine from IntPatch;

    SetWLine(me: in out; OnFirst: Boolean from Standard; Line: WLine from IntPatch)
    	is static;

    SetRLine(me: in out; OnFirst: Boolean from Standard; Line: RLine from IntPatch)
      	is static;

    Prepare(me: in out)
      	is static private;

    ResetError(me: in out);

    NbPoints(me) returns Integer;
  
    Point(me; Index : Integer) 
    	returns Pnt2d from gp;
                                      	    	 

fields

    pnt      : Pnt2d   from gp;
    typ      : IType   from IntPatch;
    onfirst  : Boolean from Standard;
    wpoly    : WLine from IntPatch;
    rpoly    : RLine from IntPatch;

end PolyLine;
