-- Created on: 1999-04-15
-- Created by: Denis PASCAL
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class DocumentStorageDriver from MDocStd inherits StorageDriver from PCDM

	---Purpose: storage driver for  a standard document


uses Document           from TDocStd,
     Document           from PDocStd,
     SRelocationTable   from MDF,
     Document           from CDM, 
     MessageDriver      from CDM,       
     Document           from PCDM,
     ExtendedString from  TCollection,
     ASDriverTable from MDF


is


    Create
    returns mutable  DocumentStorageDriver from MDocStd;
    
    CreateDocument (me: mutable) returns Document from PCDM
    ---Purpose: returns an empty PDocStd_Document. may be redefined;
    is virtual;
    	     
    Paste (me : mutable; TDOC   : Document from TDocStd;
                         PDOC   : Document from PDocStd;
			 aReloc : SRelocationTable from MDF);
  

    ---Purpose: virtual  methods of StorageDriver from PCDM
    --          ============================================
    
    Make (me: mutable; aDocument: Document from CDM)
    returns Document from PCDM 
    is redefined;
    
    ---Purpose: virtual methods (may be redefined by specialized application)
    --          =============================================================
    
    SchemaName(me) 
    returns   ExtendedString from  TCollection
    is virtual;
    
    AttributeDrivers(me : mutable; theMessageDriver : MessageDriver from CDM)
    returns ASDriverTable from MDF
    is virtual;
    
fields

    myDrivers : ASDriverTable from MDF;
    
end DocumentStorageDriver;
