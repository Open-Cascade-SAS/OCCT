-- Created by: Peter KURNEV
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


package BOPCol 

	---Purpose:  
    	-- The package contains collection classes 
	-- that are used by  
    	-- partition and  boolean operation algorithms     
uses 
    TCollection
 
is 
    imported BaseAllocator from BOPCol; 
    imported DataMapOfShapeInteger from BOPCol; 
    imported MapOfInteger from BOPCol; 
    imported ListOfInteger from BOPCol; 
    imported PInteger from BOPCol; 
    imported DataMapOfIntegerInteger from BOPCol; 
    imported DataMapOfIntegerListOfInteger from BOPCol; 
    imported IndexedDataMapOfShapeBox from BOPCol; 
    imported IndexedMapOfInteger from BOPCol; 
    imported ListOfShape from BOPCol;   
    imported DataMapOfShapeAddress from BOPCol;   
    imported DataMapOfTransientAddress from BOPCol;   
    imported PListOfInteger from BOPCol;  
    imported VectorOfInteger from BOPCol;  
    imported MapOfShape from BOPCol;  
    imported DataMapOfShapeShape from BOPCol;  
    imported DataMapOfShapeListOfShape from BOPCol;  
    imported MapOfOrientedShape from BOPCol;  
    imported IndexedDataMapOfShapeListOfShape from BOPCol;  
    imported IndexedMapOfShape from BOPCol;  
    imported ListOfListOfShape from BOPCol;  
    imported SequenceOfShape from BOPCol;  
    imported SequenceOfPnt2d from BOPCol;  
    imported DataMapOfIntegerListOfShape from BOPCol;
    imported IndexedDataMapOfIntegerListOfInteger from BOPCol;
    imported IndexedDataMapOfShapeInteger from BOPCol;  
    
end BOPCol;
