-- Created on: 1995-03-15
-- Created by: Robert COUBLANC
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Modified by rob jun 25 98 : Add Method : Reactivate projector...

class ViewerSelector3d from StdSelect inherits ViewerSelector from SelectMgr

    ---Purpose: Selector Usable by Viewers from V3d
    --          Accepts Only Sensitive Entities inheriting Select3D entities...

uses
    View                 from V3d,
    Selection            from SelectMgr,
    EntityOwner          from SelectMgr,
    Projector            from Select3D,
    Group                from Graphic3d,
    Structure            from Graphic3d,
    SequenceOfHClipPlane from Graphic3d,
    Array1OfReal         from TColStd, 
    Array1OfPnt2d        from TColgp,
    SensitivityMode      from StdSelect,
    Lin                  from gp,
    Pnt                  from gp,
    Dir                  from gp,
    XYZ                  from gp

is

    Create  returns ViewerSelector3d from StdSelect;
    ---Purpose: Constructs an empty 3D selector object.

    Create (theProj : Projector from Select3D) returns ViewerSelector3d from StdSelect;
    ---Purpose: Constructs a 3D selector object defined by the projector <theProj>.

    Convert (me : mutable; theSel : Selection from SelectMgr)
    is redefined static;
        ---Level: Public 
        ---Purpose: Processes the projection of the sensitive  primitives
        --          in the active view ; to be done before the selection action...

    Set (me : mutable; theProj : Projector from Select3D) is static;
    ---Purpose: Sets the new projector <theProj> to replace the one used at construction time.

    SetSensitivityMode (me      : mutable;
                        theMode : SensitivityMode from StdSelect) is static;
        ---Purpose: Sets the selection sensitivity mode. SM_WINDOW mode
        -- uses the specified pixel tolerance to compute the sensitivity
        -- value, SM_VIEW mode allows to define the sensitivity manually.

    SensitivityMode (me) returns SensitivityMode from StdSelect;
        ---C++: inline
        ---Purpose: Returns the selection sensitivity mode.

    SetPixelTolerance (me           : mutable;
                       theTolerance : Integer) is static;
    ---Purpose: Sets the pixel tolerance <theTolerance>.

    PixelTolerance (me) returns Integer from Standard;
        ---C++: inline
        ---Purpose: Returns the pixel tolerance.

    Pick (me           : mutable; theXPix, theYPix : Integer;
          theView      : View from V3d) is static;
    ---Level: Public 
    ---Purpose: Picks the sensitive entity at the pixel coordinates of
    -- the mouse <theXPix> and <theYPix>. The selector looks for touched areas and owners.

    Pick (me : mutable; theXPMin, theYPMin, theXPMax, theYPMax : Integer; theView : View from V3d) is static;
    ---Purpose: Picks the sensitive entity according to the minimum
    -- and maximum pixel values <theXPMin>, <theYPMin>, <theXPMax>
    -- and <theYPMax> defining a 2D area for selection in the 3D view aView.

    Pick (me : mutable; thePolyline : Array1OfPnt2d from TColgp; theView : View from V3d) is static;
    ---Level: Public 
    ---Purpose: pick action - input pixel values for polyline selection for selection.

    ---Category: Inquire Methods

    Projector (me) returns Projector from Select3D;
    ---Level: Public 
    ---Purpose: Returns the current Projector.
    ---C++: inline
    ---C++: return const&

    ---Category: Internal Methods
    --           -----------------

    UpdateProj (me      : mutable;
                theView : View from V3d) returns Boolean is static private;
    ---Level: Internal

    DisplayAreas (me      : mutable;
                  theView : View from V3d) is static;
    ---Purpose: Displays sensitive areas found in the view <theView>.

    ClearAreas (me      : mutable;
                theView : View from V3d) is static;
    ---Purpose: Clears the view aView of sensitive areas found in it.

    DisplaySensitive (me : mutable; theView : View from V3d) is static;
    --- Purpose: Displays sensitives in view <theView>.

    ClearSensitive (me : mutable; theView : View from V3d) is static;

    DisplaySensitive (me               : mutable;
                      theSel           : Selection from SelectMgr;
                      theView          : View from V3d;
                      theToClearOthers : Boolean from Standard = Standard_True)
    is static;

    DisplayAreas (me               : mutable;
                  theSel           : Selection from SelectMgr;
                  theView          : View from V3d;
                  theToClearOthers : Boolean from Standard = Standard_True)
    is static;

    ComputeSensitivePrs (me : mutable; theSel: Selection from SelectMgr)
    is static private;
    ---Level: Internal

    ComputeAreasPrs (me : mutable; theSel : Selection from SelectMgr)
    is static private;
    ---Level: Internal

    SetClipping (me : mutable; thePlanes : SequenceOfHClipPlane from Graphic3d) is protected;
    ---Level: Internal
    ---Purpose: Set view clipping for the selector.
    -- @param thePlanes [in] the view planes.

    ComputeClipRange (me; thePlanes : SequenceOfHClipPlane from Graphic3d;
                      thePickLine : Lin from gp;
                      theDepthMin, theDepthMax : out Real from Standard)
      is protected;
    ---Level: Internal
    ---Purpose: Computed depth boundaries for the passed set of clipping planes and picking line.
    -- @param thePlanes [in] the planes.
    -- @param thePickLine [in] the picking line.
    -- @param theDepthMin [out] minimum depth limit.
    -- @param theDepthMax [out] maximum depth limit.

    PickingLine (me; theX, theY : Real from Standard)
      returns Lin from gp
      is redefined protected;
    ---Level: Internal
    ---Purpose: For more details please refer to base class.

    DepthClipping (me; theX, theY : Real from Standard;
                   theMin, theMax : out Real from Standard)
      is redefined protected;
    ---Level: Internal
    ---Purpose: For more details please refer to base class.

    DepthClipping (me; theX, theY : Real from Standard;
                   theOwner : EntityOwner from SelectMgr;
                   theMin, theMax : out Real from Standard)
      is redefined protected;
    ---Level: Internal
    ---Purpose: For more details please refer to base class.

    HasDepthClipping (me; theOwner : EntityOwner from SelectMgr)
      returns Boolean is redefined protected;
    ---Level: Internal
    ---Purpose: For more details please refer to base class.
    
fields

    myProjector         : Projector from Select3D;
    myPrevAt            : Real from Standard[3];
    myPrevUp            : Real from Standard[3];
    myPrevProj          : Real from Standard[3];
    myPrevAxialScale    : Real from Standard[3];
    myPrevFOV           : Real from Standard;
    myPrevScale         : Real from Standard;
    myPrevOrthographic  : Boolean from Standard;
    mySensMode          : SensitivityMode from StdSelect;
    myPixelTolerance    : Integer from Standard;
    myToUpdateTolerance : Boolean from Standard;

    --areas verification...

    myareagroup  : Group                from Graphic3d;
    mysensgroup  : Group                from Graphic3d;
    mystruct     : Structure            from Graphic3d;
    myClipPlanes : SequenceOfHClipPlane from Graphic3d;

end ViewerSelector3d;
