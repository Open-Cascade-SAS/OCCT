-- Created on: 1997-08-01
-- Created by: SMO
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class NamedShapeDriver from TPrsStd inherits Driver from TPrsStd
---Purpose: An implementation of TPrsStd_Driver for named shapes.
uses

  GUID               from Standard,
  Label              from TDF,
  InteractiveObject  from AIS
is

    Create
    returns mutable NamedShapeDriver from TPrsStd;
---Purpose: Constructs an empty named shape driver.
    Update (me : mutable ;
           aLabel      : Label from TDF;
	   anAISObject : in out InteractiveObject from AIS)
    returns Boolean from Standard
    is  redefined virtual;
    --- Purpose: Build the AISObject (if null) or update it.
    --           No compute is done.
    --           Returns <True> if informations was found
    --           and AISObject updated. 
	   

end NamedShapeDriver;

