-- Created on: 1996-04-10
-- Created by: Joelle CHAUVET
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Modified:	Mon Dec  9 10:30:56 1996
--    by:	Joelle CHAUVET
--		G1135 : Empty constructor

class Framework from AdvApp2Var

uses

    Boolean,Real,NoSuchObject from Standard,
    HArray1OfReal from TColStd,
    IsoType from GeomAbs,
    SequenceOfNode,SequenceOfStrip,Iso,Node from AdvApp2Var

raises NoSuchObject from Standard

is

    Create returns Framework;
    Create(Frame : SequenceOfNode; 
           UFrontier, VFrontier : SequenceOfStrip)  
    returns Framework;
    
    FirstNotApprox(me; IndexIso,IndexStrip : out Integer; 
                       anIso : out Iso) 
    ---Purpose: search the Index of the first Iso not approximated,
    --          if all Isos are approximated Standard_False is returned.
    returns Boolean; 

    FirstNode(me; Type : IsoType; IndexIso,IndexStrip : Integer) 
    returns Integer;
    
    LastNode(me; Type : IsoType; IndexIso,IndexStrip : Integer) returns Integer; 
    
    ChangeIso(me: in out; IndexIso,IndexStrip : Integer; anIso : Iso);
    
    Node(me; IndexNode : Integer)
    ---C++: return const&
    ---C++: inline    
    returns Node
    raises NoSuchObject from Standard;
	
    Node(me; U,V : Real) 
    ---C++: return const&
    returns Node
    raises NoSuchObject from Standard;
	
    IsoU(me; U,V0,V1 : Real) 
    ---C++: return const&
    returns Iso
    raises NoSuchObject from Standard;
	
    IsoV(me; U0,U1,V : Real) 
    ---C++: return const&    
    returns Iso
    raises NoSuchObject from Standard;
	
    ChangeNode(me: in out; IndexNode : Integer)
    ---C++: return &
    ---C++: inline    
    returns Node;

    
    UpdateInU(me: in out; CuttingValue : Real);
    
    UpdateInV(me: in out; CuttingValue : Real);
    
    UEquation(me; IndexIso,IndexStrip : Integer) 
    ---C++: return const &
    returns HArray1OfReal; 
    
    VEquation(me; IndexIso,IndexStrip : Integer)
    ---C++: return const & 
     returns HArray1OfReal;
 

fields

    myNodeConstraints    : SequenceOfNode;
    myUConstraints       : SequenceOfStrip;
    myVConstraints       : SequenceOfStrip;

end Framework;

