-- Created on: 1997-04-01
-- Created by: Christian CAILLET
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class FieldListN  from StepData    inherits FieldList  from StepData

    ---Purpose : Describes a list of fields, in a general way
    --           This basic class is for a null size list
    --           Subclasses are for 1, N (fixed) or Dynamic sizes

uses Field from StepData, Array1OfField from StepData

raises OutOfRange

is

    Create (nb : Integer) returns FieldListN;
    ---Purpose : Creates a FieldListN of <nb> Fields

    NbFields (me) returns Integer  is redefined;
    ---Purpose : Returns the count of fields. Here, returns starting <nb>

    Field  (me; num : Integer) returns Field
    ---Purpose : Returns the field n0 <num> between 1 and NbFields (read only)
	raises OutOfRange
    --           Error if <num> out of range
    	is redefined;
    ---C++ : return const &

    CField (me : in out; num : Integer) returns Field
    ---Purpose : Returns the field n0 <num> between 1 and NbFields, in order to
    --           modify its content
	raises OutOfRange
    --           Error if <num> out of range
    	is redefined;
    ---C++ : return &

    Destroy (me: in out) is virtual;
    ---C++ : alias "Standard_EXPORT virtual ~StepData_FieldListN() { Destroy(); }"


fields

    thefields : Array1OfField;

end FieldListN;
