-- Created on: 1997-03-19
-- Created by: Prestataire Mary FABIEN
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Mesure from TestTopOpeTools

uses

    AsciiString from TCollection,
    Array1OfPnt from TColgp,
    HArray1OfPnt from TColgp,
    Pnt from gp

is

    Create returns Mesure from TestTopOpeTools;

    Create(name : AsciiString from TCollection)
    returns Mesure from TestTopOpeTools;

    Create(Pnts : HArray1OfPnt from TColgp)
    returns Mesure from TestTopOpeTools;

    Add(me :in out; n : in Integer from Standard; t : in Real from Standard);

    SetName(me : in out; Name : AsciiString from TCollection);

    Name(me) returns AsciiString from TCollection;
    ---C++: return const&

    Pnts(me) returns Array1OfPnt from TColgp;
    ---C++: return const&

    Pnt(me; I : in Integer) returns Pnt from gp;
    ---C++: return const&

    NPnts(me) returns Integer from Standard;

    Clear(me : in out);

fields

    myName  : AsciiString from TCollection;
    myPnts  : HArray1OfPnt from TColgp;
    myNPnts : Integer from Standard;

end Mesure from TestTopOpeTools;
