-- Created on: 2006-12-05
-- Created by: Sergey  KOCHETKOV
-- Copyright (c) 2006-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class HPackedMapOfInteger from TColStd inherits TShared from MMgt 
 
	  ---Purpose: Extension of TColStd_PackedMapOfInteger class to be manipulated by handle. 
 
uses 
    PackedMapOfInteger from TColStd 
 
is 
    Create( NbBuckets: Integer from Standard = 1 ) returns mutable HPackedMapOfInteger from TColStd;    
     
    Create( theOther:  PackedMapOfInteger from TColStd ) returns mutable HPackedMapOfInteger from TColStd; 
     
    Map( me ) returns PackedMapOfInteger from TColStd 
	---C++: return const &
        ---C++: inline      
    is static;	    	
	  
    ChangeMap( me: mutable ) returns PackedMapOfInteger from TColStd 
    	---C++: return &
        ---C++: inline 
    is static; 	    	
 
fields     
    myMap : PackedMapOfInteger from TColStd; 
 
end HPackedMapOfInteger;     
