-- Created on: 1997-09-03
-- Created by: Christian CAILLET
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class IntVal  from Interface    inherits TShared  from MMgt

    ---Purpose : An Integer through a Handle (i.e. managed as TShared)

uses Integer

is

    Create returns IntVal;

    Value (me) returns Integer;

    CValue (me : mutable) returns Integer;
    ---C++ : return &

fields

    theval : Integer;

end IntVal;
