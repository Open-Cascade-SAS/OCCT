-- Created by: DAUTRY Philippe
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

--      	------------

---Version:	0.0
--Version	Date		Purpose
--		0.0	Mar 13 1997	Creation


class Data from PDF
    inherits Persistent from Standard

	---Purpose: Persistent equivalent of Data from TDF.

uses

    HArray1OfInteger from PColStd,
    HAttributeArray1 from PDF

-- raises

is

    Create
    	returns mutable Data from PDF;

    Create(aVersionNumber : Integer from Standard)
    	returns mutable Data from PDF;

    VersionNumber(me)
    	returns Integer from Standard;
	---Purpose: Returns the value of the field <myVersion>.
	---C++: inline


    Labels(me : mutable;
    	   theLabels : HArray1OfInteger from PColStd);
	---Purpose: Sets the field <myLabels> with <theLabels>.
	---C++: inline

    Labels(me)
    	returns HArray1OfInteger from PColStd;
	---Purpose: Returns the value of the field <myLabels>.
	---C++: inline

    Attributes(me : mutable;
    	   theAttributes : HAttributeArray1 from PDF);
	---Purpose: Sets the field <myAttributes> with <theAttributes>.
	---C++: inline

    Attributes(me)
    	returns HAttributeArray1 from PDF;
	---Purpose: Returns the value of the field <myAttributes>.
	---C++: inline

fields

    myVersion    : Integer          from Standard;
    myLabels     : HArray1OfInteger from PColStd;
    myAttributes : HAttributeArray1 from PDF;

end Data;
