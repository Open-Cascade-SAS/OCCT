-- File:	IGESGraph_ToolHighLight.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolHighLight  from IGESGraph

    ---Purpose : Tool to work on a HighLight. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses HighLight from IGESGraph,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolHighLight;
    ---Purpose : Returns a ToolHighLight, ready to work


    ReadOwnParams (me; ent : mutable HighLight;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : HighLight;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : HighLight;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a HighLight <ent>, from
    --           its specific (own) parameters

    OwnCorrect (me; ent : mutable HighLight) returns Boolean  is static;
    ---Purpose : Sets automatic unambiguous Correction on a HighLight
    --           (NbPropertyValues forced to 1)

    DirChecker (me; ent : HighLight) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : HighLight;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : HighLight; entto : mutable HighLight;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : HighLight;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolHighLight;
