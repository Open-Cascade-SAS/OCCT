-- Created on: 1998-08-20
-- Created by: Philippe MANGIN
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class  Curve3d  from  Approx 

uses
    HCurve         from  Adaptor3d, 
    BSplineCurve   from  Geom, 
    Shape          from  GeomAbs,
    OutOfRange     from  Standard          
    
raises  OutOfRange   from Standard, 
        ConstructionError  from  Standard

is
 
    Create(Curve:  HCurve  from Adaptor3d; 
    	    Tol3d:  Real; 
    	    Order:  Shape  from  GeomAbs; 
    	    MaxSegments:  Integer; 
    	    MaxDegree:  Integer)  returns  Curve3d  from  Approx; 
        ---Purpose: Approximation  of  a  curve  with respect of the  
    --          requiered tolerance Tol3D. 
     
    Curve(me)  returns  BSplineCurve  from  Geom; 
     
    IsDone(me)  returns  Boolean  from  Standard; 
    ---Purpose:  returns  Standard_True  if  the  approximation  has   
    -- been  done  within  requiered tolerance 
     
    HasResult(me) returns Boolean; 
    ---Purpose: returns  Standard_True if the approximation did come out 
    -- with a result that  is not NECESSARELY within the required 
    -- tolerance

    MaxError(me)  returns  Real  from  Standard; 
    ---Purpose:  returns  the  Maximum  Error  (>0 when an approximation 
    --  has  been  done, 0  if  no  approximation) 
     
    Dump(me;  o:  in  out  OStream); 
    ---Purpose:  Print on the stream  o  information about the object

fields
    myIsDone    : Boolean         from  Standard; 
    myHasResult : Boolean         from  Standard;     
    myBSplCurve : BSplineCurve    from  Geom; 
    myMaxError  : Real            from  Standard; 
    
end Curve3d;
