-- Created on: 1997-04-18
-- Created by: JLF, CAL
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


deferred class Plotter from Graphic3d inherits TShared from MMgt

	---Version:

	---Purpose: This class allows the definition of a plotter

	---Keywords:

	---Warning:
	---References:

uses

	DataStructureManager	from Graphic3d

raises

	PlotterDefinitionError	from Graphic3d

is

	Initialize
	---Level: Public
	---Purpose: Initialise the constructor of the plotter.
	--  Warning: Raises InitialisationError if the initialisation
	--	    of the plotter failed.
	raises PlotterDefinitionError from Graphic3d;
	-- if the initialisation of the plotter failed.

	Destroy ( me     : mutable )
		is virtual;
	---Level: Public
	---Purpose: Deletes the plotter <me>.
	---C++: alias ~

	---------------------------------------------------
	-- Category: Methods to modify the class definition
	---------------------------------------------------

	BeginPlot ( me		: mutable;
		    aProjector	: DataStructureManager from Graphic3d )
        	returns Boolean from Standard
        	raises PlotterDefinitionError from Graphic3d
		is virtual;
        ---Level: Public
	---Purpose:
        --  Warning: Returns Standard_True if plotting is enabled in the view.
        --	    Raises PlotterDefinitionError from Graphic3d
        --	    if plotting has already started.
        ---Category: Methods to modify the class definition

	EndPlot ( me	: mutable )
        	raises PlotterDefinitionError from Graphic3d
		is virtual;
        ---Level: Public
        ---Purpose: Stops the plotting.
        --  Warning: Raises PlotterDefinitionError from Graphic3d
        --	    if plotting has not started yet.
        ---Category: Methods to modify the class definition

	----------------------------
	-- Category: Inquire methods
	----------------------------

	PlottingState ( me )
		returns Boolean from Standard
		is deferred;
        ---Level: Public
        ---Purpose: 
        ---Category: Inquire methods

--

fields

--
-- Class	:	Graphic3d_Plotter
--
-- Purpose	:	Declaration of variables specific to plotters
--
-- Reminder	:	A plotter 

	-- the update display mode
	MyPlottingState		:	Boolean from Standard is protected;

end Plotter from Graphic3d;
