-- Created on: 1993-01-11
-- Created by: CKY / Contract Toubro-Larsen ( Arun MENON )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Node from IGESAppli  inherits IGESEntity

        ---Purpose: defines Node, Type <134> Form <0>
        --          in package IGESAppli
        --          Geometric point used in the definition of a finite element.

uses

    	XYZ  from gp,
	Pnt  from gp,
        TransfEntity         from IGESData,
        TransformationMatrix from IGESGeom

is

        Create returns mutable Node;

        -- Specific Methods pertaining to the class

        Init (me           : mutable;
              aCoord       : XYZ;
              aCoordSystem : TransformationMatrix);
        ---Purpose : This method is used to set the fields of the class Node
        --       - aCoord       : Nodal Coordinates
        --       - aCoordSystem : the Nodal Displacement Coordinate
        --                        System Entity (default 0 is Global 
        --                        Cartesian Coordinate system)

        Coord (me) returns Pnt;
        ---Purpose : returns the nodal coordinates

        System (me) returns TransfEntity;
        ---Purpose : returns TransfEntity if a Nodal Displacement Coordinate
        --           System Entity is defined
        -- else (for Global Cartesien) returns Null Handle

    	SystemType (me) returns Integer;
	---Purpose : Computes & returns the Type of Coordinate System :
	-- 0 GlobalCartesian, 1 Cartesian, 2 Cylindrical, 3 Spherical

        TransformedNodalCoord (me) returns Pnt;
        ---Purpose : returns the Nodal coordinates after transformation

fields

--
-- Class    : IGESAppli_Node
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class Node.
--
-- Reminder : A Node instance is defined by :
--            - Nodal Coordinates
--            - the Nodal Displacement Coordinate System Entity

        theCoord  : XYZ;
        theSystem : TransformationMatrix;

end Node;
