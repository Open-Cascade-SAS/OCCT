-- Created on: 1998-07-08
-- Created by: Stephanie HUMEAU
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred  class TrihedronWithGuide from GeomFill  
inherits TrihedronLaw from GeomFill

	---Purpose: To define Trihedron along one Curve with a guide
	--          
	--          
	--          
      
uses 
    HCurve from  Adaptor3d, 
    Real   from  Standard,
    Pnt    from  gp

raises 
    OutOfRange,  NotImplemented   

is  
     
    Guide(me) 
    returns  HCurve  from  Adaptor3d 
    is  deferred;  
     
    Origine(me  :  mutable; 
    	    Param1  :  Real; 
    	    Param2  :  Real) 
    is deferred;
          
    CurrentPointOnGuide(me) 
     ---Purpose: Returns the current point on guide
     --          found by D0, D1 or D2.
    returns  Pnt from gp;

fields 
    myGuide  :  HCurve  from  Adaptor3d  is  protected; 
    myTrimG  :  HCurve  from  Adaptor3d  is  protected; 
    myCurPointOnGuide : Pnt from gp      is  protected;

end TrihedronWithGuide;
    
