-- Created on: 1993-01-27
-- Created by: Isabelle GRIGNON
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class PolyArc from IntPatch

inherits Polygo from IntPatch

uses Box2d         from Bnd,
     Pnt2d         from gp,
     Array1OfPnt2d from TColgp,
     Array1OfReal  from TColStd,
     HCurve2d from Adaptor2d

raises ConstructionError from Standard

is

    Create(A: HCurve2d from Adaptor2d; NbSample: Integer from Standard; 
    	   Pfirst,Plast : Real from Standard;
           BoxOtherPolygon: Box2d from Bnd)

    	---Purpose: Creates the polygon of the arc A on the surface S.
    	--          The arc is limited by the parameters Pfirst and Plast.
    	--          None of these parameters can be infinite.

    	returns PolyArc from IntPatch
	
	raises ConstructionError from Standard;
    	--- This exception is raised if Pfirst=RealFirst or Plast=RealLast or
    	--  NbSample<=1.

    Closed(me)                   returns Boolean from Standard is redefined virtual;

    NbPoints(me)                 returns Integer;
 
    Point(me; Index : Integer)   returns Pnt2d from gp;
                                      	    	 
    Parameter(me ; Index : Integer) returns Real from Standard;
     
    SetOffset(me:in out;  OffsetX,OffsetY: Real from Standard);
       
		
fields

    brise  : Array1OfPnt2d from TColgp;
    param  : Array1OfReal  from TColStd;
    offsetx: Real          from Standard;
    offsety: Real          from Standard;
    ferme  : Boolean       from Standard;

end PolyArc;
