-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class CartesianTransformationOperator from StepGeom 

inherits GeometricRepresentationItem from StepGeom 
-- WARNING : Multiple EXPRESS inheritance
-- Not yet automaticly managed
-- inherits FunctionallyDefinedTransformation from StepGeom 

uses

	Direction from StepGeom, 
	CartesianPoint from StepGeom, 
	Real from Standard, 
	Boolean from Standard, 
	HAsciiString from TCollection
is

	Create returns mutable CartesianTransformationOperator;
	---Purpose: Returns a CartesianTransformationOperator


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      hasAaxis1 : Boolean from Standard;
	      aAxis1 : mutable Direction from StepGeom;
	      hasAaxis2 : Boolean from Standard;
	      aAxis2 : mutable Direction from StepGeom;
	      aLocalOrigin : mutable CartesianPoint from StepGeom;
	      hasAscale : Boolean from Standard;
	      aScale : Real from Standard) is virtual;

	-- Specific Methods for Field Data Access --

	SetAxis1(me : mutable; aAxis1 : mutable Direction);
	UnSetAxis1 (me:mutable);
	Axis1 (me) returns mutable Direction;
	HasAxis1 (me) returns Boolean;
	SetAxis2(me : mutable; aAxis2 : mutable Direction);
	UnSetAxis2 (me:mutable);
	Axis2 (me) returns mutable Direction;
	HasAxis2 (me) returns Boolean;
	SetLocalOrigin(me : mutable; aLocalOrigin : mutable CartesianPoint);
	LocalOrigin (me) returns mutable CartesianPoint;
	SetScale(me : mutable; aScale : Real);
	UnSetScale (me:mutable);
	Scale (me) returns Real;
	HasScale (me) returns Boolean;

fields

	axis1 : Direction from StepGeom;   -- OPTIONAL can be NULL
	axis2 : Direction from StepGeom;   -- OPTIONAL can be NULL
	localOrigin : CartesianPoint from StepGeom;
	scale : Real from Standard;   -- OPTIONAL can be NULL
	hasAxis1 : Boolean from Standard;
	hasAxis2 : Boolean from Standard;
	hasScale : Boolean from Standard;

end CartesianTransformationOperator;
