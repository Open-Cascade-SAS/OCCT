-- Created on: 1991-04-03
-- Created by: Remi GILET
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Lin2dTanObl

from GccAna

	---Purpose: This class implements the algorithms used to 
	--          create 2d line tangent to a circle or a point and 
	--          making an angle with a line.
        --          The angle is in radians.
        --          The origin of the solution is the tangency point
        --          with the first argument.
        --          Its direction is making an angle Angle with the 
        --          second argument.

--inherits Storable from Standard

uses Lin2d            from gp, 
     Pnt2d            from gp, 
     QualifiedCirc    from GccEnt,
     Array1OfReal     from TColStd,
     Array1OfLin2d    from TColgp,
     Array1OfPnt2d    from TColgp,
     Position         from GccEnt,
     Array1OfPosition from GccEnt

raises OutOfRange        from Standard,
       BadQualifier      from GccEnt,
       NotDone           from StdFail

is

---------------------------------------------------------------------------

Create (ThePoint  : Pnt2d from gp      ;
        TheLine   : Lin2d from gp      ;
        TheAngle  : Real  from Standard) returns Lin2dTanObl;
    	---Purpose: This class implements the algorithms used to 
    	--          create 2d line passing through a point and 
    	--          making an angle with a line.

Create (Qualified1 : QualifiedCirc from GccEnt  ;
        TheLine    : Lin2d         from gp      ;
        TheAngle   : Real          from Standard) returns Lin2dTanObl 
raises BadQualifier;
    	---Purpose: This class implements the algorithms used to 
    	--          create 2d line tangent to a circle and 
    	--          making an angle with a line.
    	--          Exceptions
    	--          GccEnt_BadQualifier if a qualifier is inconsistent with
    	--          the argument it qualifies (for example, enclosed for a circle).

IsDone(me) returns Boolean from Standard
is static;
    	---Purpose : Returns True if the algorithm succeeded.
    	--           Note: IsDone protects against a failure arising from a
    	--           more internal intersection algorithm, which has reached
    	--           its numeric limits.
    
NbSolutions(me) returns Integer from Standard
   	---Purpose : Returns the number of  of lines, representing solutions computed by this algorithm.
    	--           Raises NotDone if the construction algorithm didn't succeed.

raises NotDone
is static;
  
ThisSolution(me                           ;
    	     Index : Integer from Standard) returns Lin2d 
    	---Purpose: Returns the solution number Index.
    	--          Be careful: the Index is only a way to get all the 
    	--          solutions, but is not associated to theses outside the 
    	--          context of the algorithm-object.
    	-- raises NotDone if the construction algorithm didn't succeed.
   	--          It raises OutOfRange if Index is greater than the   number of solutions.
raises OutOfRange, NotDone
is static;
 
WhichQualifier(me                                  ;
    	       Index   :     Integer  from Standard;
	       Qualif1 : out Position from GccEnt  )
raises OutOfRange, NotDone
is static;
    	---Purpose: Returns the qualifier Qualif1 of the tangency argument
    	-- for the solution of index Index computed by this algorithm.
    	-- The returned qualifier is:
    	-- -   that specified at the start of construction when the
    	--   solutions are defined as enclosing or outside with
    	--   respect to the argument, or
    	-- -   that computed during construction (i.e. enclosing or
    	--   outside) when the solutions are defined as unqualified
    	--   with respect to the argument, or
    	-- -   GccEnt_noqualifier if the tangency argument is a point.
    	--  Exceptions
    	-- Standard_OutOfRange if Index is less than zero or
    	-- greater than the number of solutions computed by this algorithm.
    	-- StdFail_NotDone if the construction fails. 

Tangency1(me                                     ;
          Index         : Integer   from Standard;
          ParSol,ParArg : out Real  from Standard;
          PntSol        : out Pnt2d from gp      )
    	---Purpose : Returns informations about the tangency point between the 
    	--           result number Index and the first argument.
    	--           ParSol is the intrinsic parameter of the point ParSol on 
    	--           the solution curv.
    	--           ParArg is the intrinsic parameter of the point ParArg on 
    	--           the argument curv. Raises NotDone if the construction algorithm 
    	--          didn't succeed.
    	--          It raises OutOfRange if Index is greater than the  number of solutions.
raises OutOfRange, NotDone
is static;
  

Intersection2 (me                                     ;
               Index         : Integer   from Standard;
               ParSol,ParArg : out Real  from Standard;
               PntSol        : out Pnt2d from gp      )
    	---Purpose : Returns informations about the intersection between the
    	--           result number Index and the third argument.
    	-- Raises NotDone if the construction algorithm  didn't succeed.
    	--          It raises OutOfRange if Index is greater than the number of solutions.
raises OutOfRange, NotDone
is static;
  
fields

    WellDone : Boolean from Standard;
    	---Purpose : True if the algorithm succeeded.

    NbrSol   : Integer from Standard;
    	---Purpose : The number of possible solutions. We have to decide about the
    	--           status of the multiple solutions...

    linsol   : Array1OfLin2d from TColgp;
    	---Purpose : The solutions.

    qualifier1 : Array1OfPosition from GccEnt;
    	---Purpose: The qualifiers of the first argument.

    pnttg1sol   : Array1OfPnt2d from TColgp;
    	---Purpose: The tangency point between the solution and the first argument on 
   	-- the solution.

    pntint2sol   : Array1OfPnt2d from TColgp;
    	---Purpose: The tangency point between the solution and the second argument on 
    	-- the solution.

    par1sol   : Array1OfReal from TColStd;
    	---Purpose: The parameter of the tangency point between the solution and the 
    	-- first argument on the solution.

    par2sol   : Array1OfReal from TColStd;
       	---Purpose: The parameter of the tangency point between the solution and the 
	-- second argument on the solution.

    pararg1   : Array1OfReal from TColStd;
    	---Purpose: The parameter of the tangency point between the solution and the first 
    	-- argument on the first argument.

    pararg2   : Array1OfReal from TColStd;
    	---Purpose: The parameter of the tangency point between the solution and the second
    	-- argument on the second argument.

end Lin2dTanObl;

