-- Created on: 1997-10-22
-- Created by: Jean-Louis Frenkel
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


private class Reference from CDM  inherits Transient from Standard

uses Document from CDM, DocumentPointer from CDM, Application from CDM, MetaData from CDM

is

    Create(aFromDocument: Document from CDM; aToDocument: Document from CDM; aReferenceIdentifier: Integer from Standard; aToDocumentVersion: Integer from Standard)
    returns mutable Reference from CDM
    is private;

    Create(aFromDocument: Document from CDM; aMetaData: MetaData from CDM; aReferenceIdentifier: Integer from Standard; anApplication: Application from CDM; aToDocumentVersion: Integer from Standard; UseStorageConfiguration: Boolean from Standard)
    returns mutable Reference from CDM
    is private;
    

    

    FromDocument(me: mutable) returns Document from CDM;

    ToDocument(me: mutable) returns Document from CDM;
	    
    ReferenceIdentifier(me: mutable) returns Integer from Standard;
    
    
---Category: methods to modifiy the reference.


    Update(me: mutable; aMetaData: MetaData from CDM)
    is private;

    IsUpToDate(me) returns Boolean from Standard
    is private;
    ---Purpose: compares the actual document version with the 
    --          document version at the creation of the reference
    SetIsUpToDate(me: mutable)
    is private;

    UnsetToDocument(me: mutable; aMetaData: MetaData from CDM; anApplication: Application from CDM) is private;
    
    IsOpened(me) returns Boolean from Standard is private;
    ---Purpose: returns  true if the  ToDocument has been retrieved
    --          and opened.

    DocumentVersion(me) returns Integer from Standard;
    
    IsReadOnly(me) returns Boolean from Standard;

    Document(me) returns Document from CDM
    is private;

    MetaData(me) returns MetaData from CDM
    is private;
    
    Application(me) returns Application from CDM
    is private;

    UseStorageConfiguration(me) returns Boolean from Standard
    is private;
    
    IsInSession(me) returns Boolean from Standard
    is private;
    
    IsStored(me) returns Boolean from Standard
    is private;
    
fields

    myToDocument: Document from CDM;
    myFromDocument: DocumentPointer from CDM;
    myReferenceIdentifier: Integer from Standard;
    
    myApplication: Application from CDM;
    myMetaData: MetaData from CDM;
    myDocumentVersion: Integer from Standard;    
    myUseStorageConfiguration: Boolean from Standard;
friends class Document from CDM
end Reference from CDM;
