-- Created on: 1994-04-01
-- Created by: Modelistation
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



package BRepTopAdaptor 

	---Purpose: 
	--          
	--          
	--          *** Class2d    : Low level algorithm for 2d classification
	--          
	--          *** FClass2d   : 2d classification on a Face from TopoDS
	--                           A face is first loaded and then every 
	--                           classification is computed as a rejection.                        
	--                           (call BRepClass algorithms if necessary,
	--                           ie, when the rejection is not efficient)
	--                           
	--          *** TopolTool :  Several tools used by the intersection
	--                           algorithm and topology.
	--         
	--          

	---Level: Internal

uses Adaptor3d, TopExp, TopoDS, BRepAdaptor, gp, TopAbs,  Adaptor2d  ,
     TColgp,TColStd,TCollection,TopTools, CSLib

is

    --class Class2d;

    alias SeqOfPtr is SequenceOfAddress from TColStd;

    class FClass2d; 

    class HVertex; -- inherits HVertex from Adaptor3d

    class TopolTool; -- inherits TopolTool from Adaptor3d
    


    --- the folowing classes are used to compute and store 
    --  informations on shapes. ( TopolTool , Bnd_Box ... )
    
    class Tool; 
    
    class MapOfShapeTool  instantiates DataMap from TCollection
        (Shape          from TopoDS,
         Tool           from BRepTopAdaptor,
         ShapeMapHasher from TopTools);


end BRepTopAdaptor;
