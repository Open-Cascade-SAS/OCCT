-- Created on: 1994-12-02
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class ModifyShape from BRepBuilderAPI inherits MakeShape from BRepBuilderAPI

	---Purpose: Implements   the  methods   of MakeShape for   the
	--          constant  topology modifications.  The methods are
	--          implemented  when the modification uses a Modifier
	--          from BRepTools. Some of  them have to be redefined
	--          if  the  modification is  implemented with another
	--          tool (see Transform from BRepBuilderAPI for example).
    	-- The BRepBuilderAPI package provides the following
    	-- frameworks to perform modifications of this sort:
    	-- -   BRepBuilderAPI_Copy to produce the copy of a shape,
    	-- -   BRepBuilderAPI_Transform and
    	--   BRepBuilderAPI_GTransform to apply a geometric
    	--   transformation to a shape,
    	-- -   BRepBuilderAPI_NurbsConvert to convert the
    	--   whole geometry of a shape into NURBS geometry,
    	-- -   BRepOffsetAPI_DraftAngle to build a tapered shape.

uses
    Shape             from TopoDS,
    Face              from TopoDS,
    Edge              from TopoDS,
    ShapeModification from BRepBuilderAPI,
    ListOfShape       from TopTools,
    
    Modifier          from BRepTools,
    Modification      from BRepTools

raises
    NullObject   from Standard,
    NoSuchObject from Standard
is

    Initialize;
	---Purpose: Empty constructor.
    

    Initialize(S:Shape from TopoDS);
	---Purpose: Initializes the modifier with  the Shape  <S>, and
	--          set the field <myInitialShape> to <S>.


    Initialize(M: Modification from BRepTools);
	---Purpose: Set the field <myModification> with <M>.


    Initialize(S: Shape from TopoDS; M: Modification from BRepTools);
	---Purpose: Initializes the modifier with  the Shape  <S>, and
	--          set the field <myInitialShape> to <S>, and set the
	--          field <myModification> with  <M>, the performs the
	--          modification.


    DoModif(me: in out; S: Shape from TopoDS)
	---Purpose: Performs the previously  given modification on the
	--          shape <S>.
    
    	raises NullObject from Standard
	--- The  exception is raised if no modification has been given.
	is static protected;


    DoModif(me: in out; M: Modification from BRepTools)
	---Purpose: Performs the  modification   <M> on a   previously
	--          given shape.
    
    	raises NullObject from Standard
	--- The  exception is raised if no shape has been given.
	is static protected;


    DoModif(me: in out; S: Shape from TopoDS;
                        M: Modification from BRepTools)
	---Purpose: Performs the  modification <M> on the shape <S>.
    
    	is static protected;


--- Private implementation method

    DoModif(me: in out)
    
	is static private;

---Category: Querying isg-attention il faudrait passer en modified que
--            les faces  dont les  bornes  sont modifiees et les faces
--           inclinees en generated (pas disponible aujourd 'hui dans BRepTools_modifier
--           a reprendre
--           
    Modified (me: in out; S : Shape from TopoDS)
    	---Purpose: Returns the list  of shapes modified from the shape
    	--          <S>. 
        ---C++: return const & 
        ---Level: Public
    returns ListOfShape from TopTools
    is redefined virtual;

 
    ModifiedShape(me; S: Shape from TopoDS)
    	returns Shape from TopoDS
	---Purpose: Returns the modified shape corresponding to <S>.
    	-- S can correspond to the entire initial shape or to its subshape.
    	-- Exceptions
    	-- Standard_NoSuchObject if S is not the initial shape or
    	-- a subshape of the initial shape to which the
    	-- transformation has been applied. Raises NoSuchObject from Standard
    	-- if S is not the initial shape or a sub-shape
    	-- of the initial shape.
	---C++: return const&
	raises NoSuchObject from Standard
             
    is virtual;

fields

    myModifier     : Modifier     from BRepTools is protected;
    myInitialShape : Shape        from TopoDS    is protected;
    myModification : Modification from BRepTools is protected;
    
end ModifyShape;
