-- Created on: 1992-08-20
-- Created by: Christophe MARION
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Coincidence from HLRAlgo

	---Purpose: The Coincidence class is used in an Inteference to
	--          store informations on the "hiding" edge.
	--          
	--          2D  Data : The  tangent  and the  curvature of the
	--          projection of the edge  at the intersection point.
	--          This is necesserary  when the intersection  is  at
	--          the extremity of the edge.
	--          
	--          3D   Data  :  The   state of  the   edge  near the
	--          intersection   with  the face (before  and after).
	--          This is necessary  when the  intersection is  "ON"
	--          the face.

uses
    Integer from Standard,
    Real    from Standard,
    State   from TopAbs

is
    Create returns Coincidence from HLRAlgo;
    
    Set2D(me : in out; FE    : Integer from Standard;
                       Param : Real    from Standard)
    	---C++: inline
    is static;
    
    SetState3D(me : in out; stbef,staft : State from TopAbs)
    	---C++: inline
    is static;

    Value2D(me; FE    : out Integer from Standard;
                Param : out Real    from Standard)
    	---C++: inline
    is static;
    
    State3D(me; stbef,staft : out State from TopAbs)
    	---C++: inline
    is static;
	    
fields
    myFE    : Integer from Standard;
    myParam : Real    from Standard;
    myStBef : State from TopAbs;
    myStAft : State from TopAbs;

end Coincidence;
