-- Created on: 1996-10-21
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package TestTopOpe

uses 
 
    Draw,
    TopOpeBRepBuild,
    TopOpeBRepDS,
    TopoDS
    
is

    AllCommands(I : in out Interpretor from Draw);
    ---Purpose: Defines all Top. Ope. test commands

    TOPOCommands(I : in out Interpretor from Draw);

    BOOPCommands(I : in out Interpretor from Draw);

    HDSCommands(I : in out Interpretor from Draw);
    ---Purpose: commands on a HDS involved in topological operations

    CurrentHB(HDS : HBuilder from TopOpeBRepBuild);
    ---Purpose : Defines the HBuilder on which BOOPCommands will operate.

    CurrentDS(HDS : HDataStructure from TopOpeBRepDS);
    ---Purpose : Defines the HDS on which HDSCommands/BOOPCommands will operate.

    Shapes(S1,S2 : Shape from TopoDS);
    ---Purpose: Defines current shapes of current topological operation

    MesureCommands(I : in out Interpretor from Draw);

    CORCommands(I : in out Interpretor from Draw);

    DSACommands(I : in out Interpretor from Draw);

    OtherCommands(I : in out Interpretor from Draw);

    Factory (theDI : out Interpretor from Draw);
    ---Purpose: Loads all Draw commands of TKDrawDEB. Used for plugin.

end TestTopOpe;
