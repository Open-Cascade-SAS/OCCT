-- Created on: 1996-10-23
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class FFDumper from TopOpeBRep inherits TShared from MMgt

uses

    DataMapOfShapeInteger from TopTools,
    PFacesFiller from TopOpeBRep,
    LineInter from TopOpeBRep, 
    VPointInter from TopOpeBRep,
    VPointInterIterator from TopOpeBRep,
    Kind from TopOpeBRepDS,    
    Shape from TopoDS,
    Face from TopoDS
    
is 

    Create(PFF:PFacesFiller) returns mutable FFDumper from  TopOpeBRep; 
    Init(me:mutable;PFF:PFacesFiller); 
    DumpLine(me:mutable;I:Integer);
    DumpLine(me:mutable;L:LineInter);
    DumpVP(me:mutable;VP:VPointInter);
    DumpVP(me:mutable;VP:VPointInter;ISI:Integer); 
    ExploreIndex(me;S:Shape;ISI:Integer) returns Integer; 
    DumpDSP(me;VP:VPointInter;GK:Kind;G:Integer;newinDS:Boolean);
    PFacesFillerDummy(me) returns PFacesFiller;

fields

    myPFF:PFacesFiller from TopOpeBRep;
    myF1,myF2:Face from TopoDS;
    myEM1,myEM2:DataMapOfShapeInteger from TopTools; 
    myEn1,myEn2:Integer;
    myLineIndex : Integer;

end FFDumper from TopOpeBRep;
