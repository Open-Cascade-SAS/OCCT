-- File:	BOPTools_IteratorOfCoupleOfShape.cdl
-- Created:	Mon Nov 27 16:31:08 2000
-- Author:	Michael KLOKOV
--		<mkk@nizhnox.nnov.matra-dtv.fr>
---Copyright:	 Matra Datavision 2000

class IteratorOfCoupleOfShape from BOPTools

    	---Purpose: The class IteratorOfCoupleOfShape provides the iteration
    	---         on the couples of shapes stored in ShapesDataStructure 
	---         according to the given types of shapes and
	---         status of their intersection.
	---         The statuses are stored in 2 dimension array.

uses
    ShapeEnum from TopAbs,
    HArray2OfIntersectionStatus from BOPTools,
    PShapesDataStructure from BooleanOperations,
    IntersectionStatus from BOPTools, 
    ListOfCoupleOfInteger from BOPTools, 
    ListIteratorOfListOfCoupleOfInteger from BOPTools,    
    NoSuchObject from Standard 
    
raises NoSuchObject from Standard 

is

    Create  
    	returns IteratorOfCoupleOfShape from BOPTools;
    	---Purpose: 
    	--- Empty Constructor 
    	---

    Create(PDS: PShapesDataStructure from BooleanOperations;
	   Type1: ShapeEnum from TopAbs;
    	   Type2: ShapeEnum from TopAbs)
    	returns IteratorOfCoupleOfShape from BOPTools;
    	---Purpose: 
    	--- Initializes iterator by ShapesDataStructure and
    	--- shape types
	---

    Destroy(me: in out) is virtual;
        ---C++: alias "Standard_EXPORT virtual ~BOPTools_IteratorOfCoupleOfShape(){Destroy();}"

    Initialize(me: in out; Type1: ShapeEnum from TopAbs;
    	    	    	   Type2: ShapeEnum from TopAbs) 
							    
	raises NoSuchObject from Standard 
    	is virtual;
    	---Purpose: 
    	--- Initializes iterator with shape types. 
    	--- The iterator uses PDS assigned in constructor or in SetDataStructure().
    	--- Raises the exception if myPDS is null.
	---


    SetDataStructure(me: in out; PDS: PShapesDataStructure from BooleanOperations)
    	raises
	    NoSuchObject from Standard;
    	---Purpose: 
    	--- Initialize iterator with ShapeDataStructure.
	---
    

    More(me)  
    	returns Boolean from Standard 
    	is virtual;
	---Purpose:
	--- Returns True if there are still not
	--- treated couples of shapes
	---
    
    Next(me: in out) 
    	is virtual;
    	---Purpose:
	--- Moves to the next couple of iteration
	---
    
    Current(me; Index1: in out Integer from Standard;
    	    	Index2: in out Integer from Standard;
    	    	WithSubShape: out Boolean from Standard) 
    	is virtual;
    	---Purpose: 
    	--- Returns current couple of indices and
    	--- flag WithSubShape which is true 
    	--- if bounding boxes of subshapes
    	--- are intersected
	---

    ListOfCouple(me) 
    	returns  ListOfCoupleOfInteger from BOPTools;  
    	---C++:  return const &
	---Purpose:
	--- Returns a list of couples of shape indices
	--- according to shape types by which
	--- the iterator was initialized
	---
	
    MoreP(me)  
    	returns Boolean from Standard   
    	is protected;
    
    NextP(me: in out) 
    	is protected;
    
    CurrentP(me;Index1: in out Integer from Standard;
    	    	Index2: in out Integer from Standard)
    	raises NoSuchObject from Standard 
    	is protected;

    SetIntersectionStatus(me: in out; Index1: Integer from Standard;
		        	      Index2: Integer from Standard;
    	    	    	    	      theStatus: IntersectionStatus from BOPTools);
    	---Purpose:
	--- Sets status to array according to Index1 and Index2
	---

    GetTableOfIntersectionStatus(me)
    	returns HArray2OfIntersectionStatus from BOPTools;
	---C++: return const &
	---Purpose:
	--- Returns 2 dimension array of intersection statuses
	---
    
    DumpTableOfIntersectionStatus(me);
    	---Purpose:
	--- For internal use
	---
    
fields
    myPDS: PShapesDataStructure from BooleanOperations is protected;
    myTableOfStatus: HArray2OfIntersectionStatus from BOPTools is protected;
    myCurrentIndex1: Integer from Standard is protected;
    myCurrentIndex2: Integer from Standard is protected;
    myType1:         ShapeEnum from TopAbs is protected;
    myType2:         ShapeEnum from TopAbs is protected;
--  
    myFirstLowerIndex :Integer from Standard is protected; 
    myFirstUpperIndex :Integer from Standard is protected; 
    mySecondLowerIndex:Integer from Standard is protected; 
    mySecondUpperIndex:Integer from Standard is protected; 
    myListOfCouple    :ListOfCoupleOfInteger from BOPTools is protected;  
    myIterator        :ListIteratorOfListOfCoupleOfInteger from BOPTools is protected;  
--  
end IteratorOfCoupleOfShape from BOPTools;
