-- Created on: 2002-10-29
-- Created by: Michael SAZONOV
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class ADriver from BinMDF inherits TShared from MMgt

        ---Purpose: Attribute Storage/Retrieval Driver.

uses
    ExtendedString   from TCollection,
    MessageDriver    from CDM,
    AsciiString      from TCollection,
    Attribute        from TDF,
    RRelocationTable from BinObjMgt,
    SRelocationTable from BinObjMgt,
    Persistent       from BinObjMgt

is
    Initialize (theMsgDriver: MessageDriver from CDM;
                theName     : CString from Standard = NULL);

    NewEmpty    (me)
        returns mutable Attribute from TDF
        is deferred;
        ---Purpose: Creates a new attribute from TDF.

    SourceType  (me) returns Type from Standard;
        ---C++: return const &
	---C++: inline
        ---Purpose: Returns the type of source object,
        --          inheriting from Attribute from TDF.

    TypeName    (me)
        returns AsciiString from TCollection
        is static;
        ---C++: return const &
	---C++: inline
        ---Purpose: Returns the type name of the attribute object

    Paste       (me; aSource     : Persistent from BinObjMgt;
                     aTarget     : mutable Attribute from TDF;
                     aRelocTable : out RRelocationTable from BinObjMgt)
        returns Boolean from Standard is deferred;
        ---Purpose: Translate the contents of <aSource> and put it
        --          into <aTarget>, using the relocation table
        --          <aRelocTable> to keep the sharings.

    Paste       (me; aSource     : Attribute from TDF;
                     aTarget     : in out Persistent from BinObjMgt;
                     aRelocTable : out SRelocationTable from BinObjMgt)
        is deferred;
        ---Purpose: Translate the contents of <aSource> and put it
        --          into <aTarget>, using the relocation table
        --          <aRelocTable> to keep the sharings.

    WriteMessage (me; theMessage : ExtendedString from TCollection);
        ---Purpose: Send message to Application (usually when error occurres)

fields

    myMessageDriver : MessageDriver from CDM;
    myTypeName      : AsciiString   from TCollection is protected;

end ADriver;
