-- Created on: 1992-05-27
-- Created by: Remi LEQUETTE
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.





class TEdge from BRep inherits TEdge from TopoDS

	---Purpose: The TEdge from BRep is  inherited from  the  TEdge
	--          from TopoDS. It contains the geometric data.
	--          
	--          The TEdge contains :
	--           
	--           * A tolerance.
	--           
	--           * A same parameter flag.
	--           
	--           * A same range flag.
	--           
	--           * A Degenerated flag.
	--           
	--           *  A  list   of curve representation.

uses
    TShape                    from TopoDS,
    ListOfCurveRepresentation from BRep

is
    Create returns mutable TEdge from BRep;
	---Purpose: Creates an empty TEdge.
	
    Tolerance(me) returns Real
	---C++: inline
    is static;
    	
    Tolerance(me : mutable; T : Real)
	---C++: inline
    is static;
    
    UpdateTolerance(me : mutable; T : Real)
	---Purpose: Sets the tolerance  to the   max  of <T>  and  the
	--          current  tolerance.
	--          
	---C++: inline
    is static;
    
    SameParameter(me) returns Boolean
    is static;
    
    SameParameter(me : mutable; S : Boolean)
    is static;
    
    SameRange(me) returns Boolean
    is static;
    
    SameRange(me : mutable; S : Boolean)
    is static;
    
    Degenerated(me) returns Boolean
    is static;
    
    Degenerated(me : mutable; S : Boolean)
    is static;
    
    Curves(me) returns ListOfCurveRepresentation from BRep
	---C++: return const &
	---C++: inline
    is static;
    
    ChangeCurves(me : mutable) returns ListOfCurveRepresentation from BRep
	---C++: return &
	---C++: inline
    is static;
    
    EmptyCopy(me) returns mutable TShape from TopoDS;
	---Purpose: Returns a copy  of the  TShape  with no sub-shapes.
    
fields

    myTolerance     : Real;
    myFlags         : Integer;
    myCurves        : ListOfCurveRepresentation from BRep;

end TEdge;
