-- Created on: 1996-05-31
-- Created by: Laurent BUCHARD
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package IntCurvesFace

----------------------------------------------------------------------
-- This package provide algorithms to  compute the intersection points
-- between a Face [a  Shape] and a set of  curves (The face [shape] is
-- loaded, then for each curve is given to compute the intersection).
-- 
-- Intersector [  ShapeIntersector ] can be  used when the caller have
-- to intersect more than one curve with the face [the shape].
-- 
-- 
-- If there is  only one curve, or  if  the face  has no restrictions,
-- someother algorithms can be called. 
--    
-- see for example the packages : 
-- 
--      ** BRepIntCurveSurface :  ( One Curve   <->   One  Shape )
--      ** IntCurveSurface     :  ( One Curve   <->   One  Surface)
--     
----------------------------------------------------------------------


uses 
    gp              ,
    TopAbs          ,
    TopoDS          ,
    BRepTopAdaptor  ,
    BRepAdaptor     ,
    Adaptor3d         ,
    Bnd             ,
    IntCurveSurface ,
    TColStd         ,
    GeomAbs
    
is

    class Intersector;            -- Intersection between a Face and a set of curves 
    
    class ShapeIntersector;       -- Intersection between a Shape and a set of curves 
                                  -- Note ( has an empty constructor )
    
end;

