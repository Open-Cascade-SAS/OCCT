-- Created on: 1999-10-11
-- Created by: Atelier CAS2000
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package  BRepOffsetAPI 

uses   
    Standard, 
    StdFail,
    gp, 
    GeomAbs,
    Geom,
    GeomFill,
    Approx,
    TopoDS,
    TopTools, 
    BRepAlgo,
    BRepBuilderAPI, 
    BRepSweep, 
    BRepPrimAPI,  	     
    BRepFill, 
    Law, 
    Draft, 
    BRepOffset, 
     
    TColStd,
    TCollection

is 


    --
    -- Sweeping
    -- 

    class MakePipe;        ---  inherits MakeSweep from BRepPrimAPI    
	---Purpose: To create shape by pipe
	          
    class MakePipeShell;  ---  inherits MakeSweep from BRepPrimAPI
    	---Purpose: Numerous posibilities to create shell by sweeping          
     


    class  MakeDraft; ---  inherits MakeShape from BRepBuilderAPI
    
    class DraftAngle; ---  inherits MakeShape from BRepBuilderAPI




    class FindContigousEdges;
      ---Purpose: find the contigous edges of shapes for control
      --          (continuity C0, C1, ...)

    alias Sewing  is  Sewing from BRepBuilderAPI;
      ---Purpose: sew the shapes along their common edges
   


    --
    -- Evolved and Offseting
    -- 
    
    class MakeOffset;     ---  inherits MakeShape from BRepBuilderAPI
	---Purpose: Offsets to a set of plane wires.
    
    class MakeOffsetShape; ---  inherits MakeShape from BRepBuilderAPI
    	--Purpose: Offset shape to shells or solids.

    class MakeThickSolid;    ---   inherits MakeOffsetShape from BRepOffsetAPI
	---Purpose: Thick solid to shells or solids.

    class MakeEvolved;    ---  inherits MakeShape from BRepBuilderAPI

 
    --
    -- Construction of Shape through sections.
    -- 

    class ThruSections;	      ---  inherits  MakeShape  from  BRepBuilderAPI

    class NormalProjection ;  ---  inherits  MakeShape  from  BRepBuilderAPI

    class MiddlePath;	      ---  inherits  MakeShape  from  BRepBuilderAPI
    
    -- 
    --   Plate
    --     
    class MakeFilling;  ---  inherits MakeShape from BRepBuilderAPI

	---Purpose: N-Side Filling
	--  This algorithm avoids to build a face from:
	--  * a set of edges defining the bounds of the face and some
	--    constraints the surface of the face has to satisfy
	--  * a set of edges and points defining some constraints
	--    the support surface has to satisfy
	--  * an initial surface to deform for satisfying the constraints
	--  * a set of parameters to control the constraints.
     
    class SequenceOfSequenceOfReal instantiates 
    	Sequence from TCollection (SequenceOfReal from TColStd);

    class SequenceOfSequenceOfShape instantiates 
    	Sequence from TCollection (SequenceOfShape from TopTools);

end;
