-- Created on: 1996-07-26
-- Created by: Maria PUMBORIOS
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



package FilletSurf 

	---Purpose:  This package contains the API giving 
	--           only geometric informations about fillets
	--           for Toyota Project UV4. 
        
uses
    TopoDS,
    TopTools,
    ChFi3d,
    ChFiDS,
    BRepAdaptor,
    Adaptor3d,
    math,
    Geom,
    Geom2d,
    gp,
    StdFail,
    TopAbs
is

---------------------------------------------------------- 
--  enumeration used to describe the status of start and end section
--  of the fillet 
--   TwoExtremityOnEdge
--   OneExtremityOnEdge
--   NoExtremityOnEdge
----------------------------------------------------------
--                                                               
--    
enumeration StatusType  is  TwoExtremityOnEdge, OneExtremityOnEdge, 
                            NoExtremityOnEdge  
end  StatusType;
    
---------------------------------------------------------- 
--  enumeration used to describe the status of the computation of the fillet
-- IsOk  
-- IsNotOk 
-- IsPartial    
--   
----------------------------------------------------------

enumeration StatusDone  is  IsOk, IsNotOk,IsPartial 
                      
end  StatusDone;

---------------------------------------------------------- 
--  enumeration used to describe the  status error  
--   EmptyList 
--   EdgeNotG1 
--   FacesNotG1
--    EdgeNotOnShape    
--    NotSharpEdge
--    PbFilletCompute
----------------------------------------------------------

enumeration ErrorTypeStatus  is  EmptyList, EdgeNotG1,FacesNotG1,EdgeNotOnShape,
                                 NotSharpEdge, PbFilletCompute                    
end  ErrorTypeStatus ;



--  this class is the API giving geometric informations about fillets:
 
    class Builder; 


-- this class is private and is only used by the class Builder:


    private class InternalBuilder;
    

end FilletSurf;
















