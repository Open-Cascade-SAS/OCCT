-- Created by: DAUTRY Philippe
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

--      	----------------------

---Version:	0.0
--Version	Date		Purpose
--		0.0	Sep  8 1997	Creation



deferred class AttributeDelta from TDF inherits TShared from MMgt

	---Purpose: This class discribes the services we need to
	--           implement Delta and Undo/Redo services.
	--           
	--          AttributeDeltas are applied in an unpredictable
	--          order. But by the redefinition of the method
	--          IsNowApplicable, a condition can be verified
	--          before application. If the AttributeDelta is not
	--          yet applicable, it is put at the end of the
	--          AttributeDelta list, to be treated later. If a
	--          dead lock if found on the list, the
	--          AttributeDeltas are forced to be applied in an
	--          unpredictable order.


uses

    Label     from TDF,
    Attribute from TDF
    
is

    Initialize(anAttribute: Attribute from TDF);
    

    Apply(me : mutable)
    	is deferred;
    	---Purpose: Applies the delta to the attribute.
    
    Label(me)
    	returns Label from TDF;
	---Purpose: Returns the label concerned by <me>.

    Attribute(me)
    	returns Attribute from TDF;
	---Purpose: Returns the reference attribute.

    ID(me)
    	returns GUID from Standard;
	---Purpose: Returns the ID of the attribute concerned by <me>.


    ---Category: Miscelleaneous
    --           --------------------------------------------------------------

    Dump(me; OS : in out OStream from Standard)
    	returns OStream from Standard
    	is virtual;
	---Purpose: Dumps the contents.
	--          
	---C++: return &
	---C++: alias operator<<

fields

    myAttribute : Attribute from TDF;
    myLabel     : Label from TDF;

end AttributeDelta;




