-- Created by: DAUTRY Philippe
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

--      	------------------

---Version:	0.0
--Version	Date		Purpose
--		0.0	Feb  4 1998	Creation


class Shape1 from PTopoDS inherits Storable from Standard

    ---Purpose: The PTopoDS_Shape1 is the Persistent view of a TopoDS_Shape.
    --          
    --  a  Shape1 contains :
    --          
    --          - a reference to a TShape1.
    --          
    --          - a Location  to put the TShape1 in  a local coordinate
    --          system.
    --          
    --          - an Orientation.
    --          
    --          It inherits from ExternShareable, so that it can be shared
    --          by other objects located outside the container.
    
uses

    Orientation   from TopAbs,
    TShape1       from PTopoDS,
    Location      from PTopLoc
    
is
    Create returns Shape1 from PTopoDS;
    ---Level: Internal 

    Nullify(me : in out)
    is static;

    TShape(me) returns any TShape1 from PTopoDS
    ---Level: Internal 
    ---C++: return const &
    is static;

    TShape(me : in out; T : TShape1 from PTopoDS)
    ---Level: Internal 
    is static;

    Location(me) returns Location from PTopLoc
    ---Level: Internal 
    is static;
	
    Location(me : in out; L : Location from PTopLoc)
    ---Level: Internal 
    is static;
	
    Orientation(me) returns Orientation from TopAbs
    ---Level: Internal 
    is static;

    Orientation(me: in out; O : Orientation from TopAbs)
    ---Level: Internal 
    is static;
    
fields

    myTShape   : TShape1     from PTopoDS;
    myLocation : Location    from PTopLoc;
    myOrient   : Orientation from TopAbs;

end Shape1;
