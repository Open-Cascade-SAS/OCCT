-- Created on: 1994-03-25
-- Created by: model
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class HVertex from Adaptor3d 

	---Purpose: 


inherits TShared from MMgt

uses Pnt2d       from gp,
     Orientation from TopAbs,
     HCurve2d    from Adaptor2d

is

    Create
    
    	returns mutable HVertex from Adaptor3d;


    Create(P: Pnt2d from gp; Ori: Orientation from TopAbs;
           Resolution: Real from Standard)

    	returns mutable HVertex from Adaptor3d;


    Value(me: mutable)
    
    	returns Pnt2d from gp
    is virtual;


    Parameter(me: mutable; C: HCurve2d from Adaptor2d)
    
    	returns Real from Standard
    is virtual;


    Resolution(me: mutable; C: HCurve2d from Adaptor2d)
    
	---Purpose: Parametric resolution (2d).

    	returns Real from Standard
    is virtual;


    Orientation(me: mutable)
    
    	returns Orientation from TopAbs
    is virtual;


    IsSame(me: mutable; Other: mutable like me)
    
    	returns Boolean from Standard
    is virtual;


fields

    myPnt : Pnt2d       from gp;
    myTol : Real        from Standard;
    myOri : Orientation from TopAbs;

end HVertex;
