-- Created on: 1993-03-10
-- Created by: JCV
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class OffsetCurve from Geom inherits Curve from Geom

    
        ---Purpose :
        --  This class implements the basis services for an offset curve
        --  in 3D space. The Offset curve in this package can be a self
        --  intersecting curve even if the basis curve does not 
        --  self-intersect. The self intersecting portions are not deleted
        --  at the construction time.
        --  An offset curve is a curve at constant distance (Offset) from
        --  a basis curve in a reference direction V. The offset curve 
        --  takes its parametrization from the basis curve.
        --  The Offset curve is in the direction of of the normal N 
        --  defined with the cross product  V^T where the vector T
        --  is given by the first derivative on the basis curve with 
        --  non zero length.
        --  The distance offset may be positive or negative to indicate the
        --  preferred side of the curve :
        --  . distance offset >0 => the curve is in the direction of N
        --  . distance offset >0 => the curve is in the direction of - N
        --  
        --  On the Offset curve :
        --  Value (U) = BasisCurve.Value(U) + (Offset * (T ^ V)) / ||T ^ V||
        --  
        --  At any point the Offset direction V must not be parallel to the
        --  vector T and the vector T must not have null length else the
        --  offset curve is not defined. So the offset curve has not the 
        --  same continuity as the basis curve.
        -- 
        --   Warnings :
        --  
        --  In this package we suppose that the continuity of the offset
        --  curve is one degree less than the continuity of the basis 
        --  curve and we don't check that at any point ||T^V|| != 0.0
        --  
        --  So to evaluate the curve it is better to check that the offset
        --  curve is well defined at any point because an exception could 
        --  be raised. The check is not done in this package at the creation
        --  of the offset curve because the control needs the use of an
        --  algorithm which cannot be implemented in this package.
        -- 
        --  The OffsetCurve is closed if the first point and the last point
        --  are the same (The distance between these two points is lower or
        --  equal to the Resolution sea package gp) . The OffsetCurve can be
        --  closed even if the basis curve is not closed. 


uses Dir      from gp,
     Pnt      from gp,
     Trsf     from gp,
     Vec      from gp,
     Curve    from Geom,
     Geometry from Geom,
     Shape    from GeomAbs


raises ConstructionError   from Standard,
       RangeError          from Standard,
       NoSuchObject        from Standard,
       UndefinedDerivative from Geom,
       UndefinedValue      from Geom




is




  Create (C : Curve from Geom; Offset : Real;  V : Dir)
     returns mutable OffsetCurve
        ---Purpose :
        --  C is the basis curve, Offset is the distance between <me> and
        --  the basis curve at any point. V defines the fixed reference 
        --  direction (offset direction). If P is a point on the basis
        --  curve and T the first derivative with non zero length
        --  at this point, the corresponding point on the offset curve is
        --  in the direction of the vector-product N = V ^ T   where
        --  N is a unitary vector.
        --  Warnings :
        --  In this package the entities are not shared. The OffsetCurve is
        --  built with a copy of the curve C. So when C is modified the
        --  OffsetCurve is not modified
     raises ConstructionError;
        ---Purpose :
        --  Raised if the basis curve C is not at least C1.
        --  Warnings :
        --  No check is done to know if ||V^T|| != 0.0 at any point.
        


  Reverse (me : mutable);
        ---Purpose  : Changes the orientation of this offset curve.
    	-- As a result:
    	-- - the basis curve is reversed,
    	-- - the start point of the initial curve becomes the
    	--   end point of the reversed curve,
    	-- - the end point of the initial curve becomes the
    	--   start point of the reversed curve, and
    	-- - the first and last parameters are recomputed.
  

  ReversedParameter(me; U : Real) returns Real;
	---Purpose: Computes the parameter on the reversed curve for
    	-- the point of parameter U on this offset curve.
 

  SetBasisCurve (me : mutable; C : Curve from Geom)
     raises ConstructionError;
        ---Purpose :  Changes this offset curve by assigning C as the basis curve from which it is built.
    	-- Exceptions
    	-- Standard_ConstructionError if the curve C is not at least "C1" continuous.
      

  SetDirection (me : mutable; V : Dir);
    	---Purpose : Changes this offset curve by assigning V as the
    	-- reference vector used to compute the offset direction.

  SetOffsetValue (me : mutable; D : Real);
        ---Purpose :  Changes this offset curve by assigning D as the offset value.


  BasisCurve (me) returns Curve from Geom;
    	---Purpose : Returns the basis curve of this offset curve.
    	-- Note: The basis curve can be an offset curve.


  Continuity (me)  returns Shape from GeomAbs;
    	---Purpose : Returns the global continuity of this offset curve as a
    	-- value of the GeomAbs_Shape enumeration.
    	-- The degree of continuity of this offset curve is equal
    	-- to the degree of continuity of the basis curve minus 1.
        --  Continuity of the Offset curve :
        --  C0 : only geometric continuity,
        --  C1 : continuity of the first derivative all along the Curve,
        --  C2 : continuity of the second derivative all along the Curve,
        --  C3 : continuity of the third derivative all along the Curve,
        --  G1 : tangency continuity all along the Curve,
        --  G2 : curvature continuity all along the Curve,
        --  CN : the order of continuity is infinite.
        --  Warnings :
        --  Returns the continuity of the basis curve - 1. 
        --  The offset curve must have a unique offset direction defined
        --  at any point.


  Direction (me)  returns Dir;
        ---Purpose : Returns the reference vector of this offset curve.
     	---C++: return const&
   
        ---Purpose  : Value and derivatives
        --  Warnings :
        --  The exception UndefinedValue or UndefinedDerivative is 
        --  raised if it is not possible to compute a unique offset
        --  direction.
        --  If T is the first derivative with not null length and
        --  V the offset direction the relation ||T(U) ^ V|| != 0
        --  must be satisfied to evaluate the offset curve.
        --  No check is done at the creation time and we suppose
        --  in this package that the offset curve is well defined.


  D0(me; U : Real; P : out Pnt);
        ---Purpose:  Warning! this should not be called 
        --          if the basis curve is not at least C1. Nevertheless
        --          if used on portion where the curve is C1, it is OK


  D1 (me; U : Real; P : out Pnt; V1 : out Vec)
     raises UndefinedDerivative;
        ---Purpose:  Warning! this should not be called 
        --           if the continuity of the basis curve is not C2.
        --           Nevertheless, it's OK to use it  on portion 
        --           where the curve is C2


  D2 (me; U : Real; P : out Pnt; V1, V2 : out Vec)
     raises UndefinedDerivative;
        ---Purpose:  Warning! this should not be called 
        --           if the continuity of the basis curve is not C3.
        --           Nevertheless, it's OK to use it  on portion 
        --           where the curve is C3  
       


  D3 (me; U : Real; P : out Pnt; V1, V2, V3 : out Vec)
     raises UndefinedDerivative;
     	---Warning:
        --         this should not be called 
        --           if the continuity of the basis curve is not C4.
        --           Nevertheless, it's OK to use it  on portion 
        --           where the curve is C4  
       

        

  DN (me; U : Real; N : Integer)   returns Vec
        ---Purpose :
        --  The returned vector gives the value of the derivative
        --  for the order of derivation N.    
     	--Warning!
        --         this should not be called 
        --           if the continuity of the basis curve is not CN+1.
        --           Nevertheless, it's OK to use it  on portion 
        --           where the curve is CN+1  
       
     raises UndefinedDerivative,




        ---Purpose  : 
        --  The following functions compute the value and derivatives
        --  on the offset curve and returns the derivatives on the
        --  basis curve too.  
        --  The computation of the value and derivatives on the basis
        --  curve are used to evaluate the offset curve
        --  
        --  Warning:
        --  The exception UndefinedValue or UndefinedDerivative is 
        --  raised if it is not possible to compute a unique offset
        --  direction.
    
    	    RangeError;
        ---Purpose : Raised if N < 1.
        --         

  Value (me; U : Real; P, Pbasis : out Pnt; V1basis : out Vec)
     raises UndefinedValue;

    	---Purpose:  Warning! this should not be called 
        --          if the basis curve is not at least C1. Nevertheless
        --          if used on portion where the curve is C1, it is OK 
  
  D0 (me; U : Real; P, Pbasis : out Pnt; V1basis : out Vec)
     raises UndefinedValue;
     	---Purpose:  Warning! this should not be called 
        --           if the continuity of the basis curve is not C1.
        --           Nevertheless, it's OK to use it  on portion 
        --           where the curve is C1

  

  D1 (me; U : Real; P, Pbasis : out Pnt; V1, V1basis, V2basis : out Vec)
     raises UndefinedDerivative;
        ---Purpose:  Warning! this should not be called 
        --           if the continuity of the basis curve is not C1.
        --           Nevertheless, it's OK to use it  on portion 
        --           where the curve is C1

  D2 (me; U : Real; P, Pbasis : out Pnt;  V1, V2, V1basis, V2basis, 
      V3basis : out Vec)
     raises UndefinedDerivative;

    	---Purpose:  Warning!  this should not be called 
        --           if the continuity of the basis curve is not C3.
        --           Nevertheless, it's OK to use it  on portion 
        --           where the curve is C3  
  FirstParameter (me)  returns Real;

  LastParameter (me)   returns Real;

    	--- Purpose: Returns the value of the first or last parameter of this
    	-- offset curve. The first parameter corresponds to the
    	-- start point of the curve. The last parameter
    	-- corresponds to the end point.
    	-- Note: the first and last parameters of this offset curve
    	-- are also the ones of its basis curve.
    
  Offset (me)          returns Real;
    	---Purpose: Returns the offset value of this offset curve.
    
  IsClosed (me)   returns Boolean;
        ---Purpose : Returns True if the distance between the start point 
        --  and the end point of the curve is lower or equal to 
        --  Resolution from package gp.


  IsCN (me; N : Integer)  returns Boolean
        ---Purpose : Returns true if the degree of continuity of the basis
    	-- curve of this offset curve is at least N + 1.
        --  This method answer True if the continuity of the basis curve 
        --  is N + 1.  We suppose in this class that a normal direction
        --  to the basis curve (used to compute the offset curve) is 
        --  defined at any point on the basis curve.
     raises RangeError;
        ---Purpose : Raised if N < 0.


  IsPeriodic (me)  returns Boolean;
    	---Purpose : Returns true if this offset curve is periodic, i.e. if the
    	-- basis curve of this offset curve is periodic.


  Period (me) returns Real from Standard
	---Purpose: Returns the period of this offset curve, i.e. the period
    	-- of the basis curve of this offset curve.
    	-- Exceptions
    	-- Standard_NoSuchObject if the basis curve is not periodic.
  raises
    	NoSuchObject from Standard
  is redefined;


  Transform (me : mutable; T : Trsf);
        --- Purpose: Applies the transformation T to this offset curve.
    	-- Note: the basis curve is also modified.

  TransformedParameter(me; U : Real; T : Trsf from gp) returns Real
    	---Purpose: Returns the  parameter on the  transformed  curve for
    	--       the transform of the point of parameter U on <me>.
    	--      me->Transformed(T)->Value(me->TransformedParameter(U,T))
	--          is the same point as
	--          me->Value(U).Transformed(T)
	--          This methods calls the basis curve method.
     is redefined;  

  ParametricTransformation(me; T : Trsf from gp) returns Real
    	---Purpose: Returns a  coefficient to compute the parameter on
    	--          the transformed  curve  for  the transform  of the
	--          point on <me>.
	--          
    	--          Transformed(T)->Value(U * ParametricTransformation(T))
	--          is the same point as
	--          Value(U).Transformed(T)
	--          This methods calls the basis curve method.
     is redefined;  

	     

  Copy (me)  returns mutable like me;
    	---Purpose: Creates a new object which is a copy of this offset curve.

fields

  basisCurve  : Curve from Geom;
  direction   : Dir;
  offsetValue : Real;

end;
