-- Created on: 2000-08-15
-- Created by: data exchange team
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



package MXCAFDoc 

	---Purpose: 

uses
    TopLoc,
    PTopLoc,
    TDF,
    PDF,
    MDF,
    MDataStd,
    CDM

is
    class DocumentToolRetrievalDriver;
    class DocumentToolStorageDriver;
    class ColorToolRetrievalDriver;
    class ColorToolStorageDriver;
    class ShapeToolRetrievalDriver;
    class ShapeToolStorageDriver;

    class LayerToolRetrievalDriver;
    class LayerToolStorageDriver;
    
    class LocationStorageDriver;
    class LocationRetrievalDriver;
    class ColorStorageDriver;
    class ColorRetrievalDriver;
    class VolumeStorageDriver;
    class VolumeRetrievalDriver;
    class AreaStorageDriver;
    class AreaRetrievalDriver;
    class CentroidStorageDriver;
    class CentroidRetrievalDriver;
    
    class GraphNodeStorageDriver;
    class GraphNodeRetrievalDriver;

    class DatumStorageDriver;
    class DatumRetrievalDriver;
    class DimTolStorageDriver;
    class DimTolRetrievalDriver;
    class DimTolToolRetrievalDriver;
    class DimTolToolStorageDriver;
    class MaterialStorageDriver;
    class MaterialRetrievalDriver;
    class MaterialToolRetrievalDriver;
    class MaterialToolStorageDriver;

    AddStorageDrivers(aDriverSeq : ASDriverHSequence from MDF; theMsgDriver : MessageDriver from CDM);
	---Purpose: Adds the attribute storage drivers to <aDriverSeq>.


    AddRetrievalDrivers(aDriverSeq : ARDriverHSequence from MDF; theMsgDriver : MessageDriver from CDM);
	---Purpose: Adds the attribute retrieval drivers to <aDriverSeq>.


end MXCAFDoc;
