-- Created on: 1997-11-20
-- Created by: Philippe MANGIN
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



deferred class SectionLaw from GeomFill inherits TShared from MMgt  

	---Purpose: To define section law in  sweeping        

uses 
 BSplineSurface   from Geom,  
 Curve            from Geom, 
 HCurve           from Adaptor3d, 
 Shape            from GeomAbs,
 Pnt              from gp, 
 Array1OfPnt      from TColgp,
 Array1OfVec      from TColgp, 
 Array1OfInteger  from TColStd,
 Array1OfReal     from TColStd  

raises NotImplemented , 
       DomainError,
       OutOfRange from  Standard 
is  
-- 
--========== To compute Sections and derivatives Sections
--      

   D0(me : mutable; 
      Param: Real;
      Poles    : out Array1OfPnt   from TColgp;
      Weigths  : out Array1OfReal  from TColStd)
      ---Purpose: compute the section for v = param           
   returns Boolean  is  deferred;
	
   D1(me : mutable;
      Param: Real;
      Poles    : out Array1OfPnt   from TColgp;
      DPoles   : out Array1OfVec   from TColgp;
      Weigths  : out Array1OfReal  from TColStd;
      DWeigths : out Array1OfReal  from TColStd)
      ---Purpose: compute the first  derivative in v direction  of the
      --           section for v =  param 
      --  Warning : It used only for C1 or C2 aproximation
   returns Boolean  
   raises  NotImplemented 
   is  virtual; 
   
    D2(me : mutable;
      Param: Real;
      Poles     : out Array1OfPnt   from TColgp;
      DPoles    : out Array1OfVec   from TColgp;
      D2Poles   : out Array1OfVec   from TColgp;
      Weigths   : out Array1OfReal  from TColStd;
      DWeigths  : out Array1OfReal  from TColStd;
      D2Weigths : out Array1OfReal  from TColStd)      
      ---Purpose: compute the second derivative  in v direction of the
      --          section  for v = param  
      --  Warning : It used only for C2 aproximation
   returns Boolean 
   raises  NotImplemented  
   is  virtual; 
    
   BSplineSurface(me) 
   ---Purpose: give if possible an bspline Surface, like iso-v are the
   --          section.   If it is  not possible this  methode have to
   --          get an Null Surface. It is the default  implementation.
   returns BSplineSurface  from  Geom
   is  virtual;

    SectionShape(me; NbPoles   : out Integer from Standard;
                     NbKnots   : out Integer from Standard;
                     Degree    : out Integer from Standard) 
	---Purpose: get the format of an  section
    is  deferred;  
    
    Knots(me; TKnots: out Array1OfReal from TColStd)
	---Purpose: get the Knots of the section 
	is deferred;

    Mults(me; TMults: out Array1OfInteger from TColStd)
	---Purpose: get the Multplicities of the section          
	is deferred;   

    IsRational(me)
	---Purpose: Returns if the sections are rationnal or not         
    returns Boolean  is deferred;  
     
    IsUPeriodic(me)  
        ---Purpose: Returns if the sections are periodic or not       
    returns Boolean  is deferred;  
     
    IsVPeriodic(me)  
        ---Purpose: Returns if law is periodic or not       
    returns Boolean  is deferred;  
--
--  =================== Management  of  continuity  ===================
--                 
    NbIntervals(me; S : Shape from GeomAbs) 
	---Purpose: Returns  the number  of  intervals for  continuity
	--          <S>. 
        --          May be one if Continuity(me) >= <S>
   returns Integer  is  deferred;

   Intervals(me; T : in out Array1OfReal from TColStd; 
    	         S : Shape from GeomAbs)
	---Purpose: Stores in <T> the  parameters bounding the intervals
	--          of continuity <S>.
	--          
	--          The array must provide  enough room to  accomodate
	--          for the parameters. i.e. T.Length() > NbIntervals()
    raises
    	OutOfRange from Standard 
    is deferred;  
     
    	
   SetInterval(me: mutable; First, Last: Real from Standard)    
	---Purpose: Sets the bounds of the parametric interval on 
	--          the function
	--          This determines the derivatives in these values if the
	--          function is not Cn.
   is deferred; 
   
   GetInterval(me; First, Last: out Real from Standard)    
	---Purpose: Gets the bounds of the parametric interval on 
	--          the function
   is deferred;  
    
   GetDomain(me; First, Last: out  Real from Standard)  
    	---Purpose: Gets the bounds of the function parametric domain.
    	--  Warning: This domain it is  not modified by the
    	--          SetValue method         
   is  deferred; 
   
--  ===================== To  help  computation  of  Tolerance ======
--      Evaluation of error, in 2d space, or on rational function, is
--      difficult.  The following methods can help the approximation to
--      make good evaluation and use good tolerances.
--      
--       It is not necessary for the following informations to be very
--       precise. A fast evaluation is sufficient.
      
  GetTolerance(me;  
    	       BoundTol, SurfTol, AngleTol : Real;
	       Tol3d : out Array1OfReal)
	---Purpose: Returns the tolerances associated at each poles to
	--          reach  in approximation, to satisfy: BoundTol error
	--          at the   Boundary  AngleTol tangent error  at  the
	--          Boundary  (in radian)  SurfTol   error inside the
	--          surface.
  is  deferred; 
   
  
  SetTolerance(me :  mutable; Tol3d, Tol2d  :  Real) 
  ---Purpose: Is  usefull, if (me)  have to run  numerical
  --          algorithm  to perform D0,  D1 or D2 
  -- The default implementation make nothing.
        
  is virtual; 
   
  BarycentreOfSurf(me) 
   ---Purpose:  Get the barycentre of Surface.   
   --          An   very  poor estimation is sufficent. 
   --          This information is usefull to perform well 
   --          conditioned rational approximation.
   --  Warning: Used only if <me> IsRational         
   returns Pnt from gp    
   raises  NotImplemented   
   is  virtual; 
      
	
   MaximalSection(me) returns Real
    	---Purpose: Returns the   length of the greater section. This
    	--          information is usefull to G1's control.
        --  Warning: With an little value, approximation can be slower.
   is deferred;
    
   GetMinimalWeight(me; Weigths  : out Array1OfReal  from TColStd)
    	---Purpose: Compute the minimal value of weight for each poles
    	--          in all  sections.  
        --          This information is  usefull to control error
    	--          in rational approximation.
        --  Warning: Used only if <me> IsRational        
   raises  NotImplemented   
   is virtual;  
    
--- Particular case  

    IsConstant(me;  Error  :  out  Real)   
	---Purpose: Say if all sections are equals          
    returns  Boolean   
    is  virtual;

    ConstantSection(me)  
     	---Purpose:  Return a  copy of the  constant Section,  if me
     	--          IsConstant
     	--               
    returns  Curve  from  Geom 
    raises  DomainError  --  If  <me>  is  not  Constante
    is  virtual;
  
    IsConicalLaw(me;  Error  :  out  Real) 
    ---Purpose:  Returns True if all section  are circle, with same 
    --          plane,same center and  linear  radius  evolution
    --          Return False by Default.
    returns  Boolean 
    is  virtual;     
     
    CirclSection(me;  Param  :  Real)  
      ---Purpose:  Return the circle section  at parameter <Param>, if
      --          <me> a  IsConicalLaw
    returns  Curve  from  Geom  
    raises  DomainError  --  If  <me>  is  not  a  Conical  Law
    is  virtual;

end SectionLaw;
