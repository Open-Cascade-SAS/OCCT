-- File:	BRepBndLib.cdl
-- Created:	Thu Jul 22 16:12:28 1993
-- Author:	Isabelle GRIGNON
--		<isg@nonox>
---Copyright:	 Matra Datavision 1993


package BRepBndLib 

	---Purpose: This package provides the bounding boxes for curves
	--          and surfaces from BRepAdaptor. 
-- Functions to add a topological shape to a bounding box
uses BRepAdaptor,
     Bnd,
     TopoDS,
     Geom,
     GeomAbs,
     TColgp,
     gp

is

    --
    -- 	 Package methods for shapes
    -- 	 

    Add(S : Shape from TopoDS; B : in out Box from Bnd);
    	---Purpose:Adds the shape S to the bounding box B.
-- More precisely are successively added to B:
-- -   each face of S; the triangulation of the face is used if it exists,
-- -   then each edge of S which does not belong to a face,
--   the polygon of the edge is used if it exists
-- -   and last each vertex of S which does not belong to an edge.
--   After each elementary operation, the bounding box B is
-- enlarged by the tolerance value of the relative sub-shape.
-- When working with the triangulation of a face this value of
-- enlargement is the sum of the triangulation deflection and
-- the face tolerance. When working with the
-- polygon of an edge this value of enlargement is
-- the sum of the polygon deflection and the edge tolerance.
-- Warning
-- -   This algorithm is time consuming if triangulation has not
--   been inserted inside the data structure of the shape S.
-- -   The resulting bounding box may be somewhat larger than the object.
	
	
    AddClose(S : Shape from TopoDS; B : in out Box from Bnd);
    	---Purpose: Adds the shape S to the bounding box B.
-- This is a quick algorithm but only works if the shape S is
-- composed of polygonal planar faces, as is the case if S is
-- an approached polyhedral representation of an exact
-- shape. Pay particular attention to this because this
-- condition is not checked and, if it not respected, an error
-- may occur in the algorithm for which the bounding box is built.
-- Note that the resulting bounding box is not enlarged by the
-- tolerance value of the sub-shapes as is the case with the
-- Add function. So the added part of the resulting bounding
-- box is closer to the shape S.
	
		     
end BRepBndLib;




