-- Created on: 1993-02-10
-- Created by: Mireille MERCIEN
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

generic class HQueue from PCollection (Item as Storable)
inherits Persistent

     ---Purpose: A queue is a sequence of items in which items 
     -- are added at one end (called the back of the
     -- queue) and removed at the other end (called
     -- the front)
     -- The Queue is empty if there are no elements.

raises   NoSuchObject from Standard


    class QueueNode instantiates HSingleList from PCollection(Item);

    class QueueIterator from PCollection 
    	    	    	    	    	   
        ---Purpose: Iterator of the class Queue.

    raises NoMoreObject from Standard,
           NoSuchObject from Standard
    is     
 
     	Create(Q : HQueue from PCollection) 
    	returns QueueIterator from PCollection;
        ---Purpose: Creates an iterator on the queue Q.
        -- Sets the iterator at the beginning of the Queue Q.

     	More(me) returns Boolean from Standard;
        ---Level: Public
        ---Purpose: Returns True if there are other items.

     	Next(me: in out) raises NoMoreObject from Standard;
        ---Level: Public
	---Purpose: Sets the iterator to the next item.
	    
     	Value(me) returns any Item raises NoSuchObject from Standard;
        ---Level: Public
	---Purpose: Returns the item value corresponding to 
	-- the current position of the iterator.

    fields
    	 TheIterator : QueueNode;
    end;


is	
     Create returns mutable HQueue from PCollection;
	---Purpose: Creates an empty queue.

     Length(me) returns Integer from Standard;
        ---Level: Public
	---Purpose: Returns the number of items in the queue.
	---Example: before
	--   me = (A B C) 
	-- returns 3

     IsEmpty(me) returns Boolean from Standard;
        ---Level: Public
	---Purpose: Returns True if the queue contains no element.

     Front(me) returns any Item raises NoSuchObject from Standard; 
        ---Level: Public
	---Purpose: Returns the item at the front of the queue.
	-- Raises an exception if the queue is empty.
        ---Example: before
	--   me = (A B C) 
        -- after
	--   me = (A B C)
       	-- returns 
	--   A
     
     FFront(me) returns QueueNode; 
        ---Level: Public
	---Purpose: Returns the field TheFront(the front of the queue).

     FBack(me) returns QueueNode; 
        ---Level: Public
	---Purpose: Returns the field Theback(the back of the queue).

     Clear(me : mutable);
        ---Level: Public
	---Purpose: Removes all the elements from the queue
	---Example: before
	--   me = (A B C) 
        -- after
        --   me = ()

     Push(me : mutable; T : Item);
        ---Level: Public
	---Purpose: Inserts an item at the back of the queue.
	---Example: before
	--   me = (A B) , T = C
        -- after
	--   me = (A B C)

     Pop(me : mutable) raises NoSuchObject from Standard;
        ---Level: Public
	---Purpose: Removes an item from the front of the queue.
	-- Raises an exception if the queue is empty
	---Example: before
	--   me = (A B C)
        -- after
	--   me = (B C)
	-- returns 
	--   A
 
     ChangeFront(me:mutable ; T : Item) raises NoSuchObject from Standard;
        ---Level: Public
	---Purpose: Replaces the front element of the queue with T.
	-- Raises an exception if the queue is empty.
	---Example: before
	--   me = (A B C) , T = D
        -- after
	--   me = (D B C)

     ShallowCopy(me) 
        returns mutable like me 
        is redefined;
        ---Level: Advanced
	---C++: function call


     ShallowDump (me; s: in out OStream) 
        is redefined;
        ---Level: Advanced
    	---C++: function call


    Destroy(me : mutable);
    ---C++: alias ~
    
fields
     TheFront   : QueueNode;
     TheBack    : QueueNode;
     TheLength  : Integer from Standard;  
end; 






