-- Created on: 1996-03-07
-- Created by: Stagiaire Frederic CALOONE
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Modified:	Wed Mar  5 09:45:42 1997
--    by:	Joelle CHAUVET
--              G1134 : convertion of a GeomPlate_Surface to a Geom_BSplineSurface
--                      by approximation with G0 or G1 criterion
--              + no more reference to TopoDS

package GeomPlate
 
uses gp,
     Adaptor3d,
     Adaptor2d,
     Law,
     GeomFill,
     TColgp,
     Plate,
     Geom,
     math,
     TColGeom,
     TColGeom2d,
     GeomAbs,
     TCollection,
     ElSLib,
     StdFail,   
     ProjLib,
     TColStd,
     AdvApp2Var, 
     Geom2d, 
     Extrema, 
     GeomLProp
     
     
is

    class BuildPlateSurface ; 

    imported Array1OfHCurveOnSurface;     
     
    imported transient class HArray1OfHCurveOnSurface;
     
    class  CurveConstraint; 
     
    class  PointConstraint;  
     
     
    imported Array1OfSequenceOfReal;

    imported transient class HArray1OfSequenceOfReal;

    imported SequenceOfCurveConstraint; 
     
    imported SequenceOfPointConstraint; 
	
    imported transient class HSequenceOfCurveConstraint;
    
    imported transient class HSequenceOfPointConstraint;  


    class BuildAveragePlane;

    class Surface;

    class MakeApprox;

    class PlateG0Criterion;

    class PlateG1Criterion;

    class Aij;

    imported SequenceOfAij;
    
end;






