-- Created on: 1993-05-07
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class WPointInterIterator from TopOpeBRep

uses

    LineInter from TopOpeBRep,
    PLineInter from TopOpeBRep,
    WPointInter from TopOpeBRep
    
is

    -- ==========================
    -- Restriction Point iterator
    -- ==========================

    Create returns WPointInterIterator from TopOpeBRep;
    Create (LI : LineInter from TopOpeBRep) 
    returns WPointInterIterator from TopOpeBRep; 

    Init(me:in out; LI : LineInter from TopOpeBRep) is static;
    Init(me:in out) is static;
    More(me) returns Boolean from Standard is static;
    Next(me:in out) is static;
 
    CurrentWP(me:in out) returns WPointInter from TopOpeBRep 
    ---C++: return const &
    is static;

    PLineInterDummy(me) returns PLineInter from TopOpeBRep;

fields

    myLineInter : PLineInter from TopOpeBRep;
    myWPointIndex : Integer from Standard;
    myWPointNb : Integer from Standard;
    
end WPointInterIterator from TopOpeBRep;
