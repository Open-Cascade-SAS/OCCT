
-- File:	Graphic2d_Paragraph.cdl
-- Created:	Mon Jun 12 16:36:51 1995
-- Author:	Gerard GRAS
--		<gg@azimox>
-- Update:	GG 20/08/98 PERFORMANCE
--		Change Update() method by ComputeMinMax() method 

---Copyright:	 Matra Datavision 1993

class Paragraph from Graphic2d inherits Primitive from Graphic2d

	---Version:

	---Purpose: The primitive Paragraph
	--	    contains a row column of editable texts
	--	    each text can have a different color and font index.

	---Keywords: Primitive, Paragraph, Text
	---Warning:
	---References:

uses
	Drawer				from Graphic2d,
	GraphicObject			from Graphic2d,
	TypeOfAlignment			from Graphic2d,
	PlaneAngle			from Quantity,
	Ratio				from Quantity,
	Factor				from Quantity,
	Length				from Quantity,
	ExtendedString			from TCollection,
	SequenceOfInteger		from TColStd,
	SequenceOfShortReal		from TShort,
	SequenceOfExtendedString	from TColStd,
	CardinalPoints			from Aspect,
	FStream				from Aspect,
	IFStream			from Aspect

raises
	OutOfRange from Standard

is
	-------------------------
	-- Category: Constructors
	-------------------------

	Create (aGraphicObject: GraphicObject from Graphic2d;
		X, Y: Real from Standard;
		anAngle: PlaneAngle from Quantity = 0.0;
		anOffset: CardinalPoints from Aspect = Aspect_CP_Center;
                aScale: Factor from Quantity = 1.0)
	returns mutable Paragraph from Graphic2d;
	---Level: Public
	---Purpose: Creates a paragraph in a graphic object <aGraphicObject>
	--	    The reference point is <X>, <Y>.
	--	    The orientation angle is <anAngle>.
	--	    The offset position of the reference point is <aPosition> 
	--	    depending of the size of paragraph.
	--	    The paragraph scale.
	--	    Angles are measured counterclockwise with 0 radian
	--	    at 3 o'clock.
	--  Warning: a paragraph can be orientable.slantable and zoomable 
	-- only when this options are enable regardless of the graphic driver.
	-- i.e: Xw driver does not,but Xdps or PS driver does.
	---Category: Constructors

	---------------------------------------------------
	-- Category: Methods to modify the class definition
	---------------------------------------------------

	SetSlant (me: mutable; aSlant: PlaneAngle from Quantity = 0.0)
	is static;
	---Level: Public
	---Purpose: Sets the slant angle of the paragraph <me>.
        ---Category: Paragraph management

	SetSpacing(me: mutable; aSpacing: Ratio from Quantity = 0.5)
	is static;
	---Level: Public
	---Purpose: Sets the line spacing ratio for the paragraph <me>.
	--	    the spacing height between two lines depends of
	--	    the spacing factor apply on the height of the line currently	--	    writen.
        ---Category: Paragraph management

	SetMargin(me: mutable; aMargin: Length from Quantity = 0.0)
	is static;
	---Level: Public
	---Purpose: Sets the fixed margin for the paragraph <me>.
        ---Category: Paragraph management

        SetZoomable (me: mutable; aFlag: Boolean from Standard = Standard_False)
        is static;
	---Level: Public
        ---Purpose: The paragraph <me> follows the scale factor of the view
        --          if the flag is Standard_True.
        ---Category: Zoom management


	SetFrameColorIndex (me:mutable; anIndex: Integer from Standard = 0)
	is static;
	---Level: Public
	---Purpose: Sets the frame color index for the paragraph <me>.
        --  Warning: Note that the paragraph frame is drawn only when index 
	--	   is > 0.
        ---Category: Paragraph management

        SetFrameWidthIndex (me:mutable; anIndex: Integer from Standard = 0)
        is static;
        ---Level: Public
        ---Purpose: Sets the width index for the frame of the paragraph <me>.
        --          default width is 0 (1 pixel out line frame is drawn).

	SetHidingColorIndex (me:mutable; anIndex: Integer from Standard = 0)
	is static;
	---Level: Public
	---Purpose: Sets the hiding color index for the paragraph <me>.
        --  Warning: Note that the paragraph background is filled only when index 
	--	is >= 0.
	--	 A value of 0 permits to drawn the paragraph background with
	--	the current view background color.
        ---Category: Paragraph management

	SetCurrentColorIndex (me:mutable; anIndex: Integer from Standard = 1)
	is static;
	---Level: Public
	---Purpose: Sets the current color index for the paragraph <me>.
        --  Warning: Note that the index 0 can be undefined as a ColorMapEntry,
        --        in this case the default color is taken.
        ---Category: Paragraph management

        SetCurrentFontIndex (me:mutable; anIndex: Integer from Standard = 0;
                                aHScale: Length from Quantity = 1.0;
                                aWScale: Length from Quantity = 1.0)
        is static;
        ---Level: Public
        ---Purpose: Sets the current font index and scales for the paragraph <me>.
        --  Warning: Note that the index 0 can be undefined as a FontMapEntry ,
        --         in this case the default system text font is taken.
        ---Category: Paragraph management

	SetCurrentAlignment (me:mutable; anAlignment: TypeOfAlignment from Graphic2d = 
							Graphic2d_TOA_LEFT)
	is static;
	---Level: Public
	---Purpose: Sets the current text alignment for the paragraph <me>.
        ---Category: Paragraph management

	SetCurrentUnderline (me:mutable; isUnderlined: Boolean from Standard =
						Standard_False)
	is static;
	---Level: Public
	---Purpose: Sets the current text underline flag for the paragraph <me>.
        ---Category: Paragraph management

	AddText (me: mutable; aText: ExtendedString from TCollection;
	     		      aRow: Integer from Standard = 0;
	     		      aColumn: Integer from Standard = 0)
        is static;
	---Level: Public
	---Purpose: Adds a text at a row-column position in the paragraph <me>
	-- with the current Color,Font,Alignment attributes
	-- at the position <aColumn,aRow> if <aColumn> and <aRow> are > 0
	--  or at the end of the line if <aColumn> is 0, 
	--  or at the end of the paragraph if <aRow> is 0.
        ---Category: Paragraph management

	ChangeText (me: mutable; aText: ExtendedString from TCollection;
	     		      aRow: Integer from Standard;
	     		      aColumn: Integer from Standard)
        is static;
	---Level: Public
	---Purpose: Changes a text in the paragraph at a row-column position,
	--	    don't change the attributes of the text.
	--  Warning: May do nothing if the row-column don't exist in the
	--	   paragraph.
        ---Category: Paragraph management

        Clear (me: mutable) is static;
        ---Level: Public   
        ---Purpose: Clear ALL the text in the paragraph <me>.
        ---Category: Paragraph management

	--------------------------
	-- Category: Draw and Pick
	--------------------------

	Draw (me : mutable; aDrawer: Drawer from Graphic2d)
	is static protected;
	---Level: Internal
	---Purpose: Draws the paragraph <me>.

	Pick (me : mutable; X, Y: ShortReal from Standard;
		aPrecision: ShortReal from Standard;
		aDrawer: Drawer from Graphic2d)
	returns Boolean from Standard
	is static protected;
	---Level: Internal
	---Purpose: Returns Standard_True if the paragraph <me> is picked,
	--	    Standard_False if not.

    
        ----------------------------
        -- Category: Inquire methods
        ----------------------------
 
        IsZoomable (me)
                returns Boolean from Standard is static;
        ---Level: Internal
        ---Purpose: Returns Standard_True if the Paragraph <me> follows
        --          the scale factor of the view.
        ---Category: Zoom management

        Size (me; aWidth,aHeight: out Length from Quantity) is static;
        ---Level: Public
        ---Purpose: Returns the size of the paragraph <me> .
        ---Category: Paragraph management

        Position (me; X,Y: out Length from Quantity) is static;
        ---Level: Public
        ---Purpose: Returns the paragraph position.

        Offset (me; Dx,Dy: out Length from Quantity) 
	returns CardinalPoints from Aspect is static;
        ---Level: Public
        ---Purpose: Returns the paragraph Offset.

        Angle (me) returns PlaneAngle from Quantity is static;
        ---Level: Public
        ---Purpose: Returns the paragraph orientation.

        Slant (me) returns PlaneAngle from Quantity is static;
        ---Level: Public
        ---Purpose: Returns the paragraph slant.

        Spacing (me) returns Ratio from Quantity is static;
        ---Level: Public
        ---Purpose: Returns the paragraph spacing ratio.

        Margin (me) returns Length from Quantity is static;
        ---Level: Public
        ---Purpose: Returns the paragraph margin value.

        HidingColorIndex (me) returns Integer from Standard is static;
        ---Level: Public
        ---Purpose: Returns the paragraph hiding color index.

        FrameColorIndex (me) returns Integer from Standard is static;
        ---Level: Public
        ---Purpose: Returns the paragraph frame color index.

        FrameWidthIndex (me) returns Integer from Standard is static;
        ---Level: Public
        ---Purpose: Returns the paragraph frame width index.

	    Text( me; aRank: Integer from Standard;
		      aRow,aColumn: out Integer from Standard;
		      aColorIndex,aFontIndex: out Integer from Standard;
		      anAlignment: out TypeOfAlignment from Graphic2d)
        returns ExtendedString from TCollection
	    ---Level: Public
	    ---Purpose: Returns the text string and attributes of rank <aRank>.
	       raises OutOfRange is static;
	    ---Trigger: if aRank is < 1 or > Length().
        ---Category: Paragraph management

        TextSize (me; aRank: Integer from Standard;
	              aWidth,aHeight,anXoffset,anYoffset: out Length from Quantity)
                returns Boolean from Standard
        ---Level: Public
        ---Purpose: Returns Standard_True if the current Driver used is enabled
        --         to get the right size and offsets in the
        --         world size parameter <aWidth>,<aHeight>,<anXoffset>,<anYoffset>
        --         depending of the attributes of the paragraph text position
    	--	    <aRank> and the current scale of the view.
        --          NOTE that the text offsets defines the relative position of the
        --         of the text string origin from the lower left corner of the text
        --         boundary limits.
	       raises OutOfRange is static;
	    ---Trigger: if aRank is < 1 or > Length().
        ---Category: Paragraph management

	    Length (me) returns Integer is static;
	    ---Level: Public
	    ---Purpose: Returns the number of Text of the paragraph <me>.

	    MaxRow (me) returns Integer is static;
	    ---Level: Public
	    ---Purpose: Returns the number of Row of the paragraph <me>.

	    MaxColumn (me) returns Integer is static;
	    ---Level: Public
	    ---Purpose: Returns the number of Column of the paragraph <me>.

        ----------------------------
        -- Category: Private methods
        ----------------------------

        ComputeMinMax (me : mutable)
                returns Boolean from Standard is redefined static;
        ---Level: Internal
        ---Purpose: Computes the MinMax of the paragraph if possible.

	----------------------------------------------------------------------

	Save( me; aFStream: in out FStream from Aspect ) is virtual;
--	Retrieve( me; aIFStream: in out IFStream from AIS2D ) is virtual;

fields

	myX:		ShortReal from Standard;
	myY:		ShortReal from Standard;
	myXoffset:	ShortReal from Standard;
	myYoffset:	ShortReal from Standard;
	myOffset:	CardinalPoints from Aspect;
	myWidth:	ShortReal from Standard;
	myHeight:	ShortReal from Standard;
	myAngle:	ShortReal from Standard;
	mySlant:	ShortReal from Standard;
	mySpacing:	ShortReal from Standard;
	myMargin:	ShortReal from Standard;
	myScale:	ShortReal from Standard;
    myIsZoomable:           Boolean from Standard;
	myFrameColorIndex:	    Integer from Standard;
	myFrameWidthIndex:	    Integer from Standard;
	myHidingColorIndex:	    Integer from Standard;
	myCurrentColorIndex:	Integer from Standard;
	myCurrentFontIndex:	    Integer from Standard;
    myCurrentFontHScale:    ShortReal from Standard;
    myCurrentFontWScale:    ShortReal from Standard;
	myCurrentAlignment:	    TypeOfAlignment from Graphic2d;
	myCurrentUnderline:	    Boolean from Standard;
	myTextStringList:	    SequenceOfExtendedString from TColStd;
	myTextDescriptorList:	SequenceOfInteger from TColStd;
	myTextXpositionList:	SequenceOfShortReal from TShort;
	myTextYpositionList:	SequenceOfShortReal from TShort;
	myTextFheightList:	    SequenceOfShortReal from TShort;
	myTextFoffsetList:	    SequenceOfShortReal from TShort;
    myTextHScaleList:       SequenceOfShortReal from TShort;
    myTextWScaleList:       SequenceOfShortReal from TShort;

end Paragraph from Graphic2d;
