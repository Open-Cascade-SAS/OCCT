-- Created on: 1992-04-07
-- Created by: Christian CAILLET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



deferred class ViewKindEntity  from IGESData  inherits IGESEntity

    ---Purpose : defines required type for ViewKind in directory part
    --           that is, Single view or Multiple view
    --           An effective ViewKind entity must inherit it and define
    --           IsSingle (True for Single, False for List of Views),
    --           NbViews and ViewItem (especially for a List)

uses Boolean

raises OutOfRange

is

    IsSingle (me) returns Boolean  is deferred;
    ---Purpose : says if "me" is a Single View (True) or a List of Views (False)

    NbViews (me) returns Integer  is deferred;
    ---Purpose : Returns the count of Views for a List of Views. For a Single
    --           View, may return simply 1

    ViewItem (me; num : Integer) returns ViewKindEntity
    raises OutOfRange  is deferred;
    ---Purpose : Returns the View n0. <num> for a List of Views. For a Single
    --           Views, may return <me> itself

end ViewKindEntity;
