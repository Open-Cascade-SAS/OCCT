-- Created on: 1997-04-23
-- Created by: Alexander BRIVIN
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PointAspect from VrmlConverter inherits TShared from MMgt

	---Purpose: qualifies the aspect properties for  
	--          the VRML conversation of points. 

uses 

    Material    from   Vrml

is

    Create
    returns mutable PointAspect from VrmlConverter;

    ---Purpose: create a default PointAspect. 
    --  Default value: HasMaterial  =  False  - a  line  hasn't  own  material (color) 

    Create  (aMaterial: Material from Vrml; 
    	    	 OnOff: Boolean from Standard)
    returns mutable PointAspect from VrmlConverter;
 
    SetMaterial(me: mutable; aMaterial: Material from Vrml)
    is static;
 
    Material(me) returns mutable Material from Vrml 
    is  static; 

    SetHasMaterial(me: mutable; OnOff: Boolean from Standard)
    ---Purpose: defines the necessary of writing  own  Material from Vrml into  output  OStream. 
    --          By default False  -  the material is not writing into OStream, 
    --          True  -  the material is writing. 
    is  static; 

    HasMaterial(me) returns Boolean from Standard 
    ---Purpose: returns True if the  materials is  writing into OStream.
    is static;
 
    
fields
     
    myMaterial		:	Material    from   Vrml;    
    myHasMaterial       :       Boolean  from  Standard;
    
end PointAspect;
