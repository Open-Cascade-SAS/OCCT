-- Created on: 1993-04-06
-- Created by: Philippe DAUTRY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Direction from PGeom2d inherits Vector from PGeom2d

        ---Purpose :  The class Direction  specifies a vector that  is
        --         never null. It is a unit vector.
        --         
	---See Also : Direction from Geom2d.

uses  Vec2d from gp

is


  Create returns mutable Direction from PGeom2d;
        --- Purpose : Creates a unit vector with default values.
	---Level: Internal 


  Create (aVec: Vec2d from gp) returns mutable Direction from PGeom2d;
        ---Purpose : Create a unit vector with <aVec>.
	---Level: Internal 


end;
