-- Created on: 1993-03-23
-- Created by: BBL
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class XAlienImage from AlienImage inherits AlienUserImage from AlienImage

    	---Purpose: Defines an X11 Alien image, i.e. an image file to be
    	-- used with X11 xwd utility.

uses
	File 			from OSD,
	AsciiString 		from TCollection,
	ColorImage 		from Image,
	PseudoColorImage 	from Image,
	Image			from Image,
	X11XWDAlienData 	from AlienImage

is
	Create returns mutable XAlienImage from AlienImage;
    	---Purpose: Constructs an empty X11 alien image.
	Clear( me : in out mutable) ;
	---Level: Public
	---Purpose: Frees memory allocated by XAlienImage
	---C++: alias ~

	SetName( me : in out mutable;
		 aName : in AsciiString from TCollection) ;
	---Purpose: Sets the Image name for the Name function.

	Name( me : in immutable ) returns AsciiString from TCollection ;
	---C++: return const &
        ---Purpose: Returns the Image name.

	ToImage( me : in immutable ) 
	  returns mutable Image from Image ;
	---Level: Public
	---Purpose : Converts an XAlienImage object to a Image object.

	FromImage( me : in out mutable ; anImage : in Image from Image ) ;
	---Level: Public
	---Purpose : Converts an Image object to a XAlienImage object.

	Read ( me : in out mutable; afile : in out File from OSD )
	  returns Boolean from Standard ;
	---Level: Public
	---Purpose: Reads the content of a  XAlienImage object from a file .
	--          Returns True if file is a XWD file .

	Write( me : in immutable; afile : in out File from OSD )
	  returns Boolean from Standard ;
	---Level: Public
	---Purpose: Writes the content of a  XAlienImage object to a file .

fields
	myData : X11XWDAlienData  from  AlienImage;

end ;
 
