-- Created on: 1996-01-11
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class WiresOnShape from LocOpe inherits ProjectedWires from LocOpe

	---Purpose: 

uses Shape               from TopoDS,
     Face                from TopoDS,
     Wire                from TopoDS,
     Compound            from TopoDS,
     Edge                from TopoDS,
     Vertex              from TopoDS,
     DataMapOfShapeShape from TopTools,
--     DataMapIteratorOfDataMapOfShapeShape from TopTools
     IndexedDataMapOfShapeShape from TopTools,
     MapOfShape          from TopTools


is

    Create(S: Shape from TopoDS)

    	returns mutable WiresOnShape from LocOpe;


    Init(me: mutable; S: Shape from TopoDS)
    
    	is static;

    SetCheckInterior(me: mutable; ToCheckInterior: Boolean from Standard)
	---Purpose: Set the flag of check internal intersections
	--          default value is True (to check)
	---C++: inline      
    	is static;

    Bind(me: mutable; W: Wire from TopoDS;
                      F: Face from TopoDS)
		     
	is static;

    Bind(me: mutable; Comp: Compound from TopoDS;
                      F:    Face from TopoDS)
		     
	is static;

    Bind(me: mutable; E: Edge from TopoDS;
                      F: Face from TopoDS)
		      
    	is static;


    Bind(me: mutable; EfromW: Edge from TopoDS;
    	              EonFace: Edge from TopoDS)
		      
	is static;


    BindAll(me: mutable)
    
    	is static;


    IsDone(me)
    
    	returns Boolean from Standard
	---C++: inline
	is static;


    InitEdgeIterator(me: mutable)
    
    	;


    MoreEdge(me: mutable)
    	returns Boolean from Standard
	;


    Edge(me: mutable)
    	returns Edge from TopoDS
	;


    OnFace(me: mutable)
	---Purpose: Returns the face of the shape on which the current
	--          edge is projected.
    	returns Face from TopoDS
	;

    
    OnEdge(me: mutable; E: out Edge from TopoDS)
	---Purpose: If the   current  edge is  projected  on  an edge,
	--          returns <Standard_True> and sets the value of <E>.
	--          Otherwise, returns <Standard_False>.
    	returns Boolean from Standard
	;


    NextEdge(me: mutable)
    
    	;


    OnVertex(me: mutable; Vwire :     Vertex from TopoDS;
    	                  Vshape: out Vertex from TopoDS)
			  
	returns Boolean from Standard
	;


    OnEdge(me: mutable; V: Vertex from TopoDS;
                        E: out Edge from TopoDS;
			P: out Real from Standard)
	---Purpose: If the vertex <V> lies on  an edge of the original
	--          shape,  returns     <Standard_True> and   sets the
	--          concerned edge in  <E>,  and the parameter on  the
	--          edge in <P>.
	--          Else returns <Standard_False>.
	returns Boolean from Standard
	;
	
    IsFaceWithSection(me; aFace : Shape from TopoDS)
	---Purpose: tells is the face to be split by section or not
	---C++: inline
	returns Boolean from Standard
	;


fields

    myShape : Shape                      from TopoDS;
    myMapEF : IndexedDataMapOfShapeShape from TopTools;
    myFacesWithSection : MapOfShape      from TopTools;
    myCheckInterior : Boolean            from Standard;
    myMap   : DataMapOfShapeShape        from TopTools;
    myDone  : Boolean                    from Standard;
    myIndex : Integer                    from Standard;

end WiresOnShape;
