-- Created on: 1999-07-29
-- Created by: Roman LYGIN
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package Message 

    	---Purpose: Defines
   	--          - tools to work with messages
    	--          - basic tools intended for progress indication

uses

    MMgt,
    TColStd,
    TCollection,
    Standard

is

    enumeration Gravity is
    	---Purpose: Defines gravity level of messages
	-- - Trace: low-level details on algorithm execution (usually for debug purposes)
	-- - Info: informative message
	-- - Warning: warning message
	-- - Alarm: non-critical error
	-- - Fail: fatal error 
	Trace,
        Info,
        Warning,
        Alarm,
	Fail
    end Gravity;

    imported Status;
    imported StatusType;
    imported ExecStatus;

    class Msg;
    	---Purpose: Defines message.
    class MsgFile;
    	---Purpose: Defines file storing messages.
	
    class Messenger;
    	---Purpose: Messenger is API class providing general-purpose interface for 
	--          libraries that may issue text messages without knowledge
	--          of how these messages will be further processed.
	
    class Algorithm;
	---Purpose: Class Message_Algorithm is the root class for all algorithms.
	--          It provides generic mechanism for management execution status,
	--          collection and output of corresponding error/warning messages

    deferred class Printer;
    	---Purpose: Defines basic message printer.
	
	class PrinterOStream;
	    ---Purpose: Defines printer associated with an ostream
    
    class ListOfMsg instantiates List from TCollection (Msg from Message);
    
    class SequenceOfPrinters instantiates 
    Sequence from TCollection (Printer from Message);

    -- Progress indication
    deferred class ProgressIndicator;
    class ProgressScale;
    class ProgressSentry;
    class SequenceOfProgressScale instantiates
         Sequence from TCollection (ProgressScale from Message);
    
    DefaultMessenger returns Messenger from Message;
        ---Purpose: Defines default messenger for OCCT applications.
        --          This is global static instance of the messenger.
	--          By default, it contains single printer directed to cout.
	--          It can be customized according to the application needs.
	---C++: return const &

    FillTime (Hour, Minute: Integer; Second: Real) returns AsciiString from TCollection;
    	---Purpose: Returns the string filled with values of hours, minutes and seconds.
	-- Example:
    	--          1. (5, 12, 26.3345) returns "05h:12m:26.33s",
	--          2. (0,  6, 34.496 ) returns "06m:34.50s",
	--          3. (0,  0,  4.5   ) returns "4.50s"

end Message;
