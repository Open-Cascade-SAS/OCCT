-- Created on: 1993-03-23
-- Created by: BBL,JLF
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class MemoryOperations from AlienImage

	---Version: 0.0

	---Level: Public
	---Purpose: This class defines class method for
	--          memory mangement .
	---Keywords:
	---Warning:
	---References:
--uses

raises
      NullObject

is
   SwapLong ( myclass ; Data : in Address from Standard
		      ; Size : in Integer from Standard ) 
	---Level: Internal
   ---Purpose: Swap byte in a long word ( 32 Bit )
   --	       Size is the number of long word to swap
   --          ex : SwapLong( "abcd". 1 ) gives "dcba"  
   --          
	raises NullObject;

   SwapShort( myclass ; Data : in Address from Standard
		      ; Size : in Integer from Standard )
	---Level: Internal
   ---Purpose: Swap byte in a short word ( 16 Bit )
   --	       Size is the number of short word to swap
   --          ex : SwapShort( "ab". 1 ) gives "ba"  
   --          
	raises NullObject;

end MemoryOperations;
 
