-- Created on: 1997-11-05
-- Created by: Francois PONTET
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Document from PDocStd inherits Document from PCDM

	---Purpose: 

uses

      Data from PDF

is

    Create
    returns Document from PDocStd;   

    Create (data : Data from PDF)
    returns Document from PDocStd;


    SetData (me : mutable; data : Data from PDF);

    GetData (me) 
    returns Data from PDF;

fields

     myData :  Data from PDF;

end Document;
