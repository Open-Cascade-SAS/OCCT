-- Created on: 2000-01-28
-- Created by: data exchange team
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MsgRegistrator from ShapeExtend inherits BasicMsgRegistrator from ShapeExtend

    ---Purpose: Attaches messages to the objects (generic Transient or shape).
    --          The objects of this class are transmitted to the Shape Healing
    --          algorithms so that they could collect messages occurred during
    --          processing.
    --
    --          Messages are added to the Maps (stored as a field) that can be
    --          used, for instance, by Data Exchange processors to attach those
    --          messages to initial file entities.

uses

    Shape                       from TopoDS,
    Gravity                     from Message,
    Msg                         from Message,
    ListOfMsg                   from Message,
    DataMapOfTransientListOfMsg from ShapeExtend,
    DataMapOfShapeListOfMsg     from ShapeExtend

is

    Create returns MsgRegistrator from ShapeExtend;
    	---Purpose: Creates an object.
	
    
    Send (me: mutable; object : Transient;
    	    	       message: Msg from Message;
    	    	       gravity: Gravity from Message) is redefined;
    	---Purpose: Sends a message to be attached to the object.
	--          If the object is in the map then the message is added to the
    	--          list, otherwise the object is firstly added to the map.

    Send (me: mutable; shape  : Shape from TopoDS;
    	    	       message: Msg from Message;
    	    	       gravity: Gravity from Message) is redefined;
    	---Purpose: Sends a message to be attached to the shape.
	--          If the shape is in the map then the message is added to the
    	--          list, otherwise the shape is firstly added to the map.

    MapTransient (me) returns DataMapOfTransientListOfMsg from ShapeExtend;
    	---C++    : inline
    	---C++    : return const&
	---Purpose: Returns a Map of objects and message list
	
    MapShape (me) returns DataMapOfShapeListOfMsg from ShapeExtend;
    	---C++    : inline
    	---C++    : return const&
	---Purpose: Returns a Map of shapes and message list

fields

    myMapTransient: DataMapOfTransientListOfMsg from ShapeExtend;
    myMapShape: DataMapOfShapeListOfMsg from ShapeExtend;
    
end MsgRegistrator;
