-- Created on: 2000-05-18
-- Created by: Peter KURNEV
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.
 
package BOPTest 
---Purpose: 

uses
    gp,
    Draw,
    DBRep, 
    TopAbs,    	     
    TopoDS,
    TopTools, 
    BOPCol,    
    BOPDS,    
    BOPAlgo 
     
is  
    
    class Objects; 
    class DrawableShape; 
    -- 
    AllCommands        (aDI:out Interpretor from Draw);
    BOPCommands        (aDI:out Interpretor from Draw); 
    CheckCommands      (aDI:out Interpretor from Draw); 
    TolerCommands      (aDI:out Interpretor from Draw); 
    LowCommands        (aDI:out Interpretor from Draw); 
    ObjCommands        (aDI:out Interpretor from Draw);
    PartitionCommands  (aDI:out Interpretor from Draw);
    APICommands        (aDI:out Interpretor from Draw); 
    OptionCommands     (aDI:out Interpretor from Draw); 
    HistoryCommands    (aDI:out Interpretor from Draw); 

    Factory            (aDI:out Interpretor from Draw);
    
end BOPTest;
