-- Created on: 2000-02-07
-- Created by: data exchange team
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package ShapeAlgo 

    ---Purpose: 

uses

    MMgt,
    Geom,
    Geom2d,
    TColGeom,
    TColGeom2d,
    TopoDS,
    ShapeExtend,
    ShapeAnalysis,
    ShapeFix,
    GeomAbs

is

    class ToolContainer;

    class AlgoContainer;
    	---Purpose: Provides initerface to the algorithms from Shape Healing.

    Init;
    	---Purpose: Creates and initializes default AlgoContainer.
    
    SetAlgoContainer (aContainer: AlgoContainer from ShapeAlgo);
    	---Purpose: Sets default AlgoContainer

    AlgoContainer returns AlgoContainer from ShapeAlgo;
    	---Purpose: Returns default AlgoContainer

end ShapeAlgo;
