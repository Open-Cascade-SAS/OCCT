-- File:	BRepBlend_SurfRstConstRad.cdl
-- Created:	Thu Feb  6 16:22:22 1997
-- Author:	Jacques GOUSSARD
-- Author:	Laurent BOURESCHE
--		<lbo@pomalox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1997

class SurfRstConstRad from BRepBlend
inherits SurfRstFunction from Blend


uses Vector          from math,
     Matrix          from math,
     Ax1             from gp,
     Vec             from gp,
     Vec2d           from gp,
     Pnt             from gp,
     Pnt2d           from gp,
     Circ            from gp,
     Array1OfPnt     from TColgp,
     Array1OfVec     from TColgp,
     Array1OfPnt2d   from TColgp,
     Array1OfVec2d   from TColgp,
     Array1OfReal    from TColStd,
     Array1OfInteger from TColStd,
     Shape           from GeomAbs,
     Point           from Blend,
     SectionShape    from BlendFunc,
     HSurface        from Adaptor3d,
     HCurve          from Adaptor3d,
     HCurve2d        from Adaptor2d,
     CurveOnSurface  from Adaptor3d,
     ParameterisationType from Convert


is

    Create(Surf    : HSurface from Adaptor3d;
    	   SurfRst : HSurface from Adaptor3d;
    	   Rst     : HCurve2d from Adaptor2d; 
    	   CGuide  : HCurve   from Adaptor3d)
    returns SurfRstConstRad from BRepBlend;

    NbVariables(me)
    ---Purpose: Returns 3.
    returns Integer from Standard;

    NbEquations(me)
    ---Purpose: Returns 3.
    returns Integer from Standard;

    Value(me: in out; X: Vector; F: out Vector)
    ---Purpose: computes the values <F> of the Functions for the 
    --          variable <X>.
    --          Returns True if the computation was done successfully, 
    --          False otherwise.
    returns Boolean from Standard;
    
    Derivatives(me: in out; X: Vector; D: out Matrix)
    ---Purpose: returns the values <D> of the derivatives for the 
    --          variable <X>.
    --          Returns True if the computation was done successfully, 
    --          False otherwise.
    returns Boolean from Standard;
    
    Values(me: in out; X: Vector; F: out Vector; D: out Matrix)
    ---Purpose: returns the values <F> of the functions and the derivatives
    --          <D> for the variable <X>.
    --          Returns True if the computation was done successfully, 
    --          False otherwise.
    returns Boolean from Standard;

    Set(me      : in out; 
        SurfRef : HSurface from Adaptor3d;
    	RstRef  : HCurve2d from Adaptor2d);
    	   
    Set(me: in out; Param: Real from Standard);

    Set(me: in out; First, Last: Real from Standard);
    ---Purpose: Sets the bounds of the parametric interval on 
    --          the guide line.
    --          This determines the derivatives in these values if the
    --          function is not Cn.

    GetTolerance(me; Tolerance: out Vector from math; Tol: Real from Standard);

    GetBounds(me; InfBound,SupBound: out Vector from math);

    IsSolution(me: in out; Sol: Vector from math; Tol: Real from Standard)
    returns Boolean from Standard;

     GetMinimalDistance(me) 
        ---Purpose: Returns   the    minimal  Distance  beetween   two
        --          extremitys of calculed sections.          
   	returns  Real  from  Standard 
	is redefined;

--- TheFollowing methods are called only when 
--  IsSolution returns Standard_True.

    PointOnS(me)
    ---C++: return const&
    returns Pnt from gp;

    PointOnRst(me)
    ---C++: return const&
    returns Pnt from gp;

    Pnt2dOnS(me)
    ---Purpose: Returns U,V coordinates of the point on the surface.
    ---C++: return const&
    returns Pnt2d from gp;

    Pnt2dOnRst(me)
    ---Purpose: Returns  U,V coordinates of the point  on the curve on
    --          surface.
    ---C++: return const&
    returns Pnt2d from gp;

    ParameterOnRst(me)
    ---Purpose: Returns parameter of the point on the curve.
    returns Real from Standard;

    IsTangencyPoint(me)
    returns Boolean from Standard;

    TangentOnS(me)
    ---C++: return const&
    returns Vec from gp;

    Tangent2dOnS(me)
    ---C++: return const&
    returns Vec2d from gp;

    TangentOnRst(me)
    ---C++: return const&
    returns Vec from gp;

    Tangent2dOnRst(me)
    ---C++: return const&
    returns Vec2d from gp;

    Decroch(me; 
    	    Sol    : Vector from math;
    	    NS,TgS : out Vec from gp)
    ---Purpose: Enables  implementation  of  a criterion of  decrochage
    --          specific to  the function. 
    --  Warning: Can  be  called  without  previous  call  of  issolution
    --          but the values  calculated can  be  senseless.    
    returns Boolean from Standard
    is static;

-- methodes hors template (en plus du create)

    Set(me     : in out; 
    	Radius : Real from Standard; 
    	Choix  : Integer from Standard)
    is static;

    Set(me: in out; TypeSection: SectionShape from BlendFunc)
    ---Purpose: Sets  the  type  of   section generation   for the
    --          approximations. 
    is static;

    Section(me        : in out; 
            Param     : Real from Standard;
            U,V,W     : Real from Standard;
            Pdeb,Pfin : out Real from Standard;
            C         : out Circ from gp)
    is static;

-- Methods for the approximation
-- 
    IsRational(me) returns Boolean
    ---Purpose: Returns  if the section is rationnal
    is static;

    GetSectionSize(me) returns Real
    ---Purpose:  Returns the length of the maximum section
    is static;
    
    GetMinimalWeight(me; Weigths  : out Array1OfReal  from TColStd)
    ---Purpose: Compute the minimal value of weight for each poles
    --          of all sections.
    is static;

    NbIntervals(me; S : Shape from GeomAbs) returns Integer
    ---Purpose: Returns  the number  of  intervals for  continuity
    --          <S>. May be one if Continuity(me) >= <S>
    is static;
    
    Intervals(me; T : in out Array1OfReal from TColStd; 
    	          S : Shape from GeomAbs)
    ---Purpose: Stores in <T> the  parameters bounding the intervals
    --          of continuity <S>.        
    --          The array must provide  enough room to  accomodate
    --          for the parameters. i.e. T.Length() > NbIntervals()
    is static;

    GetShape(me        : in out;
             NbPoles   : out Integer from Standard;
    	     NbKnots   : out Integer from Standard;
             Degree    : out Integer from Standard;
             NbPoles2d : out Integer from Standard)
    is static;

    GetTolerance(me; 
    	    	 BoundTol, SurfTol, AngleTol : Real;
		 Tol3d : out Vector;
		 Tol1D : out Vector )
    ---Purpose: Returns the tolerance to reach in approximation
    --          to respecte
    --          BoundTol error at the Boundary
    --          AngleTol tangent error at the Boundary
    --          SurfTol error inside the surface.
    is static;

    Knots(me: in out; TKnots: out Array1OfReal from TColStd)
    is static;

    Mults(me: in out; TMults: out Array1OfInteger from TColStd)
    is static;

    Section(me       : in out ; 
    	    P        : Point from Blend;
            Poles    : out Array1OfPnt   from TColgp;
	    DPoles   : out Array1OfVec   from TColgp;
  	    Poles2d  : out Array1OfPnt2d from TColgp;
	    DPoles2d : out Array1OfVec2d from TColgp;
	    Weigths  : out Array1OfReal  from TColStd;
	    DWeigths : out Array1OfReal  from TColStd)
    ---Purpose: Used for the first and last section 
    returns Boolean from Standard
    is static;

    Section(me: in out; P: Point from Blend;
			Poles     : out Array1OfPnt   from TColgp;
			DPoles    : out Array1OfVec   from TColgp;
			D2Poles   : out Array1OfVec   from TColgp;
    	                Poles2d   : out Array1OfPnt2d from TColgp;
			DPoles2d  : out Array1OfVec2d from TColgp;
			D2Poles2d : out Array1OfVec2d from TColgp;
			Weigths   : out Array1OfReal  from TColStd;
			DWeigths  : out Array1OfReal  from TColStd;
                        D2Weigths : out Array1OfReal  from TColStd)
    ---Purpose: Used for the first and last section
    --          The method returns Standard_True if the derivatives
    --          are computed, otherwise it returns Standard_False.
    returns Boolean from Standard
    is static;

    Section(me       : in out ; 
    	    P        : Point from Blend;
            Poles    : out Array1OfPnt   from TColgp;
    	    Poles2d  : out Array1OfPnt2d from TColgp;
	    Weigths  : out Array1OfReal  from TColStd)
    is static;

    Resolution(me; 
    	       IC2d : Integer from Standard;
	       Tol  : Real from Standard;
	       TolU, TolV : out Real from Standard);

fields

    surf     : HSurface             from Adaptor3d;
    surfrst  : HSurface             from Adaptor3d;
    rst      : HCurve2d             from Adaptor2d;
    cons     : CurveOnSurface       from Adaptor3d;
    guide    : HCurve               from Adaptor3d; 
    tguide   : HCurve               from Adaptor3d; 
    pts      : Pnt                  from gp;
    ptrst    : Pnt                  from gp;
    pt2ds    : Pnt2d                from gp;
    pt2drst  : Pnt2d                from gp;
    prmrst   : Real                 from Standard;
    istangent: Boolean              from Standard;
    tgs      : Vec                  from gp;
    tg2ds    : Vec2d                from gp;
    tgrst    : Vec                  from gp;
    tg2drst  : Vec2d                from gp;

    ray      : Real                 from Standard;
    choix    : Integer              from Standard;
    ptgui    : Pnt                  from gp;
    d1gui    : Vec                  from gp;
    d2gui    : Vec                  from gp;
    nplan    : Vec                  from gp;
    normtg   : Real                 from Standard;
    theD     : Real                 from Standard;
       
    surfref  : HSurface             from Adaptor3d;
    rstref   : HCurve2d             from Adaptor2d;

    maxang   : Real                 from Standard;
    minang   : Real                 from Standard;   
    distmin  : Real                 from Standard;   
    mySShape : SectionShape         from BlendFunc;
    myTConv  : ParameterisationType from Convert;

end SurfRstConstRad;
