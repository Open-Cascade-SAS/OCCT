-- Created on: 1999-03-09
-- Created by: data exchange team
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PersonAndOrganizationItem from StepAP214 inherits ApprovalItem from StepAP214

	-- <PersonAndOrganizationItem> is an EXPRESS Select Type construct translation.
	-- it gathers : ApprovalPersonOrganization, AutoDesignDateAndPersonAssignment

uses

    	AppliedOrganizationAssignment from StepAP214
	
is

	Create returns PersonAndOrganizationItem;
	---Purpose : Returns a PersonAndOrganizationItem SelectType

	CaseNum (me; ent : Transient) returns Integer is redefined;
	---Purpose: Recognizes a APersonAndOrganizationItem Kind Entity that is :
    	--        1 -> AppliedOrganizationAssignment
    	--        2 -> AssemblyComponentUsageSubstitute
	--        3 -> DocumentFile
    	--        4 -> MaterialDesignation
    	--        5 -> MechanicalDesignGeometricPresentationRepresentation
	--        6 -> PresentationArea
    	--        7 -> Product
	--        8 -> ProductDefinition
    	--        9 -> ProductDefinitionFormation
	--    	  10 -> ProductDefinitionRelationship
	--        11 -> PropertyDefinition
    	--        12 -> ShapeRepresentation
    	--        13 -> SecurityClassification
	--        0 else


    	AppliedOrganizationAssignment (me) returns any AppliedOrganizationAssignment;
    	---Purpose : returns Value as a AppliedOrganizationAssignment (Null if another type)

	
end PersonAndOrganizationItem;
