-- File:	MeshDS_Node.cdl
-- Created:	Thu Sep  9 18:28:16 1993
-- Author:	Didier PIFFAULT
--		<dpf@zerox>
---Copyright:	 Matra Datavision 1993


deferred generic class Node from MeshDS (dummyarg as any)

	---Purpose: Describes the  necessary services of a node to use
	---         it in a Mesh data structure.

uses DegreeOfFreedom from MeshDS

is      Movability     (me)
    	    returns DegreeOfFreedom from MeshDS;


    	SetMovability  (me: in out; canMove : DegreeOfFreedom from MeshDS);


    	Domain         (me)
    	    returns Integer from Standard;


---Purpose: For maping the Nodes.
--          Same Node -> Same HashCode
--          Different Nodes -> Not IsEqual but can have same HashCode 

	HashCode       (me;
    	    	    	Upper : Integer from Standard)
	---C++: function call
	    returns Integer from Standard;


	IsEqual        (me; Other : Node from MeshDS)
	---C++: alias operator ==
	    returns Boolean from Standard;

end Node;
