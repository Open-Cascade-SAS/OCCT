-- File:	IGESSolid_ToolBooleanTree.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolBooleanTree  from IGESSolid

    ---Purpose : Tool to work on a BooleanTree. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses BooleanTree from IGESSolid,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolBooleanTree;
    ---Purpose : Returns a ToolBooleanTree, ready to work


    ReadOwnParams (me; ent : mutable BooleanTree;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : BooleanTree;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : BooleanTree;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a BooleanTree <ent>, from
    --           its specific (own) parameters

    DirChecker (me; ent : BooleanTree) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : BooleanTree;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : BooleanTree; entto : mutable BooleanTree;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : BooleanTree;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolBooleanTree;
