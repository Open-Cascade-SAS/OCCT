-- Created on: 2001-05-03
-- Created by: Igor FEOKTISTOV
-- Copyright (c) 2001-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

package QANewModTopOpe 

    	---Purpose:  QANewModTopOpe  package  provides  classes  for  limitation, gluing 
	--           and removing "floating" shapes.
uses 
  
    BRepAlgoAPI,
    TopoDS, 
    TopTools, 
    TopAbs,
    BRepTools, 
    gp,
    BOPAlgo, 
    BOPDS
 
is 
  
    enumeration  ModeOfLimitation  is  Forward,   
    	    	                       Reversed, 
				       BothParts;  
				       
    pointer  CutPtr  to  Cut  from  BRepAlgoAPI;
    pointer  CommonPtr  to  Common  from  BRepAlgoAPI;
				       
    class Tools; 
        ---Purpose: to  provide  several  tools  for  porting  to  OCC  5.0  (mkk)

    class  Limitation;  
    	---Purpose: to  provide  cutting  object  by  face  or  shell. 

    class  Intersection;  
    	---Purpose: to  provide  intersection  of  two  topological  objects.  
	 
    class Glue;                     ---  inherits BooleanOperation from BRepAlgoAPI
    	---Purpose: to  provide  topological  sewing  of  two  topological  objects.  

    class ReShaper;
    	---Purpose: to remove  "floating" objects from compound.
	-- "floating" objects are wires, edges, vertices that do not belong
	-- solids, shells or faces.
     
    IsValid(TheS : Shape  from  TopoDS; GeomControls : Boolean from Standard =  Standard_True)
    	returns Boolean from Standard;
    	---Purpose: to check if TheS is valid or not. 
	-- in difference with BRepCheck_Analizer, this method allows 
	-- some  kind of  non-manifold shapes 
	
    IsManifold(TheS : Shape  from  TopoDS) returns Boolean from Standard;
    	---Purpose: to check if TheS is manifol or not.
	-- manifold shape is valid SOLID, SHELL, WIRE, EDGE, VERTEX without internal 
	-- subshapes - faces, wires, edges and vertices that have INTERNAL orientation
	-- For SHELL there are additional conditions: orientations of faces must 
	-- corresponds each other, each edge must be shared not more then two faces.
	-- COMPSOLID is non manifold by default.
	-- COMPOUND conciders to  be manifold if:
	-- 1) all shapes in compound are manifold (see above mentioned definitions)
	-- 2) all shapes are fully disconnected - there are any shapes in  compound that 
	--    share common subshapes.
	 
    IsCompoundManifold(TheS : Compound  from  TopoDS) returns Boolean from Standard;
    	---Purpose: to check if TheS is manifol or not.
	-- compound conciders to  be manifold if:
	-- 1) all shapes in compound are manifold (see comments for method IsManifold)
	-- 2) all shapes are fully disconnected - there are any shapes in  compound that 
	--    share common subshapes.
	 
	 
    TypeOfShape(TheS : Shape  from  TopoDS) returns ShapeEnum from TopAbs;	
    	---Purpose: to define if COMPOUND is homogeneous  
    	-- (consists of shapes of the same type) and return this shape type. 
	-- If COMPOUND is mixed, method returns TopAbs_COMPOUND.  
	-- If TheS is single shape (not COMPOUND), method returns its type. 
	-- If COMPOUND contains nested compounds, it concideres to be homogeneous 
	-- if all compounds consist of shapes of the same type.	 
	
    IsConnected(TheS : Shape  from  TopoDS) returns Boolean from Standard;
    	---Purpose: to check if all subshapes in TheS, when TheS is COMPOUND, COMPSOLID, SHELL or WIRE,  
    	-- are linked through common faces, edges or  vertices.
	-- SOLID, FACE, EDGE, VERTEX concider to be connected by default.  
	 

    end  QANewModTopOpe;	
