-- Created on: 1993-07-19
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Curve2dSet from GeomTools 

	---Purpose: Stores a set of Curves from Geom2d.

uses
    Curve                 from Geom2d,
    IndexedMapOfTransient from TColStd,
    ProgressIndicator     from Message
    
raises
    OutOfRange from Standard

is

    Create returns Curve2dSet from GeomTools;
	---Purpose: Returns an empty set of Curves.
	
    Clear(me : in out)
	---Purpose: Clears the content of the set.
    is static;
	
    Add(me : in out; C : Curve from Geom2d) returns Integer
	---Purpose: Incorporate a new Curve in the  set and returns
	--          its index.
    is static;
    
    Curve2d(me; I : Integer) returns Curve from Geom2d
	---Purpose: Returns the Curve of index <I>.
    raises
    	OutOfRange from Standard
    is static;

    Index(me; C : Curve from Geom2d) returns Integer
	---Purpose: Returns the index of <L>.
    is static;
    
    Dump(me; OS : in out OStream)
	---Purpose: Dumps the content of me on the stream <OS>.
    is static;
	
    Write(me; OS : in out OStream)
	---Purpose: Writes the content of  me  on the stream <OS> in a
	--          format that can be read back by Read.
    is static;
	
    Read(me : in out; IS : in out IStream)
	---Purpose: Reads the content of me from the  stream  <IS>. me
	--          is first cleared.
	--          
    is static;
    
    --
    -- 	class methods to write an read curves
    -- 	
    
    PrintCurve2d(myclass; C  : Curve from Geom2d;
    	    	    	  OS : in out OStream;
			  compact : Boolean = Standard_False);
	---Purpose: Dumps the curve on the stream,  if compact is True
	--          use the compact format that can be read back.
	
    ReadCurve2d(myclass; IS : in out IStream;
    	    	    	 C  : in out Curve from Geom2d)
    returns IStream;
	---Purpose: Reads the curve  from  the stream.  The  curve  is
	--          assumed   to have  been  writtent  with  the Print
	--          method (compact = True).
	--          
	---C++: return &
	
    SetProgress(me : in out; PR : ProgressIndicator from Message);

    GetProgress(me) returns ProgressIndicator from Message;

fields

    myMap : IndexedMapOfTransient from TColStd;
    myProgress : ProgressIndicator from Message;

end Curve2dSet;


