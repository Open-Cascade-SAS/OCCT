-- Created on: 2002-12-12
-- Created by: data exchange team
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class ParametricCurve3dElementCoordinateSystem from StepFEA
inherits FeaRepresentationItem from StepFEA

    ---Purpose: Representation of STEP entity ParametricCurve3dElementCoordinateSystem

uses
    HAsciiString from TCollection,
    ParametricCurve3dElementCoordinateDirection from StepFEA

is
    Create returns ParametricCurve3dElementCoordinateSystem from StepFEA;
	---Purpose: Empty constructor

    Init (me: mutable; aRepresentationItem_Name: HAsciiString from TCollection;
                       aDirection: ParametricCurve3dElementCoordinateDirection from StepFEA);
	---Purpose: Initialize all fields (own and inherited)

    Direction (me) returns ParametricCurve3dElementCoordinateDirection from StepFEA;
	---Purpose: Returns field Direction
    SetDirection (me: mutable; Direction: ParametricCurve3dElementCoordinateDirection from StepFEA);
	---Purpose: Set field Direction

fields
    theDirection: ParametricCurve3dElementCoordinateDirection from StepFEA;

end ParametricCurve3dElementCoordinateSystem;
