-- Created on: 1999-03-05
-- Created by: Fabrice SERVANT
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Point from IntPolyh

uses
    
    Pnt from gp,
    HSurface from Adaptor3d

is


    Create;
    
    Create(xx,yy,zz,uu,vv : Real from Standard); 

    X(me) 
    returns Real from Standard
    is static;

    Y(me) 
    returns Real from Standard
    is static;

    Z(me) 
    returns Real from Standard
    is static;

    U(me) 
    returns Real from Standard
    is static;

    V(me) 
    returns Real from Standard
    is static;
    
    PartOfCommon(me)
    returns Integer from Standard
    is static;
    
    Equal(me: in out; Pt: Point from IntPolyh)
        ---C++: alias operator =
    is static;
	
    Set(me: in out; v1,v2,v3,v4,v5: Real from Standard; II: Integer from Standard = 1)
    is static;
	
    SetX(me: in out; v: Real from Standard) 
    is static;
	
    SetY(me: in out; v: Real from Standard) 
    is static;
	
    SetZ(me: in out; v: Real from Standard) 
    is static;
	
    SetU(me: in out; v: Real from Standard) 
    is static;
	
    SetV(me: in out; v: Real from Standard) 
    is static;
    
    SetPartOfCommon(me :in out; ii: Integer from Standard)
    is static;
    
    Middle(me: in out; MySurface: HSurface from Adaptor3d; P1,P2: Point from IntPolyh)
    is static;

    Add(me; P1: Point from IntPolyh)
    	---C++: alias operator +     
    returns Point from IntPolyh
    is static;
    
    Sub(me; P1: Point from IntPolyh)
    	---C++: alias operator -     
    returns Point from IntPolyh
    is static;
    
    Divide(me; rr: Real from Standard)
    	---C++: alias operator /     
    returns Point from IntPolyh
    is static;    
    
    Multiplication(me; rr: Real from Standard)
    	---C++: alias operator *     
    returns Point from IntPolyh
    is static;    
    
    SquareModulus(me)
    returns Real from Standard
    is static;       

    SquareDistance(me; P2: Point from IntPolyh)
    returns Real from Standard
    is static;       
          
    Dot(me; P2: Point from IntPolyh)
    returns Real from Standard
    is static;   

    Cross(me:in out; P1,P2: Point from IntPolyh)
    is static;
		
    Dump(me) 
    is static;
    
    Dump(me; i: Integer from Standard)
    is static; 
    
--modified by NIZNHY-PKV Fri Jan 20 12:11:36 2012 f   
    SetDegenerated(me:out; 
    	    theFlag:Boolean from Standard);   
  
    Degenerated(me) 
    	returns Boolean from Standard; 
--modified by NIZNHY-PKV Fri Jan 20 12:12:07 2012t	 
 
fields
    x,y,z,u,v : Real from Standard;
    POC : Integer from Standard; 
    --modified by NIZNHY-PKV Fri Jan 20 12:17:39 2012f
    myDegenerated : Boolean from Standard; 
    --modified by NIZNHY-PKV Fri Jan 20 12:17:41 2012t
    
end Point from IntPolyh;



