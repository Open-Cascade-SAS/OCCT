-- File:	RWStepDimTol_RWDatumFeature.cdl
-- Created:	Wed Jun  4 13:34:35 2003 
-- Author:	Galina KULIKOVA
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWDatumFeature from RWStepDimTol

    ---Purpose: Read & Write tool for DatumFeature

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    DatumFeature from StepDimTol

is
    Create returns RWDatumFeature from RWStepDimTol;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : DatumFeature from StepDimTol);
	---Purpose: Reads DatumFeature

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: DatumFeature from StepDimTol);
	---Purpose: Writes DatumFeature

    Share (me; ent : DatumFeature from StepDimTol;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWDatumFeature;
