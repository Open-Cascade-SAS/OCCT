-- File:	IGESDimen_ToolSection.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolSection  from IGESDimen

    ---Purpose : Tool to work on a Section. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses Section from IGESDimen,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolSection;
    ---Purpose : Returns a ToolSection, ready to work


    ReadOwnParams (me; ent : mutable Section;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : Section;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : Section;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a Section <ent>, from
    --           its specific (own) parameters

    OwnCorrect (me; ent : mutable Section) returns Boolean  is static;
    ---Purpose : Sets automatic unambiguous Correction on a Section
    --           (LineFont forced to Rank = 1, DataType forced to 1)

    DirChecker (me; ent : Section) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : Section;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : Section; entto : mutable Section;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : Section;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolSection;
