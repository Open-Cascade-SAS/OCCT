-- Created by: DAUTRY Philippe
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

--      	-------------------

---Version:	0.0
--Version	Date		Purpose
--		0.0	May 26 1997	Creation


class ClosureMode from TDF

	---Purpose: This class provides options closure management.

-- uses

-- raises

is

    Create(aMode : Boolean from Standard = Standard_True)
    	returns ClosureMode from TDF;
	---Purpose: Creates an objet with all modes set to <aMode>.


    Descendants(me : in out; aStatus : Boolean from Standard);
	---Purpose: Sets the mode "Descendants" to <aStatus>.
	--          
	--          "Descendants" mode means we add to the data set
	--          the children labels of each USER GIVEN label. We
	--          do not do that with the labels found applying
	--          UpToFirstLevel option.
	--          
	---C++: inline

    Descendants(me) returns Boolean from Standard;
	---Purpose: Returns true if the mode "Descendants" is set.
	--          
	---C++: inline


    References(me : in out; aStatus : Boolean from Standard);
	---Purpose: Sets the mode "References" to <aStatus>.
	--          
	--          "References" mode means we add to the data set
	--          the descendants of an attribute, by calling the
	--          attribute method Descendants().
	--          
	---C++: inline

    References(me) returns Boolean from Standard;
	---Purpose: Returns true if the mode "References" is set.
	--          
	---C++: inline


fields

    myFlags : Integer from Standard;
    -- Bit Mask Use
    -- 0   1    Descendants
    -- 1   2    References
    -- 2   4    Unused

end ClosureMode;
