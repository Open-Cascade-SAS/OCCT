-- Created on: 2003-01-14
-- Created by: data exchange team
-- Copyright (c) 2003-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class SymmetricTensor43dMember from StepFEA inherits SelectArrReal from StepData
    
    ---Purpose: Representation of member for  STEP SELECT type SymmetricTensor43d

is
    Create returns SymmetricTensor43dMember from StepFEA;
    ---Purpose: Empty constructor

    HasName (me) returns Boolean  is redefined;
    ---Purpose: Returns True if has name

    Name (me) returns CString  is redefined;
    ---Purpose: Returns set name

    SetName (me : mutable; name : CString)  returns Boolean  is redefined;
    ---Purpose: Set name

    Matches (me; name : CString) returns Boolean  is redefined;
    ---Purpose : Tells if the name of a SelectMember matches a given one;

fields

    mycase : Integer;                                                                                                         

end SymmetricTensor43dMember;
