-- Created on: 2006-08-07
-- Created by: Galina KULIKOVA
-- Copyright (c) 2006-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class FaceDivideArea from ShapeUpgrade inherits FaceDivide from ShapeUpgrade

	---Purpose: Divides face by max area criterium.

uses
    Face from TopoDS

is

    Create returns FaceDivideArea from ShapeUpgrade; 
        ---Purpose: Creates empty  constructor.

    Create (F : Face from TopoDS) returns FaceDivideArea from ShapeUpgrade;
    
    Perform (me: mutable) returns Boolean is redefined;
        ---Purpose: Performs splitting and computes the resulting shell
	--          The context is used to keep track of former splittings
    
    MaxArea(me: mutable) returns Real;
    ---C++: inline
    ---C++: return &
    ---Purpose:Set max area allowed for faces
     
fields

    myMaxArea : Real;

end FaceDivideArea;
