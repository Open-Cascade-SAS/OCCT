-- Created on: 1994-09-15
-- Created by: Bruno DUMORTIER
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ProjectOnSurface from ProjLib 

uses

    HCurve       from Adaptor3d,
    HSurface     from Adaptor3d,
    BSplineCurve from Geom

is

    Create 
    	---Purpose:  Create an empty projector.
    returns ProjectOnSurface from ProjLib;
    

    Create( S  : HSurface from Adaptor3d)
    	---Purpose: Create a projector normaly to the surface <S>.
    returns ProjectOnSurface from ProjLib;

    Delete(me:out) is virtual;
    ---C++: alias "Standard_EXPORT virtual ~ProjLib_ProjectOnSurface(){Delete() ; }"
    
    Load(me : in out; S : HSurface from Adaptor3d)
	---Purpose: Set the Surface to <S>.
	--          To compute the projection, you have to Load the Curve.
    is static;
    
    Load(me : in out; C : HCurve from Adaptor3d; Tolerance : Real)
	---Purpose: Compute the projection of the curve <C> on the Surface.
    is static;

    IsDone(me) returns Boolean ;
    
    BSpline(me) returns BSplineCurve from Geom  
    is static ;

fields

    myCurve      : HCurve   from Adaptor3d ;
    mySurface    : HSurface from Adaptor3d ;
    myTolerance  : Real ;
    myIsDone     : Boolean ;
    myResult     : BSplineCurve from Geom ;

end ProjectOnSurface;
