-- Created on: 1992-04-03
-- Created by: Laurent BUCHARD
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



package IntRes2d


    ---Purpose: This package provides the definition of the results of
    --          the intersection between 2D curves and the definition
    --          of a domain on a 2D curve.
    ---Level: Public 
    -- 
    -- All the methods of all the classes of this package are public.
    --

uses

    Standard, TCollection, gp, StdFail

is


    class IntersectionPoint;
    
    class IntersectionSegment;

    class Transition;

    class Domain;

    deferred class Intersection;

    enumeration Position is Head,Middle,End;

    enumeration TypeTrans is In,Out,Touch,Undecided;

    enumeration Situation is Inside, Outside, Unknown;

    class SequenceOfIntersectionPoint instantiates
    	       Sequence from TCollection (IntersectionPoint);

    class SequenceOfIntersectionSegment instantiates
    	       Sequence from TCollection (IntersectionSegment);


end IntRes2d; 


