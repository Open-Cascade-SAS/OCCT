-- File:	Geom2dAdaptor_HCurve.cdl
-- Created:	Fri Aug 25 14:38:16 1995
-- Author:	Remi LEQUETTE
--		<rle@mentox>
---Copyright:	 Matra Datavision 1995



class HCurve from Geom2dAdaptor inherits GHCurve from Geom2dAdaptor

	---Purpose: Provides an interface between the services provided by any
    	-- curve from the package Geom2d and those required
    	-- of the curve by algorithms, which use it.

uses
    Curve from Geom2d,
    Curve from Geom2dAdaptor

raises
    ConstructionError from Standard

is

    Create returns mutable HCurve from Geom2dAdaptor;
    
    Create( AS : Curve from Geom2dAdaptor) returns mutable HCurve from Geom2dAdaptor;

    Create( S : Curve from Geom2d) returns mutable HCurve from Geom2dAdaptor;
    
    Create( S : Curve from Geom2d; UFirst,ULast : Real) 
    returns  mutable HCurve from Geom2dAdaptor
    raises ConstructionError from Standard;
    	---Purpose: ConstructionError is raised if UFirst>ULast or VFirst>VLast

end HCurve;
