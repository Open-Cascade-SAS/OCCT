-- Created on: 1993-01-09
-- Created by: CKY / Contract Toubro-Larsen ( Arun MENON )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class OrderedGroup from IGESBasic  inherits Group

        ---Purpose: defines OrderedGroup, Type <402> Form <14>
        --          in package IGESBasic
        --          this class defines an Ordered Group with back pointers
        --          
        --          It inherits from Group

uses

        Transient        ,
        HArray1OfIGESEntity from IGESData

raises OutOfRange

is

        Create returns mutable OrderedGroup;

        -- Specific Methods pertaining to the class : see Group

--
-- Class    : IGESBasic_OrderedGroup
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class OrderedGroup.
--
-- Reminder : A OrderedGroup instance is defined by :
--            - an array of entities
--            See Group

end OrderedGroup;
