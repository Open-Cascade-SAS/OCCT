-- Created on: 2003-08-21
-- Created by: Sergey KUUL
-- Copyright (c) 2003-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ReprItemAndLengthMeasureWithUnit from StepRepr inherits RepresentationItem from StepRepr

uses
    LengthMeasureWithUnit from StepBasic,
    MeasureRepresentationItem from StepRepr,
    MeasureWithUnit from StepBasic

is

    Create returns mutable ReprItemAndLengthMeasureWithUnit;
    
    Init(me: mutable; aMWU: mutable MeasureWithUnit; aRI : RepresentationItem);

    SetLengthMeasureWithUnit(me: mutable; aLMWU: mutable LengthMeasureWithUnit);
    
    GetLengthMeasureWithUnit(me) returns mutable LengthMeasureWithUnit;

    GetMeasureRepresentationItem(me) returns mutable MeasureRepresentationItem;

    SetMeasureWithUnit(me: mutable; aMWU: mutable MeasureWithUnit);
    
    GetMeasureWithUnit(me) returns mutable MeasureWithUnit;

    GetRepresentationItem(me) returns mutable RepresentationItem;

fields

    myLengthMeasureWithUnit: LengthMeasureWithUnit from StepBasic;
    myMeasureRepresentationItem : MeasureRepresentationItem from StepRepr;
    myMeasureWithUnit: MeasureWithUnit from StepBasic;

end ReprItemAndLengthMeasureWithUnit;
