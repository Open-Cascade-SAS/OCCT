-- Created on: 2003-01-22
-- Created by: data exchange team
-- Copyright (c) 2003-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class FeaCurveSectionGeometricRelationship from StepFEA
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity FeaCurveSectionGeometricRelationship

uses
    CurveElementSectionDefinition from StepElement,
    AnalysisItemWithinRepresentation from StepElement

is
    Create returns FeaCurveSectionGeometricRelationship from StepFEA;
	---Purpose: Empty constructor

    Init (me: mutable; aSectionRef: CurveElementSectionDefinition from StepElement;
                       aItem: AnalysisItemWithinRepresentation from StepElement);
	---Purpose: Initialize all fields (own and inherited)

    SectionRef (me) returns CurveElementSectionDefinition from StepElement;
	---Purpose: Returns field SectionRef
    SetSectionRef (me: mutable; SectionRef: CurveElementSectionDefinition from StepElement);
	---Purpose: Set field SectionRef

    Item (me) returns AnalysisItemWithinRepresentation from StepElement;
	---Purpose: Returns field Item
    SetItem (me: mutable; Item: AnalysisItemWithinRepresentation from StepElement);
	---Purpose: Set field Item

fields
    theSectionRef: CurveElementSectionDefinition from StepElement;
    theItem: AnalysisItemWithinRepresentation from StepElement;

end FeaCurveSectionGeometricRelationship;
