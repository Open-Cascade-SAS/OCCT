-- File:	StepDimTol_Datum.cdl
-- Created:	Wed Jun  4 13:34:34 2003 
-- Author:	Galina KULIKOVA
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class Datum from StepDimTol
inherits ShapeAspect from StepRepr

    ---Purpose: Representation of STEP entity Datum

uses
    HAsciiString from TCollection,
    ProductDefinitionShape from StepRepr,
    Logical from StepData

is
    Create returns Datum from StepDimTol;
	---Purpose: Empty constructor

    Init (me: mutable; aShapeAspect_Name: HAsciiString from TCollection;
                       aShapeAspect_Description: HAsciiString from TCollection;
                       aShapeAspect_OfShape: ProductDefinitionShape from StepRepr;
                       aShapeAspect_ProductDefinitional: Logical from StepData;
                       aIdentification: HAsciiString from TCollection);
	---Purpose: Initialize all fields (own and inherited)

    Identification (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Identification
    SetIdentification (me: mutable; Identification: HAsciiString from TCollection);
	---Purpose: Set field Identification

fields
    theIdentification: HAsciiString from TCollection;

end Datum;
