-- Created on: 2002-12-12
-- Created by: data exchange team
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class CurveElementInterval from StepFEA
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity CurveElementInterval

uses
    CurveElementLocation from StepFEA,
    EulerAngles from StepBasic

is
    Create returns CurveElementInterval from StepFEA;
	---Purpose: Empty constructor

    Init (me: mutable; aFinishPosition: CurveElementLocation from StepFEA;
                       aEuAngles: EulerAngles from StepBasic);
	---Purpose: Initialize all fields (own and inherited)

    FinishPosition (me) returns CurveElementLocation from StepFEA;
	---Purpose: Returns field FinishPosition
    SetFinishPosition (me: mutable; FinishPosition: CurveElementLocation from StepFEA);
	---Purpose: Set field FinishPosition

    EuAngles (me) returns EulerAngles from StepBasic;
	---Purpose: Returns field EuAngles
    SetEuAngles (me: mutable; EuAngles: EulerAngles from StepBasic);
	---Purpose: Set field EuAngles

fields
    theFinishPosition: CurveElementLocation from StepFEA;
    theEuAngles: EulerAngles from StepBasic;

end CurveElementInterval;
