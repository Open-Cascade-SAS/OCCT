-- File:	RWStl.cdl
-- Created:	Thu Oct 13 12:57:13 1994
-- Author:	Marc LEGAY
--		<mle@bourdon>
---Copyright:	 Matra Datavision 1994

package RWStl 

	---Purpose: This package contains the methods to be used in 
	--          the Stereo Lithograpy Application. The main 
	--          features of this application are ,starting from a 
	--          Shape :
	--          - mesh this shape with a maximun tolerance,
	--          - display the meshing,
	--          - write the meshing in a file (binary or ascii),
	--          - read of file (binary or ascii) and display it,
	--          - translate a binary file to an ascii file,
	--          - translate an ascii file to an binary file. 
    	    	    	    	    	    	    	    	    	
uses 

    OSD, 
    Standard, 
    StlMesh,
    Message
    
is 

	WriteBinary (aMesh : Mesh from StlMesh; aPath : Path from OSD;
	    aProgInd : ProgressIndicator from Message = NULL) 
    	    	returns Boolean from Standard;
	  ---Purpose : write the meshing in a file following the 
	  --         binary format of an STL file.
	  --         Returns false if the cannot be opened; 	    	

	WriteAscii (aMesh : Mesh from StlMesh; aPath : Path from OSD;
	    aProgInd : ProgressIndicator from Message = NULL) 
    	    	returns Boolean from Standard;
	  ---Purpose : write the meshing in a file following the 
	  --         Ascii  format of an STL file. 	    	
	  --         Returns false if the cannot be opened; 	    	


    	ReadFile   (aPath : Path from OSD;
	    aProgInd : ProgressIndicator from Message = NULL) returns
    	    	Mesh from StlMesh;
	  ---Purpose : This method will chwck if the file is a binary 
	  --         file or an AsciiFile testing  the 5 first 
	  --         characters of the file wich are :"solid" in an 
	  --         ascii file. If we do not find that word we assume 
	  --         that it is a binary file.	

    	ReadBinary (aPath : Path from OSD;
	    aProgInd : ProgressIndicator from Message = NULL) returns 
    	    	Mesh from StlMesh;
	 ---Purpose : Read a meshing from a binary file
	 --        Raises NoMoreObject from Standard if a statement 
	 --        does not contain the right number of tokens
	 --        Raises TypeMisMatch if a token has not the good 
	 --        type (often real)

    	ReadAscii (aPath : Path from OSD;
	    aProgInd : ProgressIndicator from Message = NULL) returns 
    	    	Mesh from StlMesh;
	 ---Purpose : Read a meshing from a binary file
	 --        Raises NoMoreObject from Standard if a statement 
	 --        does not contain the right number of tokens
	 --        Raises TypeMisMatch if a token has not the good 
	 --        type (often real)
	 --        Raises MoMoreObject if a file is finished before 
	 --        having found the word endsolid;

end RWStl;



