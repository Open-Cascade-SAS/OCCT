-- Created on: 1993-12-02
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



package Blend

uses IntSurf, 
    TColgp, 
    TColStd, 
    Adaptor2d, 
    gp, 
    TopAbs, 
    math, 
    TCollection, 
    MMgt, 
    StdFail,  
    GeomAbs

is

--    deferred generic class SurfaceTool;
    
    generic class Iterator;          -- template class

    deferred class AppFunction;      -- inherits FunctionSetWithDerivatives from math

    deferred class Function;         -- inherits AppFunction from Blend

    deferred class FuncInv;          -- inherits FunctionSetWithDerivatives from math

    deferred class CSFunction;       -- inherits AppFunction from Blend

    deferred class SurfRstFunction;  -- inherits AppFunction from Blend

    deferred class SurfPointFuncInv; -- inherits FunctionSetWithDerivatives from math

    deferred class SurfCurvFuncInv;  -- inherits FunctionSetWithDerivatives from math

    deferred class RstRstFunction;  -- inherits AppFunction from Blend

    deferred class CurvPointFuncInv; -- inherits FunctionSetWithDerivatives from math



    class Point;
    
    generic class Extremity;
    
    generic class PointOnRst;
    
    generic class Line;

    generic class Walking;

    generic class CSWalking;


    class SequenceOfPoint instantiates Sequence from TCollection
    	(Point from Blend);
	
    enumeration Status is 
    	StepTooLarge,
	StepTooSmall,
	Backward,
	SamePoints,
	OnRst1,
	OnRst2,
	OnRst12,
	OK
    end Status;


    enumeration DecrochStatus is 
    	NoDecroch,
	DecrochRst1,
	DecrochRst2,
	DecrochBoth
    end Status;



end Blend;
