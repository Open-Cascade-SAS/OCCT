-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PointStyle from StepVisual 

inherits TShared from MMgt

uses

	HAsciiString from TCollection, 
	MarkerSelect from StepVisual, 
	SizeSelect from StepBasic, 
	Colour from StepVisual
is

	Create returns PointStyle;
	---Purpose: Returns a PointStyle

	Init (me : mutable;
	      aName : HAsciiString from TCollection;
	      aMarker : MarkerSelect from StepVisual;
	      aMarkerSize : SizeSelect from StepBasic;
	      aMarkerColour : Colour from StepVisual) is virtual;

	-- Specific Methods for Field Data Access --

	SetName(me : mutable; aName : HAsciiString);
	Name (me) returns HAsciiString;
	SetMarker(me : mutable; aMarker : MarkerSelect);
	Marker (me) returns MarkerSelect;
	SetMarkerSize(me : mutable; aMarkerSize : SizeSelect);
	MarkerSize (me) returns SizeSelect;
	SetMarkerColour(me : mutable; aMarkerColour : Colour);
	MarkerColour (me) returns Colour;

fields

	name : HAsciiString from TCollection;
	marker : MarkerSelect from StepVisual; -- a SelectType
	markerSize : SizeSelect from StepBasic; -- a SelectType
	markerColour : Colour from StepVisual;

end PointStyle;
