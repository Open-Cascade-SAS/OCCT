-- Created on: 1997-08-07
-- Created by: VAUTHIER Jean-Claude 
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- modified     Sergey Zaritchny



package MDataStd 

	---Purpose: Storage    and  Retrieval  drivers   for modelling
	--          attributes.   Transient  attributes are defined in
	--          package TDataStd and persistent one are defined in
	--          package PDataStd

uses TDF,
     PDF,
     MDF, 
     CDM,
     TDataStd

is

    	---Purpose: Storage drivers for TDataStd attributes
    	--          =======================================

	
        class DirectoryStorageDriver;

	class UAttributeStorageDriver;
	
    	class NameStorageDriver;

    	class CommentStorageDriver;

 	class IntegerStorageDriver;
	
	class IntegerArrayStorageDriver;
	
    	class RealStorageDriver;

	class RealArrayStorageDriver;
	
	class ExtStringArrayStorageDriver;	

    	class VariableStorageDriver;

    	class ExpressionStorageDriver;

    	class RelationStorageDriver;    
	
	class NoteBookStorageDriver;

    	class TreeNodeStorageDriver;
	
    	 
    --Extension 
	class TickStorageDriver;
        class IntegerListStorageDriver;
        class RealListStorageDriver;
        class ExtStringListStorageDriver;
        class BooleanListStorageDriver;
        class ReferenceListStorageDriver;
        class BooleanArrayStorageDriver;
        class ReferenceArrayStorageDriver;
        class ByteArrayStorageDriver;
        class NamedDataStorageDriver;
        class AsciiStringStorageDriver; 
        class IntPackedMapStorageDriver; 
    
    	---Purpose: Retrieval drivers for PDataStd attributes
    	--          =========================================

        class DirectoryRetrievalDriver;

	class UAttributeRetrievalDriver;
	
    	class NameRetrievalDriver;

    	class CommentRetrievalDriver;

 	class IntegerRetrievalDriver;
	
        class IntegerArrayRetrievalDriver; 
	 
        class IntegerArrayRetrievalDriver_1;	

    	class RealRetrievalDriver;

	class RealArrayRetrievalDriver; 
	 
	class RealArrayRetrievalDriver_1;	
	
	class ExtStringArrayRetrievalDriver;

	class ExtStringArrayRetrievalDriver_1;  	

	class VariableRetrievalDriver;

    	class ExpressionRetrievalDriver;

    	class RelationRetrievalDriver;	   

	class NoteBookRetrievalDriver;

    	class TreeNodeRetrievalDriver;

	  
	--  Extension 
	class TickRetrievalDriver;
        class IntegerListRetrievalDriver;
        class RealListRetrievalDriver;
        class ExtStringListRetrievalDriver;
        class BooleanListRetrievalDriver;
        class ReferenceListRetrievalDriver;
        class BooleanArrayRetrievalDriver;
        class ReferenceArrayRetrievalDriver;
        class ByteArrayRetrievalDriver; 
	class ByteArrayRetrievalDriver_1;
        class NamedDataRetrievalDriver; 
        class AsciiStringRetrievalDriver; 
        class IntPackedMapRetrievalDriver;     
    	class IntPackedMapRetrievalDriver_1;


    AddStorageDrivers(aDriverSeq : ASDriverHSequence from MDF; theMessageDriver : MessageDriver from CDM);
	---Purpose: Adds the attribute storage drivers to <aDriverSeq>.


    AddRetrievalDrivers(aDriverSeq : ARDriverHSequence from MDF; theMessageDriver : MessageDriver from CDM);
	---Purpose: Adds the attribute retrieval drivers to <aDriverSeq>.


    ---Purpose: Translation of TDataStd enumerations to integer
    --          ===============================================

    RealDimensionToInteger (e : RealEnum from TDataStd)
    returns Integer from Standard;

    IntegerToRealDimension (i : Integer from Standard)
    returns RealEnum from TDataStd;
     
end MDataStd;
