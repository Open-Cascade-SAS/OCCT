-- File:        ColourRgb.cdl
-- Created:     Mon Dec  4 12:02:24 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWColourRgb from RWStepVisual

	---Purpose : Read & Write Module for ColourRgb

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     ColourRgb from StepVisual

is

	Create returns RWColourRgb;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable ColourRgb from StepVisual);

	WriteStep (me; SW : in out StepWriter; ent : ColourRgb from StepVisual);

end RWColourRgb;
