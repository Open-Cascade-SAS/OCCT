-- Created on: 1996-01-23
-- Created by: s:       LAVNIKOV Alexey, PLOTNIKOV Eugeny & CHABROVSKY Dmitry
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Modifications: DCB at March 1998  Porting MFT for Windows NT (95)
--                PLOTNIKOV Eugeny at July 1998 (BUC60286)

package WNT

        ---Purpose: This package contains common Windows NT graphics interface.

 uses

    Aspect,
    Image,
    Quantity,
    TCollection,
    TColStd,
    TShort,
    MMgt,
    OSD

 is


        -----------------------
        -- Category: Exceptions
        -----------------------


    exception ClassDefinitionError inherits ConstructionError;
        ---Category: Exceptions


        --------------------
        -- Category: Classes
        --------------------

    class Window;
        ---Category: Classes

    class WClass;
        ---Category: Classes

        ---------------------------
        -- Category: Enumerations
        ---------------------------

    enumeration OrientationType is

        OT_PORTRAIT,
        OT_LANDSCAPE

    end OrientationType;
---Purpose: Portrait/landscape orientation.


        ---------------------------
        -- Category: Imported types
        ---------------------------


    imported Dword;
        ---Category: Imported types

    imported Uint;
        ---Category: Imported types

        ---------------------------------
        -- Category: Pointers
        ---------------------------------

    pointer WindowPtr to Window from WNT;

end WNT;
