-- File:        SolidModel.cdl
-- Created:     Mon Dec  4 12:02:31 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWSolidModel from RWStepShape

	---Purpose : Read & Write Module for SolidModel

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     SolidModel from StepShape

is

	Create returns RWSolidModel;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable SolidModel from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : SolidModel from StepShape);

end RWSolidModel;
