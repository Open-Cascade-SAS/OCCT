-- Created on: 2018-03-15
-- Created by: Stephan GARNAUD (ARM)
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.





class Host from OSD

 ---Purpose: Carries information about a Host


uses SysType, OEMType, Error, AsciiString from TCollection
raises ConstructionError, NullObject, OSDError

 is

  Create returns Host;
    ---Purpose: Initializes current host by default.
    ---Level: Advanced

  SystemVersion (me : in out) returns AsciiString is static;
    ---Purpose: Returns system name and version
    ---Level: Advanced

  SystemId (me) returns SysType is static;
    ---Purpose: Returns the system type (UNIX System V, UNIX BSD, MS-DOS...)
    ---Level: Advanced

  HostName (me : in out) returns AsciiString is static;
    ---Purpose: Returns host name.
    ---Level: Advanced

  AvailableMemory (me : in out)  returns Integer is static;
    ---Purpose: Returns available memory in Kilobytes.
    ---Level: Obsolete syntax. Will be removed in next version

  InternetAddress (me : in out) returns AsciiString is static;
    ---Purpose: Returns Internet address of current host.
    ---Level: Advanced

  MachineType (me : in out) returns OEMType is static;
    ---Purpose: Returns type of current machine.
    ---Level: Advanced

 Failed (me) returns Boolean is static;
   ---Purpose: Returns TRUE if an error occurs
   ---Level: Advanced

 Reset (me : in out) is static;
   ---Purpose: Resets error counter to zero
   ---Level: Advanced
      
 Perror (me : in out)
   ---Purpose: Raises OSD_Error
   ---Level: Advanced
   raises OSDError is static;

 Error (me) returns Integer is static;
   ---Purpose: Returns error number if 'Failed' is TRUE.
   ---Level: Advanced

fields
  myName   : AsciiString;
  myError  : Error;
end Host from OSD;


