-- Created on: 1993-04-22
-- Created by: Christian CAILLET
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class HGraph  from Interface  inherits TShared

    ---Purpose : This class allows to store a redefinable Graph, via a Handle
    --           (usefull for an Object which can work on several successive
    --           Models, with the same general conditions)

uses Graph, InterfaceModel, GeneralLib, Protocol, GTool

raises DomainError

is

    Create (agraph : Graph) returns mutable HGraph;
    ---Purpose : Creates an HGraph directly from a Graph.
    --           Remark that the starting Graph is duplicated
    
    Create (amodel : InterfaceModel; lib : GeneralLib;
     theModeStats : Boolean = Standard_True) returns mutable HGraph;
    ---Purpose : Creates an HGraph with a Graph created from <amodel> and <lib>

    Create (amodel : InterfaceModel; protocol : Protocol from Interface;
     theModeStats : Boolean = Standard_True)
    	returns mutable HGraph;
    ---Purpose : Creates an HGraph with a graph itself created from <amodel>
    --           and <protocol>

    Create (amodel : InterfaceModel; gtool : GTool from Interface;
     theModeStats : Boolean = Standard_True)
    	returns mutable HGraph;
    ---Purpose : Creates an HGraph with a graph itself created from <amodel>
    --           and <protocol>

    Create (amodel : InterfaceModel;
     theModeStats : Boolean = Standard_True) returns mutable HGraph
    ---Purpose : Same a above, but works with the GTool in the model
    	raises DomainError;
    --           Error if no Active Protocol is defined

    Graph (me) returns Graph;
    ---Purpose : Returns the Graph contained in <me>, for Read Only Operations
    --           Remark that it is returns as "const &"
    --           Getting it in a new variable instead of a reference would be
    --           a pitty, because all the graph's content would be duplicated
    ---C++ : return const &

    CGraph (me : mutable) returns Graph;
    ---Purpose : Same as above, but for Read-Write Operations
    --           Then, The Graph will be modified in the HGraph itself
    ---C++ : return &

fields

    thegraph : Graph;

end HGraph;
