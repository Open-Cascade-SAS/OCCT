-- Created on: 1995-02-08
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

private class ParameterAndOrientation from GeomInt

	---Purpose: 

uses Orientation from TopAbs

is

    Create
    
    	returns ParameterAndOrientation from GeomInt;


    Create(P: Real from Standard; Or1,Or2: Orientation from TopAbs)
    
    	returns ParameterAndOrientation from GeomInt;


    SetOrientation1(me: in out; Or: Orientation from TopAbs)
    
    	is static;


    SetOrientation2(me: in out; Or: Orientation from TopAbs)
    
    	is static;


    Parameter(me)
    
    	returns Real from Standard
	is static;


    Orientation1(me)
    
    	returns Orientation from TopAbs
    	is static;


    Orientation2(me)
    
    	returns Orientation from TopAbs
    	is static;


fields

    prm : Real from Standard;
    or1 : Orientation from TopAbs;
    or2 : Orientation from TopAbs;

end ParameterAndOrientation;
