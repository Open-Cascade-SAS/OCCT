-- Created on: 1994-02-18
-- Created by: Bruno DUMORTIER
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Line from GeomFill

	---Purpose: 

inherits TShared from MMgt


is

    Create returns mutable Line from GeomFill;

    Create(NbPoints : Integer from Standard)
    returns mutable Line from GeomFill;

    NbPoints(me)
    returns Integer from Standard
	---C++: inline
    is static;


    Point(me; Index: Integer from Standard)
    returns Integer  from Standard
	---C++: inline
    is static;

fields

    myNbPoints : Integer from Standard;

end Line;
