-- Created on: 1998-10-29
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Hctxff2d from TopOpeBRep inherits TShared from  MMgt

uses

    Shape from TopoDS,
    Face from TopoDS,
    HSurface from BRepAdaptor,
    Surface from BRepAdaptor,
    SurfaceType from GeomAbs

is

    Create returns mutable Hctxff2d from TopOpeBRep;
    SetFaces(me:mutable; F1,F2:Face);
    SetHSurfaces(me:mutable; S1,S2:HSurface from BRepAdaptor);
    SetHSurfacesPrivate(me:mutable) is private;
    SetTolerances(me:mutable;Tol1,Tol2:Real);
    GetTolerances(me;Tol1,Tol2:out Real);
    GetMaxTolerance(me) returns Real;
    Face(me;I:Integer) returns Face;---C++ : return const &
    HSurface(me;I:Integer) returns HSurface from BRepAdaptor;
    SurfacesSameOriented(me) returns Boolean;
    FacesSameOriented(me) returns Boolean;
    FaceSameOrientedWithRef(me;I:Integer) returns Boolean;

fields

    myFace1 : Face from TopoDS;
    mySurface1 : HSurface from BRepAdaptor;
    mySurfaceType1 : SurfaceType from GeomAbs;
    myf1surf1F_sameoriented : Boolean;

    myFace2 : Face from TopoDS;
    mySurface2 : HSurface from BRepAdaptor;
    mySurfaceType2 : SurfaceType from GeomAbs;
    myf2surf1F_sameoriented : Boolean;

    mySurfacesSameOriented : Boolean;
    myFacesSameOriented : Boolean;
    
    myTol1,myTol2 : Real;
    
end Hctxff2d from TopOpeBRep;
