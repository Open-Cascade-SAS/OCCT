-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class UniformSurfaceAndRationalBSplineSurface from StepGeom 

inherits BSplineSurface from StepGeom 


	--- This classe is an implementation of EXPRESS
	--  ANDOR Subtype Declaration.
uses

	UniformSurface from StepGeom, 
	RationalBSplineSurface from StepGeom, 
	HAsciiString from TCollection, 
	Integer from Standard, 
	HArray2OfCartesianPoint from StepGeom, 
	BSplineSurfaceForm from StepGeom, 
	Logical from StepData, 
	HArray2OfReal from TColStd, 
	Real from Standard
is

	Create returns mutable UniformSurfaceAndRationalBSplineSurface;
	---Purpose: Returns a UniformSurfaceAndRationalBSplineSurface


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aUDegree : Integer from Standard;
	      aVDegree : Integer from Standard;
	      aControlPointsList : mutable HArray2OfCartesianPoint from StepGeom;
	      aSurfaceForm : BSplineSurfaceForm from StepGeom;
	      aUClosed : Logical from StepData;
	      aVClosed : Logical from StepData;
	      aSelfIntersect : Logical from StepData) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aUDegree : Integer from Standard;
	      aVDegree : Integer from Standard;
	      aControlPointsList : mutable HArray2OfCartesianPoint from StepGeom;
	      aSurfaceForm : BSplineSurfaceForm from StepGeom;
	      aUClosed : Logical from StepData;
	      aVClosed : Logical from StepData;
	      aSelfIntersect : Logical from StepData;
	      aUniformSurface : mutable UniformSurface from StepGeom;
	      aRationalBSplineSurface : mutable RationalBSplineSurface from StepGeom) is virtual;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aUDegree : Integer from Standard;
	      aVDegree : Integer from Standard;
	      aControlPointsList : mutable HArray2OfCartesianPoint from StepGeom;
	      aSurfaceForm : BSplineSurfaceForm from StepGeom;
	      aUClosed : Logical from StepData;
	      aVClosed : Logical from StepData;
	      aSelfIntersect : Logical from StepData;
	      aWeightsData : mutable HArray2OfReal from TColStd) is virtual;

	-- Specific Methods for Field Data Access --

	SetUniformSurface(me : mutable; aUniformSurface : mutable UniformSurface);
	UniformSurface (me) returns mutable UniformSurface;
	SetRationalBSplineSurface(me : mutable; aRationalBSplineSurface : mutable RationalBSplineSurface);
	RationalBSplineSurface (me) returns mutable RationalBSplineSurface;

	-- Specific Methods for ANDOR Field Data Access --

	SetWeightsData(me : mutable; aWeightsData : mutable HArray2OfReal);
	WeightsData (me) returns mutable HArray2OfReal;
	WeightsDataValue (me; num1 : Integer;  num2 : Integer) returns Real;
	NbWeightsDataI (me) returns Integer;
	NbWeightsDataJ (me) returns Integer;

	-- Specific Methods for ANDOR Field Data Access --


fields

	uniformSurface : UniformSurface from StepGeom;
	rationalBSplineSurface : RationalBSplineSurface from StepGeom;

end UniformSurfaceAndRationalBSplineSurface;
