-- Created on: 1991-05-14
-- Created by: Laurent Painnot
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.





class BracketedRoot from math
     	---Purpose: This class implements the Brent method to find the root of a function
     	-- located within two bounds. No knowledge of the derivative is required.

uses Matrix from math, 
     Vector from math, 
     Function from math,
     OStream from Standard

raises NotDone

is

    Create(F: in out Function;
    	   Bound1, Bound2, Tolerance: Real;
	   NbIterations: Integer = 100; ZEPS : Real =1.0e-12)
	---Purpose:   
    	-- The Brent method is used to find the root of the function F between 
    	-- the bounds Bound1 and Bound2 on the function F.
    	-- If F(Bound1)*F(Bound2) >0 the Brent method fails.  
    	-- The tolerance required for the root is given by Tolerance.
    	-- The solution is found when :
    	--    abs(Xi - Xi-1) <= Tolerance;
    	-- The maximum number of iterations allowed is given by NbIterations.

    returns BracketedRoot;
    
    IsDone(me)
    	---Purpose: Returns true if the computations are successful, otherwise returns false.
    	---C++: inline
    returns Boolean
    is static;


    Root(me)
        ---Purpose: returns the value of the root.
        -- Exception NotDone is raised if the minimum was not found.
     	---C++: inline
    returns Real
    raises NotDone
    is static;
    
    
    Value(me)
        ---Purpose: returns the value of the function at the root.
        -- Exception NotDone is raised if the minimum was not found.
      	---C++: inline
    returns Real
    raises NotDone
    is static;
    
    NbIterations(me)
        ---Purpose: returns the number of iterations really done during the
        -- computation of the Root.
        -- Exception NotDone is raised if the minimum was not found.
    	---C++: inline

    returns Integer
    raises NotDone
    is static;
    

    Dump(me; o: in out OStream)
	---Purpose: Prints on the stream o information on the current state 
    	--          of the object.

    is static;



fields

Done:      Boolean;
TheRoot:   Real;
TheError:  Real;
NbIter:    Integer;

end BracketedRoot;
