-- Created on: 1991-04-24
-- Created by: Arnaud BOUZY
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



package Draw 

	---Purpose: MAQUETTE DESSIN MODELISATION

uses OSD, MMgt, TCollection, TColStd, gp, Message

is
    exception Failure inherits Failure from Standard; 
     
    enumeration ColorKind is blanc,                 
    	    	    	    --white in english
    	    	    	     rouge,
                            --red in english
                             vert,
    	    	    	    --green in english
    	    	    	      bleu,
    	    	    	    --blue in english 
    	    	    	      cyan,
			    -- same in english
               	      	      or,
    	    	    	    --gold in english 
    	    	    	      magenta,
    	    	    	    --same in english 
    	    	    	      marron,
			    --brown in english
    	    	    	      orange,
    	    	    	    --same in english 
    	    	    	      rose,
			    --pink in english 
                     	      saumon,
    	    	    	    --salmon in english 
    	    	    	      violet,
			    --same in english 
                              jaune,
    	    	    	    --yellow in english 
    	    	    	      kaki,
                            --DarkOliveGreen in english 
                              corail;
			    --Coral in english 
		     
    enumeration MarkerShape is
    	Square, Losange, X, Plus, Circle, CircleZoom;
	
	---Purpose: Circle is not sensible to zoom, like 
	--          other MarkerShape, contrarily to CircleZoom
	


    deferred class Drawable3D;
    
    deferred class Drawable2D;
    
    class Color;
    
    class Display;
    
    class Segment3D;
    
    class Segment2D;
    
    class Marker3D;
    
    class Marker2D;
    
    class Axis3D;
    
    class Axis2D;
    
    class Text3D;
    
    class Text2D;
    
    class Circle3D;
    
    class Circle2D;
    
    class Number;
    
    class Chronometer;
    
    class Grid;
    
    class Box;
	---Purpose: a 3d box
    
    class SequenceOfDrawable3D instantiates 
    	Sequence from TCollection (Drawable3D);
	
    class ProgressIndicator;

    imported PInterp;
	---Purpose: typedef Tcl_Interp * Draw_PInterp;
    
    primitive CommandFunction;
	---Purpose: typedef Standard_Integer (*Draw_CommandFunction)
	--          (Draw_Interpretor&, Standard_Integer, char**)
    
    class Interpretor;
	---Purpose: Encapsulate the Tcl interpretor to add commands.

    class Printer;
	---Purpose: Implements a printer class to connect Message_Messenger 
	--          tool to Draw_Interpretor output.

    class VMap instantiates
      DataMap from TCollection(Integer,
    	    	    	       Drawable3D from Draw,
                               MapIntegerHasher from TColStd);    
        
    private class MapOfFunctions instantiates DataMap from TCollection(AsciiString from TCollection ,Function from OSD, AsciiString from TCollection);

    class MapOfAsciiString instantiates IndexedMap from TCollection(AsciiString from TCollection,AsciiString from TCollection); 
     
    Load(theDI: out Interpretor from Draw; theKey, theResourceFileName: AsciiString from TCollection)  
--    returns Transient from Standard
    raises Failure  from Draw;      
     
    Load(theDI: out Interpretor from Draw;
         theKey, theResourceFileName: AsciiString from TCollection;
         theDefaultsDirectory, theUserDefaultsDirectory: in out AsciiString from TCollection;
         Verbose :  Boolean from Standard = Standard_False)  
    raises Failure  from Draw;      

    --
    --  methods to handle variables
    --  
    
    Set(Name : CString;  
    	D : Drawable3D from Draw; 
        Disp : Boolean from Standard);
       ---Purpose: Sets a variable. Display it if <Disp> is true.
    
    Set(Name : CString;  
    	D : Drawable3D from Draw);
	---Purpose: Sets a    variable,  a  null   handle    clear the
	--          vartiable. Automatic display is context driven.
	
    Set(Name : CString;  
    	val : Real);
	---Purpose: Sets a numeric variable.
    
    Get(Name : in out CString;  
    	Complain : Boolean = Standard_True)
    	returns Drawable3D from Draw;
	---Purpose: Returns a variable  value.  Null if  the  variable
	--          does not exist, a warning  is printed if  Complain
	--          is True.
	--          
	--          The name "."   does a graphic  selection.   If the
	--          selection is a variable <Name> is overwritten with
	--          the name of the variable.
	
    Get(Name : CString;  
    	val : out Real)  
    	returns Boolean;
	---Purpose: Gets a   numeric  variable. Returns  True   if the
	--          variable exist.

    Set(Name : CString; val : CString);
	---Purpose: Sets a TCL sting variable
	
    Atof(Name : CString) returns Real;
	---Purpose: Search a  numeric  variable.  If none found converts
	--          the string to a real.
    
    Atoi(Name : CString) returns Integer;
	---Purpose: Search a  numeric  variable.  If none found converts
	--          the string to an integer.
    
    
    LastPick(view,X,Y,button : out Integer);
	---Purpose: Returns last graphic selection description.
	
    Repaint;
	---Purpose: Asks to repaint the screen after the current command.
	
    SetProgressBar(thePI: ProgressIndicator from Draw);
        ---Purpose: sets progress indicator
	
    GetProgressBar returns ProgressIndicator from Draw;
        ---Purpose: gets progress indicator


    --
    --	Draw Commands
    --		

    Commands(I : in out Interpretor from Draw);
	---Purpose: Defines all Draw commands

    BasicCommands(I : in out Interpretor from Draw);
	---Purpose: Defines Draw basic commands

    VariableCommands(I : in out Interpretor from Draw);
	---Purpose: Defines Draw variables handling commands.

    GraphicCommands(I : in out Interpretor from Draw);
	---Purpose: Defines Draw variables handling commands.

    PloadCommands(I : in out Interpretor from Draw);
	---Purpose: Defines Loads Draw plugins commands.

    UnitCommands(I : in out Interpretor from Draw);
	---Purpose: Defines Draw unit commands

end Draw;
