-- Created on: 2000-08-21
-- Created by: Andrey BETENEV
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Context from ShapeProcess inherits TShared from MMgt

    ---Purpose: Provides convenient interface to resource file
    --          Allows to load resource file and get values of
    --          attributes starting from some scope, for example
    --          if scope is defined as "ToV4" and requested parameter
    --          is "exec.op", value of "ToV4.exec.op" parameter from
    --          the resource file will be returned

uses

    Manager                 from Resource,
    AsciiString             from TCollection,
    HSequenceOfHAsciiString from TColStd,
    Messenger               from Message,
    ProgressIndicator       from Message

is

    Create;
    	---Purpose: Creates an empty tool

    Create (file: CString; scope: CString = "");
    	---Purpose: Creates a new tool and initialises by name of
	--          resource file and (if specified) starting scope
	--          Calls method Init()

    Init (me: mutable; file: CString; scope: CString = "")
    returns Boolean;
    	---Purpose: Initialises a tool by loading resource file and 
        --          (if specified) sets starting scope
	--          Returns False if resource file not found

    LoadResourceManager(me: mutable; file: CString) returns Manager from Resource;
    	---Purpose: Loading Resource_Manager object if this object not
	--          equal internal static Resource_Manager object or
	--          internal static Resource_Manager object is null

    ResourceManager (me) returns Manager from Resource;
    	---Purpose: Returns internal Resource_Manager object
	---C++: return const &

    SetScope (me: mutable; scope: CString);
    	---Purpose: Set a new (sub)scope

    UnSetScope (me: mutable);
    	---Purpose: Go out of current scope

    IsParamSet (me; param: CString) returns Boolean;
    	---Purpose: Returns True if parameter is defined in the resource file

    GetReal    (me; param: CString; val: out Real   ) returns Boolean;
    GetInteger (me; param: CString; val: out Integer) returns Boolean;
    GetBoolean (me; param: CString; val: out Boolean) returns Boolean;
    GetString  (me; param: CString; val: out AsciiString from TCollection) returns Boolean;
    	---Purpose: Get value of parameter as being of specific type
	--          Returns False if parameter is not defined or has a wrong type

    RealVal    (me; param: CString; def: Real   ) returns Real;
    IntegerVal (me; param: CString; def: Integer) returns Integer;
    BooleanVal (me; param: CString; def: Boolean) returns Boolean;
    StringVal  (me; param: CString; def: CString) returns CString;
    	---Purpose: Get value of parameter as being of specific type
	--          If parameter is not defined or does not have expected
        --          type, returns default value as specified

    SetMessenger (me: mutable; messenger: Messenger from Message);
    ---Purpose : Sets Messenger used for outputting messages.

    Messenger (me) returns Messenger from Message;
    ---Purpose : Returns Messenger used for outputting messages.
    
    SetProgress (me: mutable; theProgress: ProgressIndicator from Message);
    ---Purpose : Sets Progress Indicator.

    Progress (me) returns ProgressIndicator from Message;
    ---Purpose : Returns Progress Indicator.

    SetTraceLevel (me: mutable; tracelev: Integer);
    ---Purpose : Sets trace level used for outputting messages
    --           - 0: no trace at all
    --           - 1: errors
    --           - 2: errors and warnings
    --           - 3: all messages
    --           Default is 1 : Errors traced

    TraceLevel (me) returns Integer;
    ---Purpose : Returns trace level used for outputting messages.

fields

    myRC:        Manager from Resource;
    myScope:     HSequenceOfHAsciiString from TColStd;
    myMessenger: Messenger from Message;
    myProgress:  ProgressIndicator from Message;
    myTraceLev:  Integer;

end Context;
