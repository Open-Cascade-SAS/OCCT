-- Created on: 1993-06-14
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class BuilderON from TopOpeBRepBuild

uses

    PBuilder from TopOpeBRepBuild,
    PGTopo from TopOpeBRepBuild,
    PWireEdgeSet from TopOpeBRepBuild,
    ListOfShape from TopTools,
    Shape from TopoDS,
    Interference from TopOpeBRepDS,
    ListOfInterference from TopOpeBRepDS,
    Plos from TopOpeBRepTool

is
    -- BuilderON3d
    --------------
    Create returns BuilderON;
    Create(PB:PBuilder;F:Shape;PG:PGTopo;PLSclass:Plos;PWES:PWireEdgeSet) returns BuilderON;
    Perform(me:in out;PB:PBuilder;F:Shape;PG:PGTopo;PLSclass:Plos;PWES:PWireEdgeSet) is static;

    -- private
    GFillONCheckI(me;I:Interference) returns Boolean;
    GFillONPartsWES1(me:in out;I:Interference);
    GFillONPartsWES2(me:in out;I:Interference;EspON:Shape);


    -- BuilderON2d
    --------------
    Perform2d(me:in out;PB:PBuilder;F:Shape;PG:PGTopo;PLSclass:Plos;PWES:PWireEdgeSet) is static;
    
    -- private
    GFillONParts2dWES2(me:in out;I:Interference;EspON:Shape);
    
fields

    myPB : PBuilder from TopOpeBRepBuild;
    myPG : PGTopo from TopOpeBRepBuild;
    myPLSclass : Plos from TopOpeBRepTool;
    myPWES : PWireEdgeSet from TopOpeBRepBuild;
    myFace : Shape from TopoDS;
    
    myFEI : ListOfInterference from TopOpeBRepDS; --BuilderON2d 
    
end BuilderON from TopOpeBRepBuild;
