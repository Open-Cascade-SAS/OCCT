-- Created on: 1997-02-05
-- Created by: Alexander BRIVIN and Dmitry TARASOV
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Coordinate3 from Vrml inherits  TShared  from  MMgt

	---Purpose: defines a Coordinate3 node of VRML specifying
	--          properties of geometry and its appearance. 
    	--  This node defines a set of 3D coordinates to be used by a subsequent IndexedFaceSet,  
    	--  IndexedLineSet, or PointSet node. This node does not produce a visible result  
    	--  during rendering; it simply replaces the current coordinates in the rendering  
    	--  state for subsequent nodes to use. 
uses
 
     HArray1OfVec  from  TColgp 

is
    Create ( aPoint : HArray1OfVec  from  TColgp )
    	returns Coordinate3 from Vrml; 
     
    Create  returns Coordinate3 from Vrml;
    
    SetPoint ( me  :  mutable; aPoint : HArray1OfVec  from  TColgp );
    Point ( me )  returns  HArray1OfVec  from  TColgp; 
    
    Print  ( me;  anOStream: in out OStream from Standard) returns OStream from Standard;
    ---C++:  return  & 

fields

    myPoint  : HArray1OfVec  from  TColgp;  -- Coordinate point(s)

end Coordinate3;
