-- Created on: 1992-11-19
-- Created by: Remi LEQUETTE
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Edge from BRepClass 

	---Purpose: This class  is used to send  the  description of an
	--          Edge to the classifier. It  contains  an Edge and a
	--          Face. So the PCurve of the Edge can be found.

uses
    Edge from TopoDS,
    Face from TopoDS

is
    Create returns Edge from BRepClass;
    
    Create (E : Edge from TopoDS; F : Face from TopoDS)
    returns Edge from BRepClass;

    Edge(me : in out) returns Edge from TopoDS
	---C++: inline
	---C++: return &
	---C++: alias "const TopoDS_Edge& Edge() const;"
    is static;
    
    Face(me : in out) returns Face from TopoDS
	---C++: inline
	---C++: return &
	---C++: alias "const TopoDS_Face& Face() const;"
    is static;

fields
    myEdge : Edge from TopoDS;
    myFace : Face from TopoDS;

end Edge;
