-- Created on: 1994-06-01
-- Created by: Christian CAILLET
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class RebuildDrawings  from IGESSelect  inherits ModelModifier from IGESSelect

    ---Purpose : Rebuilds Drawings which were bypassed to produce new models.
    --           If a set of entities, all put into a same IGESModel, were
    --           attached to a same Drawing in the starting Model, this Modifier
    --           rebuilds the original Drawing, but only with the transferred
    --           entities. This includes that all its views are kept too, but
    --           empty; and annotations are not kept. Drawing Name is renewed.
    --           
    --           If the Input Selection is present, tries to rebuild Drawings
    --           only for the selected entities. Else, tries to rebuild
    --           Drawings for all the transferred entities.

uses AsciiString from TCollection,
     IGESModel, CopyTool, ContextModif

is

    Create returns mutable RebuildDrawings;
    ---Purpose : Creates an RebuildDrawings, which uses the system Date

    Performing (me; ctx : in out ContextModif;
    	        target  : mutable IGESModel;
                TC      : in out CopyTool);
    ---Purpose : Specific action : Rebuilds the original Drawings

    Label (me) returns AsciiString from TCollection;
    ---Purpose : Returns a text which is
    --           "Rebuild Drawings"

end RebuildDrawings;
