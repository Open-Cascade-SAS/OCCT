-- Created on: 1993-03-23
-- Created by: BBL,JLF
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Modified:    DCB (20-OCT-98)
--              Define ToImage()/FromName() as deferred.

deferred class AlienUserImage from AlienImage inherits AlienImage

        ---Version: 0.0

        ---Purpose: This class defines an Alien user image.
        -- Alien Image is X11 .xwd image or SGI .rgb image for examples

        ---Keywords:
        ---Warning:
        ---References:

uses
        Image   from Image,
        File    from OSD

raises
        TypeMismatch    from Standard

is
        Initialize ;

        Read ( me : in out mutable ; afile : in out File from OSD )
          returns Boolean from Standard is deferred;
        ---Level: Public
        ---Purpose: Read content of a  UserAlienImage object from a file .
        --         Returns True if sucess .

        Read ( me : in out mutable ; afile : in CString from Standard )
          returns Boolean from Standard ;
        ---Level: Public
        ---Purpose: Read content of a UserAlienImage object from a file .
        --          Returns True if file is a AlienImage file .

        Write ( me : in immutable ; afile : in out File from OSD )
          returns Boolean from Standard is deferred ;
        ---Level: Public
        ---Purpose: Write content of a UserAlienImage object to a file .

        Write ( me : in immutable ; afile : in CString from Standard )
          returns Boolean from Standard ;
        ---Level: Public
        ---Purpose: Write content of a UserAlienImage object to a file .

        ToImage ( me : in  immutable )
        returns mutable Image from Image 
        raises TypeMismatch from Standard
        is deferred;
        ---Level: Public
        ---Purpose : convert a AidaAlienData object to a Image object.

        FromImage ( me : in out mutable ; anImage : in Image from Image )
        raises TypeMismatch from Standard
        is deferred;
        ---Level: Public
        ---Purpose : convert a Image object to a AidaAlienData object.

end AlienUserImage;
 
