-- Created on: 1993-06-17
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class HDataStructure from TopOpeBRepDS inherits TShared from MMgt

uses

    AsciiString                      from TCollection,
    Orientation                      from TopAbs,
    ShapeEnum                        from TopAbs,
    ListIteratorOfListOfShape        from TopTools,
    OStream                          from Standard,
    Shape                            from TopoDS,
    SurfaceIterator                  from TopOpeBRepDS,
    CurveIterator                    from TopOpeBRepDS,
    PointIterator                    from TopOpeBRepDS,
    DataStructure                    from TopOpeBRepDS,
    Surface                          from TopOpeBRepDS,
    Curve                            from TopOpeBRepDS,
    Point                            from TopOpeBRepDS,
    Kind                             from TopOpeBRepDS,
    Config                           from TopOpeBRepDS,    	
    Check                            from TopOpeBRepDS,
    Interference                     from TopOpeBRepDS,
    ListOfInterference               from TopOpeBRepDS,
    ListIteratorOfListOfInterference from TopOpeBRepDS
    
is

    Create returns mutable HDataStructure from TopOpeBRepDS;
    
    AddAncestors(me : mutable; S : Shape from TopoDS);
    
    AddAncestors(me : mutable; S  : Shape from TopoDS;
    	    	               T1,T2 : ShapeEnum from TopAbs)
    ---Purpose: Update  the data structure with  shapes of type T1
    --          containing a subshape of type T2 which is stored
    --          in the DS.
    --          Used by the previous one.
    is static;

    Complete(me : mutable) 
    ---Purpose: perform post processing of the DS.
    is static;

    ChkIntg(me : mutable)
    ---Purpose: Check the integrity of the DS
    is static;
    
    DS(me) returns DataStructure from TopOpeBRepDS
	---C++: return const &
    is static;

    ChangeDS(me : mutable) returns DataStructure from TopOpeBRepDS
	---C++: return &
    is static;

    --
    --   The new geometries
    --   
    
    NbSurfaces(me) returns Integer
    is static;
    
    NbCurves(me) returns Integer
    is static;
    
    NbPoints(me) returns Integer
    is static;
    
    Surface(me; I : Integer) returns Surface from TopOpeBRepDS
    ---Purpose: Returns the surface of index <I>.
	---C++: return const &
    is static;
    
    SurfaceCurves(me; I : Integer) returns CurveIterator from TopOpeBRepDS
    ---Purpose: Returns an iterator  on the curves on  the surface
	--          <I>. 
    is static;
    
    Curve(me; I : Integer) returns Curve from TopOpeBRepDS
    ---Purpose: Returns the Curve of index <I>.
	---C++: return const &
    is static;

    ChangeCurve(me : mutable ; I : Integer) returns Curve from TopOpeBRepDS
    ---Purpose: Returns the Curve of index <I>.
	--          
	---C++: return &
    is static;

    CurvePoints(me; I : Integer) returns PointIterator from TopOpeBRepDS
    ---Purpose: Returns an iterator   on the points on  the  curve
	--          <I>.
    is static;
    
    Point(me; I : Integer) returns Point from TopOpeBRepDS
    ---Purpose: Returns the point of index <I>.
	---C++: return const &
    is static;
    
    
   --
   --   The topologies
   --   

   NbShapes(me) returns Integer
   is static; 

   Shape(me; I : Integer;
    	    	 FindKeep : Boolean = Standard_True)
    returns Shape from TopoDS
   ---Purpose: Returns the shape of index <I> in the DS
   ---C++: return const &
   is static;

   Shape(me; S : Shape from TopoDS;
    	    	 FindKeep : Boolean = Standard_True)
    returns Integer from Standard
   ---Purpose: Returns the index of shape <S> in the DS
       --          returns 0 if <S> is not in the DS
    is static;
    
   --
   --   Geometry attached to topology
   --   
   
    HasGeometry(me; S : Shape from TopoDS) returns Boolean
    ---Purpose: Returns True if <S> has new geometries.
    is static;
   
    HasShape(me; S : Shape from TopoDS;
    	    	 FindKeep : Boolean = Standard_True)
    returns Boolean
    ---Purpose: Returns True if <S> has new geometries (SOLID,FACE,EDGE)
	--          or if <S> (SHELL,WIRE) has sub-shape (FACE,EDGE)
	--          with new geometries
    is static;

    HasSameDomain(me; S : Shape from TopoDS;
    	    	      FindKeep : Boolean = Standard_True)
    ---Purpose: Returns True if <S> share a geometrical domain with
	--          some other shapes.
    returns Boolean is static;

    SameDomain(me; S : Shape from TopoDS) 
    returns ListIteratorOfListOfShape from TopTools
    ---Purpose: Returns an iterator on the SameDomain shapes attached
	--          to the shape <S>.
    is static;
   
    SameDomainOrientation(me; S : Shape from TopoDS) 
    returns Config from TopOpeBRepDS
    ---Purpose: Returns orientation of shape <S> compared with its 
	--          reference shape
    is static;
   
    SameDomainReference(me; S : Shape from TopoDS) 
    returns Integer from Standard
    ---Purpose: Returns orientation of shape <S> compared with its 
	--          reference shape
    is static;
   
    SolidSurfaces(me; S : Shape from TopoDS) 
    returns SurfaceIterator from TopOpeBRepDS
    ---Purpose: Returns an iterator on the  surfaces attached to the
	--          solid <S>.
    is static;
    
    SolidSurfaces(me; I : Integer from Standard) 
    returns SurfaceIterator from TopOpeBRepDS
    ---Purpose: Returns an iterator on the  surfaces attached to the
	--          solid <I>.
    is static;
    
    FaceCurves(me; F : Shape from TopoDS) 
    returns CurveIterator from TopOpeBRepDS
    ---Purpose: Returns an iterator on the  curves attached to the
	--          face <F>.
    is static;
    
    FaceCurves(me; I : Integer from Standard) 
    returns CurveIterator from TopOpeBRepDS
    ---Purpose: Returns an iterator on the  curves attached to the
	--          face <I>.
    is static;
    
    EdgePoints(me; E : Shape from TopoDS) 
    returns PointIterator from TopOpeBRepDS
    ---Purpose: Returns an iterator on the points  attached to the
	--          edge <E>.
    is static;

    MakeCurve(me : mutable; 
     	      C1 : Curve from TopOpeBRepDS;
    	      C2 : in out Curve from TopOpeBRepDS)
    returns Integer from Standard
    is static;

    RemoveCurve(me : mutable; iC : Integer from Standard)
    is static;
    
    RemoveShape(me : mutable; iS : Integer from Standard)
    is static;
    
    NbGeometry(me; K : Kind from TopOpeBRepDS) 
    returns Integer from Standard is static;

    NbTopology(me; K : Kind from TopOpeBRepDS) 
    returns Integer from Standard is static;

    NbTopology(me)
    returns Integer from Standard is static;

    EdgesSameParameter(me)
    returns Boolean from Standard is static;
    ---Purpose: returns True if all the edges stored as shapes in the DS
    --          are SameParameter, otherwise False.
    
    SortOnParameter(me; L1 : ListOfInterference from TopOpeBRepDS;  
	                L2 : out ListOfInterference from TopOpeBRepDS)
    is static;

    SortOnParameter(me; L : in out ListOfInterference from TopOpeBRepDS)
    is static;

    MinMaxOnParameter(me; L : ListOfInterference from TopOpeBRepDS;
    	                  Min,Max : out Real from Standard)
    is static;

    ScanInterfList(me; 
    	      IT  : in out ListIteratorOfListOfInterference from TopOpeBRepDS; 
    	      PDS : Point from TopOpeBRepDS)
    ---Purpose: 
    	-- Search, among a list of interferences accessed by the iterator
    	-- <IT>, a geometry <G> whose 3D point is identical to the 3D point
    	-- of the TheDSPoint <PDS>.
    	-- returns True if such an interference has been found, False else.
    	-- if True, iterator It points (by the Value() method) on the first 
    	-- interference accessing an identical 3D point.
    returns Boolean from Standard
    is static;
    
    GetGeometry(me; 
    	    	IT  : in out ListIteratorOfListOfInterference from TopOpeBRepDS;
    	    	PDS : Point from TopOpeBRepDS;
		G   : out Integer from Standard;
		K   : out Kind from TopOpeBRepDS)
    ---Purpose:
    	-- Get the geometry of a DS point <PDS>.
    	-- Search for it with ScanInterfList (previous method).
    	-- if found, set <G,K> to the geometry,kind of the interference found.
    	-- returns the value of ScanInterfList().
    returns Boolean from Standard
    is static;
        
    StoreInterference(me : mutable; 
    	    	      I  : Interference from TopOpeBRepDS;
      	    	      LI : in out ListOfInterference from TopOpeBRepDS;
    	    	      str : AsciiString from TCollection = "");
    ---Purpose: 
    -- Add interference <I> to list <LI>.

    StoreInterference(me : mutable; I : Interference from TopOpeBRepDS;
      	        	            S : Shape from TopoDS;
    	    	                    str : AsciiString from TCollection = "");
    ---Purpose: 
    -- Add interference <I> to list of interference of shape <S>.

    StoreInterference(me : mutable; I  : Interference from TopOpeBRepDS;
      	        	            IS : Integer;
    	    	                    str : AsciiString from TCollection = "");
    ---Purpose: 
    -- Add interference <I> to list of interference of shape <IS>.

    StoreInterferences(me : mutable; LI : ListOfInterference from TopOpeBRepDS;
      	        	            S : Shape from TopoDS;
    	    	                    str : AsciiString from TCollection = "");				    
    StoreInterferences(me : mutable; LI  : ListOfInterference from TopOpeBRepDS;
      	        	            IS : Integer;
    	    	                    str : AsciiString from TCollection = "");
    ClearStoreInterferences(me : mutable; LI : ListOfInterference from TopOpeBRepDS;
      	        	            S : Shape from TopoDS;
    	    	                    str : AsciiString from TCollection = "");
				    
    ClearStoreInterferences(me : mutable; LI  : ListOfInterference from TopOpeBRepDS;
      	        	            IS : Integer;
    	    	                    str : AsciiString from TCollection = "");

fields
    
    myDS                 : DataStructure from TopOpeBRepDS;
    myEdgesSameParameter : Boolean from Standard;

    -- myAscii : to avoid bug WOK (incomplete hxx incomplete for HDatatStructure users)
    myAscii : AsciiString from TCollection;
    
end HDataStructure from TopOpeBRepDS;
