-- Created on: 1997-11-06
-- Created by: Roman BORISOV
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


private  class PrjResolve from ProjLib 

	---Purpose: 

uses     
    Pnt2d     from gp,
    Surface from Adaptor3d, 
    Curve  from  Adaptor3d, 
    SurfacePtr from Adaptor3d, 
    CurvePtr  from Adaptor3d

raises   
    	DomainError from Standard, 
	ConstructionError,
    	NotDone     from StdFail

is
    Create (C: Curve  from  Adaptor3d; S: Surface from Adaptor3d;  Fix: Integer)
    	returns PrjResolve 
    	raises  ConstructionError;
    	
     
    Perform(me:  in  out;  t,  U,  V:  Real;  Tol,  Inf,  Sup:  Pnt2d;  FTol:  Real  from  Standard  =  -1;  StrictInside:  Boolean  from  Standard  =  Standard_False) 
---Purpose: Calculates the ort from  C(t)  to  S  with a close point.
    	--          The close point is defined by the parameter values
    	--          U0 and V0.
    	--          The function F(u,v)=distance(S(u,v),C(t)) has an
    	--          extremum when gradient(F)=0. The algorithm searchs
    	--          a zero near the close point.
    	raises  DomainError;
	    	-- if U0,V0 are outside the definition ranges of the 
	    	-- surface.
     
    
    IsDone (me)  returns Boolean
    	---Purpose: Returns True if the distance is found.
    	is static;
 
    Solution (me) returns Pnt2d  from  gp
    	---Purpose: Returns the point of the extremum distance.
    	raises  NotDone from StdFail
	    	-- if IsDone(me)=False.
    	is static;

fields
     
    myCurve    :  CurvePtr    from  Adaptor3d; 
    mySurface  :  SurfacePtr  from  Adaptor3d;	     
    myDone     :  Boolean     from  Standard;
    mySolution :  Pnt2d       from  gp; 
    myFix      :  Integer     from  Standard; 
     
end PrjResolve;
