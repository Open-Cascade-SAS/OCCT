-- Created on: 1992-08-28
-- Created by: Remi LEQUETTE
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package GeomTools 

	---Purpose: The GeomTools package provides  utilities for Geometry.
	--          
	--          *  SurfaceSet,  CurveSet, Curve2dSet  : Tools used
	--          for dumping, writing and reading.
	--          
	--          * Methods to dump, write, read curves and surfaces.

uses
    Geom,
    Geom2d,
    TColStd,
    Message

is

    class UndefinedTypeHandler;
    --
    --  Dump, Write, Read tools
    
    class SurfaceSet;
	---Purpose: A set of Surfaces from Geom.
    	
    class CurveSet;
	---Purpose: A set of Curves from Geom.
    	
    class Curve2dSet;
	---Purpose: A set of Curves from Geom2d.
    	
    --
    --     Methods
    --     
    
    Dump(S : Surface from Geom; OS : in out OStream);
	  ---Purpose: Dumps the surface on the stream.

    Write(S : Surface from Geom; OS : in out OStream);
	  ---Purpose: Writes the surface on the stream.

    Read(S : in out Surface from Geom; IS : in out IStream); 
	  ---Purpose: Reads the surface from the stream.


    Dump(C : Curve from Geom; OS : in out OStream);
	  ---Purpose: Dumps the Curve on the stream.

    Write(C : Curve from Geom; OS : in out OStream);
	  ---Purpose: Writes the Curve on the stream.

    Read(C : in out Curve from Geom; IS : in out IStream); 
	  ---Purpose: Reads the Curve from the stream.


    Dump(C : Curve from Geom2d; OS : in out OStream);
	  ---Purpose: Dumps the Curve on the stream.

    Write(C : Curve from Geom2d; OS : in out OStream);
	  ---Purpose: Writes the Curve on the stream.

    Read(C : in out Curve from Geom2d; IS : in out IStream); 
	  ---Purpose: Reads the Curve from the stream.
	  
    SetUndefinedTypeHandler(aHandler: UndefinedTypeHandler from GeomTools);
    
    GetUndefinedTypeHandler returns UndefinedTypeHandler from GeomTools;

end GeomTools;


