-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class BoxDomain from StepShape 

inherits TShared from MMgt

uses

	CartesianPoint from StepGeom, 
	Real from Standard
is

	Create returns mutable BoxDomain;
	---Purpose: Returns a BoxDomain

	Init (me : mutable;
	      aCorner : mutable CartesianPoint from StepGeom;
	      aXlength : Real from Standard;
	      aYlength : Real from Standard;
	      aZlength : Real from Standard) is virtual;

	-- Specific Methods for Field Data Access --

	SetCorner(me : mutable; aCorner : mutable CartesianPoint);
	Corner (me) returns mutable CartesianPoint;
	SetXlength(me : mutable; aXlength : Real);
	Xlength (me) returns Real;
	SetYlength(me : mutable; aYlength : Real);
	Ylength (me) returns Real;
	SetZlength(me : mutable; aZlength : Real);
	Zlength (me) returns Real;

fields

	corner : CartesianPoint from StepGeom;
	xlength : Real from Standard;
	ylength : Real from Standard;
	zlength : Real from Standard;

end BoxDomain;
