-- Created on: 1991-03-22
-- Created by: Philippe DAUTRY
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package GccInt

	---Purpose: This package implements the services needed by the 
	--          toolkit Gcc to use curves other than lines or circles.
	--          This package is also used for intersections and 
	--          bisecting curves.

uses gp,
     MMgt,
     Standard

is

enumeration IType is Lin, Cir, Ell, Par, Hpr, Pnt;

deferred class Bisec;

class BCirc;

class BElips;

class BLine;

class BParab;

class BPoint;

class BHyper;

end GccInt;
