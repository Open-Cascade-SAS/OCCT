-- Created on: 2000-11-23
-- Created by: Michael KLOKOV
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Curve from IntTools
      ---Purpose: class is a container of
      --          one 3d curve
      --          two 2d curves

uses
    Curve from Geom,
    Curve from Geom2d,
    Pnt  from gp, 
    CurveType from GeomAbs
is
    Create  
    	returns Curve from IntTools;
	---Purpose:
	--- Empty constructor
	---

    Create(Curve3d: Curve from Geom;  
    	   FirstCurve2d : Curve from Geom2d;
    	   SecondCurve2d: Curve from Geom2d)
    	returns Curve from IntTools;
	---Purpose:
	--- Initializes me by a 3d curve
	--- and two 2d curves
	---

    SetCurves(me: in out;  
    	      Curve3d: Curve from Geom;  
    	      FirstCurve2d  : Curve from Geom2d;
    	      SecondCurve2d : Curve from Geom2d);
    	---Purpose:
	--- Modifier
	---
    
    SetCurve(me: in out;  
    	    	Curve3d: Curve from Geom);
    	---C++: inline
	---Purpose:
	--- Modifier
	---
    
    SetFirstCurve2d(me: in out;  
    	    	FirstCurve2d: Curve from Geom2d);
    	---C++: inline
	---Purpose:
	--- Modifier
	---
    
    SetSecondCurve2d(me: in out;  
    	    	SecondCurve2d: Curve from Geom2d);
    	---C++: inline
	---Purpose:
	--- Modifier
	---

    Curve(me)  
    	returns any Curve from Geom;
    	---C++: return const &
	---C++: inline
	---Purpose:
	--- Selector
	---
    
    FirstCurve2d(me)
    	returns any Curve from Geom2d;
    	---C++: return const &
	---C++: inline
	---Purpose:
	--- Selector
	---
	    
    SecondCurve2d(me)
    	returns any Curve from Geom2d;
    	---C++: return const &
	---C++: inline 
	---Purpose:
	--- Selector
	---
	
    HasBounds (me) 
    	returns Boolean from Standard;
	---Purpose:
	--- Returns true if 3d curve is BoundedCurve from Geom
	---

    Bounds    (me; aT1:out Real from Standard;    	  
                   aT2:out Real from Standard;    	  
		   aP1:out Pnt  from gp;     
		   aP2:out Pnt  from gp);
    	---Purpose:
	--- Returns boundary parameters
	--- and corresponded 3d point.
	---
	--  Warning:
	--- If HasBounds returns false
	--- the returned parameters are equal
	--- to zero.
	---

    D0        (me;  
    	       aT1:out Real from Standard; 
               aP1:out Pnt  from gp) 
    	returns Boolean from Standard;
	---Purpose:
	--- Computes 3d point corresponded to parameter aT1
	--- Returns true if given parameter aT1
	--- is inside the boundaries of the curve
	---
     
    Type  (me) 
    	returns CurveType from GeomAbs; 
	---Purpose:
	--- Returns the type of 3d curve
	---
 
fields

    my3dCurve : Curve from Geom;
    my2dCurve1: Curve from Geom2d;
    my2dCurve2: Curve from Geom2d;
    
end Curve from IntTools;
