-- Created on: 1990-12-17
-- Created by: Remi Lequette
-- Copyright (c) 1990-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Face from TopoDS inherits Shape from TopoDS

	---Purpose: Describes a face which
-- - references an underlying face with the potential to
--   be given a location and an orientation
-- - has a location for the underlying face, giving its
--   placement in the local coordinate system
-- - has an orientation for the underlying face, in terms
--   of its geometry (as opposed to orientation in relation to other shapes).

is
    Create returns Face from TopoDS;
    ---C++: inline
	---Purpose: Undefined Face.

end Face;
