-- File:        OrientedEdge.cdl
-- Created:     Mon Dec  4 12:02:28 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWOrientedEdge from RWStepShape

	---Purpose : Read & Write Module for OrientedEdge

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     OrientedEdge from StepShape,
     EntityIterator from Interface

is

	Create returns RWOrientedEdge;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable OrientedEdge from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : OrientedEdge from StepShape);

	Share(me; ent : OrientedEdge from StepShape; iter : in out EntityIterator);

end RWOrientedEdge;
