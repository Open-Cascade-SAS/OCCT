-- Created on: 1993-02-25
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class BlockBuilder from BOP
    	 
    ---Purpose: 
    ---  auxiliary class to storage and operate with data of  
    ---  connexity blocks inside the given ShapeSet 
    --- 
     
uses
    
    Shape     from TopoDS,  
     
    ShapeSet  from BOP,
    BlockIterator from BOP,

    SequenceOfInteger         from TColStd,
    DataMapOfIntegerInteger   from TColStd,
    IndexedMapOfOrientedShape from TopTools

is

    Create  
    	returns BlockBuilder;
    	---Purpose:  
    	--- Empty  Constructor 
    	---
    Create(SS : in out ShapeSet)  
    	returns BlockBuilder;
    	---Purpose:  
    	--- Create an  object for given ShapeSet  
    	---
    MakeBlock(me : in out;  
    	      SS : in out ShapeSet)  
    	is static;
    	---Purpose:   
    	--- Compute the set of connexity blocks of elements  
    	--- for of the ShapeSet SS
    -- 
    --	
    --   I t e r a t i o n   o n   b l o c k s made by MakeBlock
    -- 
    InitBlock(me : in out)  
    	is static; 

    MoreBlock(me)  
    	returns Boolean from Standard  
    	is static; 
	
    NextBlock(me : in out)  
    	is static;
    --
    -- I t e r a t i o n   o n  on shapes inside the current block 
    --
    BlockIterator(me)  
    	returns BlockIterator from  BOP   
    	is static;
    	--- Purpose:  
    	--- Returns the BlockIterator for the current block  .
    	---
    Element(me; BI : BlockIterator from  BOP)  
    	returns Shape from TopoDS  
    	is static; 
    	---C++: return const &
    	---Purpose:  
    	--- Returns the current element of <BI>.
    	---
    Element(me; I : Integer from Standard)  
    	returns Shape from TopoDS  
    	is static;
    	---C++: return const & 
    	---Purpose:  
    	--- Returns the current element with index  <I> .
    	---
    Element(me; S : Shape from TopoDS)  
    	returns Integer from Standard;
    	---Purpose:   
    	--- Returns the index of the current element .
    	---
    ElementIsValid(me; BI : BlockIterator)  
    	returns Boolean from Standard; 
    	---Purpose:   
    	--- Internal
    	---
    ElementIsValid(me; I : Integer from Standard)  
    	returns Boolean from Standard; 
    	---Purpose:   
    	--- Internal
    	---
    AddElement(me : in out; S : Shape from TopoDS)  
    	returns Integer from Standard;
    	---Purpose:   
    	--- Internal 
    	---
    SetValid(me : in out;  
    	     BI : BlockIterator from  BOP ;  
    	     IsValid : Boolean from Standard); 
    	---Purpose:   
    	--- Internal
    	---
    SetValid(me : in out;  
    	     I : Integer from Standard;  
    	     IsValid : Boolean from Standard);
    	---Purpose:   
    	--- Internal
    	---
    CurrentBlockIsRegular(me : in out)  
    	returns Boolean from Standard;
    	---Purpose:   
    	--- Returns TRUE if all elements inside the current block 
    	--- are biconnexial          
    	---
    
fields

    myOrientedShapeMapIsValid : DataMapOfIntegerInteger from TColStd;
    myOrientedShapeMap        : IndexedMapOfOrientedShape from TopTools;
    myBlocks                  : SequenceOfInteger from TColStd;
    myBlockIndex              : Integer from Standard;
    myIsDone                  : Boolean from Standard;
    myBlocksIsRegular         : SequenceOfInteger from TColStd;

end BlockBuilder;
