-- Created on: 1993-09-23
-- Created by: Jean Louis FRENKEL
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ShadedShape from StdPrs

inherits Root from Prs3d
  --- Purpose: unknown.

uses

  Presentation from Prs3d,
  Drawer       from Prs3d,
  Shape        from TopoDS,
  Pnt2d        from gp

is

  Add (myclass;
       thePresentation : Presentation from Prs3d;
       theShape        : Shape        from TopoDS;
       theDrawer       : Drawer       from Prs3d);
  ---Purpose: Shades <theShape>.

  Add (myclass;
       thePresentation : Presentation from Prs3d;
       theShape        : Shape        from TopoDS;
       theDrawer       : Drawer       from Prs3d;
       theHasTexels    : Boolean      from Standard;
       theUVOrigin     : Pnt2d        from gp;
       theUVRepeat     : Pnt2d        from gp;
       theUVScale      : Pnt2d        from gp);
  ---Purpose: Shades <theShape> with texture coordinates.

  Tessellate (myclass;
              theShape  : Shape  from TopoDS;
              theDrawer : Drawer from Prs3d);
  ---Purpose: Validates triangulation within the shape and performs tessellation if necessary.

end ShadedShape;
