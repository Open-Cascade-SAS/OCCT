-- File:        GeometricallyBoundedSurfaceShapeRepresentation.cdl
-- Created:     Mon Dec  4 12:02:27 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWGeometricallyBoundedSurfaceShapeRepresentation from RWStepShape

	---Purpose : Read & Write Module for GeometricallyBoundedSurfaceShapeRepresentation

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     GeometricallyBoundedSurfaceShapeRepresentation from StepShape,
     EntityIterator from Interface

is

	Create returns RWGeometricallyBoundedSurfaceShapeRepresentation;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable GeometricallyBoundedSurfaceShapeRepresentation from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : GeometricallyBoundedSurfaceShapeRepresentation from StepShape);

	Share(me; ent : GeometricallyBoundedSurfaceShapeRepresentation from StepShape; iter : in out EntityIterator);

end RWGeometricallyBoundedSurfaceShapeRepresentation;
