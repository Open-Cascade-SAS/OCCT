-- Created on: 1993-09-30
-- Created by: Isabelle GRIGNON
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class ShapeTool from BRepMesh 

	---Purpose: 

uses Shape from TopoDS,
     Face from TopoDS,
     Edge from TopoDS,
     Vertex from TopoDS,
     Explorer from TopExp,
     Pnt2d from gp,
     Pnt from gp,
     Box from Bnd,
     Curve from BRepAdaptor,
     Orientation from TopAbs,
     Triangulation from Poly,
     HArray1OfInteger from TColStd

raises NoSuchObject from Standard

is
    	Create  returns ShapeTool ;
	
	Init(me : in out ; S : Shape from TopoDS)
        ---C++: inline	
    	is static;
	
	MoreFace(me: in out ) returns Boolean from Standard
        ---C++: inline		
    	is static;
	
	NextFace(me : in out) 
        ---C++: inline		
    	is static;
	
    	CurrentFace( me : in out) returns Face from TopoDS
	---C++:return const &    	
        ---C++: inline		
      	is static;
	
	Init(me : in out ; F: Face from TopoDS)
        ---C++: inline		
    	is static;
	
	MoreEdge(me: in out ) returns Boolean from Standard
        ---C++: inline		
    	is static;
	
	NextEdge(me : in out) 
        ---C++: inline		
    	is static;
	
	CurrentEdge(me     : in out) 
	    ---C++: return const &
            ---C++: inline		
    	    returns Edge from TopoDS
    	is static;

	Init(me : in out ; E : Edge from TopoDS)
        ---C++: inline		
    	is static;
	
	MoreInternalVertex(me: in out ) returns Boolean from Standard

    	is static;
	
	NextInternalVertex(me : in out) 
        ---C++: inline		
    	is static;
	
	CurrentInternalVertex( me : in out) returns Vertex from TopoDS
	---C++: return const &
        ---C++: inline		
    	is static;

	Orientation(myclass; F :Face from TopoDS ) 
        ---C++: inline		
    	    returns Orientation from TopAbs;

    	Orientation(myclass; E : Edge from TopoDS ) 
        ---C++: inline		
    	    returns Orientation from TopAbs;

	Bound(myclass; F :Face from TopoDS ) 
    	    returns Box from Bnd;

    	Bound(myclass; E : Edge from TopoDS ) 
    	    returns Box from Bnd;

	FirstVertex(myclass; E : Edge from TopoDS ) 
    	    returns Vertex from TopoDS
    	raises NoSuchObject; 
    	--if there is not first vertex (semi-infinite edge)

	LastVertex(myclass; E : Edge from TopoDS) 
    	    returns Vertex from TopoDS
    	raises NoSuchObject; 
    	--if there is not last vertex (semi-infinite edge)

	Vertices(myclass; E : Edge from TopoDS;
    	    	 Vfirst, Vlast : out Vertex from TopoDS); 
	---Purpose: If there is  not First or Last vertex (infinite or
	--          semi-infinite edge) return null shapes.

	Range(myclass; E : Edge from TopoDS;
    	    	       F : Face from TopoDS;
    	               wFirst, wLast : in out Real from Standard);
        ---C++: inline		

	UVPoints(myclass; E : Edge from TopoDS;
    	    	          F : Face from TopoDS;
    	                  uvFirst, uvLast : out Pnt2d from gp);
        ---C++: inline		

    	Degenerated(myclass; E : Edge from TopoDS)
        ---C++: inline		
    	    returns Boolean from Standard;

	Tolerance(myclass; V : Vertex from TopoDS)
        ---C++: inline		
    	    returns Real from Standard;

	Parameter(myclass; V : Vertex from TopoDS;
    	    	  E : Edge from TopoDS;
    	    	  F : Face from TopoDS) returns Real from Standard;
        ---C++: inline		

    	Parameters (myclass; 
    	    	    E  : Edge from TopoDS;
    	    	    F  : Face from TopoDS; 
    	    	    W  : Real; 
    	    	    UV : out Pnt2d);
	
    	Locate     (myclass; 
    	    	    C  : Curve from BRepAdaptor;
    	    	    W  : in Real; WFound : in out Real; 
    	    	    p3d : Pnt from gp;
    	    	    UV : out Pnt2d);
	
    	Pnt(myclass; V : Vertex from TopoDS) 
        ---C++: inline
    	    returns Pnt from gp;
	    
	    
	AddInFace(myclass;
	          F : Face                 from TopoDS;
		  T : in out Triangulation from Poly);




fields

    theFIterator : Explorer from TopExp;
    theEIterator : Explorer from TopExp;
    theVIterator : Explorer from TopExp;

end ShapeTool;

