-- Created on: 1992-11-18
-- Created by: Christian CAILLET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



generic class SelectList  from IFSelect (Entity as Transient)
    	inherits SelectInList


    ---Purpose : A SelectList kind Selection selects a part of an Entity, as
    --           well as this Entity can be described as an ordered List.
    --           That is to say, it must have two methods :
    --
    --             NbEntities (me) returns Integer;
    --             Entity (me; num : Integer) returns Transient;
    --           
    --           For each class of Entity for which we want to define a
    --           SelectList, we will instanciate this class with the
    --           desired class of Entity as definition parameter : the deferred
    --           methods NbEntities and ListedEntity are now defined to call
    --           the required methods from <Entity>
    --
    --           SelectList works as SelectInList, beeing a sub-class of it

uses AsciiString from TCollection, Transient, EntityIterator, IntParam

raises OutOfRange

is

    Create returns mutable SelectList;
    ---Purpose : Creates a SelectList (with no limit);

    KeepInputEntity (me; iter : in out EntityIterator);
    ---Purpose : Keeps Input Entity, as having required type <Entity>

    NbItems (me; ent : Transient) returns Integer;
    ---Purpose : Returns count of Entities in the list in the Entity <ent>
    --           by calling method NbEntity from parameter class Entity

    ListedEntity (me; num : Integer; ent : Transient)
    	returns Transient  raises OutOfRange;
    ---Purpose : Returns an Entity of the list in the Entity <ent>, by calling
    --           method Entity from parameter class Entity
    --           Error if <ent> has not required type, or if <num> is not in
    --           the right range (1,NbEntities),

    ListLabel (me) returns AsciiString from TCollection;
    ---Purpose : Returns the specific label for the list
    --           then, following cases :
    --           " From .. Until .." or "From .." or "Until .." or "Rank no .."
    --  Warning : it is not possible to give a character constant to instantiate
    --           a generic class, thus "List From Entity" is not adapted :
    --           redefine Label if judged necessary

end SelectList;
