-- Created on: 2000-03-01
-- Created by: Denis PASCAL
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DrawDocument from DDocStd inherits Data from DDF

	---Purpose: draw variable for TDocStd_Document.
	--          ==================================

uses Document    from TDocStd,
     Drawable3D  from Draw,
     Interpretor from Draw,
     Display     from Draw

is 


    Find (myclass; Doc : Document from TDocStd)
    returns DrawDocument from DDocStd;

    Create (Doc : Document from TDocStd)
    returns DrawDocument from DDocStd;

    GetDocument(me) returns Document from TDocStd;

    DrawOn (me; dis : in out Display from Draw);
    
    Copy (me) 
    returns Drawable3D from Draw
    is redefined;
	
    Dump (me; S : in out OStream) 
    is redefined;
    
    Whatis (me; I : in out Interpretor from Draw)
    is redefined;

fields

    myDocument : Document from TDocStd;

end DrawDocument;
