-- Created on: 1997-04-17
-- Created by: Christophe MARION
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class EdgeIList from HLRBRep

uses
    Orientation          from TopAbs,
    Interference         from HLRAlgo,
    InterferenceList     from HLRAlgo,
    EdgeInterferenceTool from HLRBRep
is
    AddInterference(myclass;
                    IL : in out InterferenceList     from HLRAlgo;
    	            I  :        Interference         from HLRAlgo;
                    T  :        EdgeInterferenceTool from HLRBRep);
	---Purpose: Add the interference <I> to the list <IL>.
    
    ProcessComplex(myclass;
                   IL : in out InterferenceList     from HLRAlgo;
                   T  :        EdgeInterferenceTool from HLRBRep);
	---Purpose: Process complex transitions on the list IL.
    
end EdgeIList;
