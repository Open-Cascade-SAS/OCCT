-- Created on: 1997-03-28
-- Created by: Christian CAILLET
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SizeMember  from StepBasic    inherits SelectReal  from StepData

    ---Purpose : For immediate members of SizeSelect, i.e. :
    --           ParameterValue (a Real)

uses CString

is

    Create returns SizeMember;

    HasName (me) returns Boolean  is redefined;
    -- returns True

    Name (me) returns CString  is redefined;
    -- returns POSITIVE_LENGTH_MEASURE

    SetName (me : mutable; name : CString)  returns Boolean  is redefined;
    -- does nothing (only one case) and returns True

end SizeMember;
