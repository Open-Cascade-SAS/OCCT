-- Created on: 1991-10-03
-- Created by: JeanClaude VAUTHIER 
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

--  Modified : 07/10/97 : JPI/RBV/SMN  : traitement des courbes offset
--  et surfaces offset par approximation 


package GeomConvert

        --- Purpose : The GeomConvert package provides some global functions as follows
    	-- -   converting classical Geom curves into BSpline curves,
    	-- -   segmenting BSpline curves, particularly at knots
    	--   values: this function may be used in conjunction with the
    	--   GeomConvert_BSplineCurveKnotSplitting
    	--   class to segment a BSpline curve into arcs which
    	--   comply with required continuity levels,
    	-- -   converting classical Geom surfaces into BSpline surfaces, and
    	-- -   segmenting BSpline surfaces, particularly at
    	--   knots values: this function may be used in conjunction with the
    	--   GeomConvert_BSplineSurfaceKnotSplitting
    	--   class to segment a BSpline surface into patches
    	--   which comply with required continuity levels.
    	--  All geometric entities used in this package are bounded.
        --  
        -- References :
        --  . Generating the Bezier Points of B-spline curves and surfaces
        --    (Wolfgang Bohm) CAGD volume 13 number 6 november 1981
        --  . On NURBS: A Survey  (Leslie Piegl) IEEE Computer Graphics and
        --    Application January 1991
        --  . Curve and surface construction using rational B-splines 
        --    (Leslie Piegl and Wayne Tiller) CAD Volume 19 number 9 november
        --    1987
        --  . A survey of curve and surface methods in CAGD (Wolfgang BOHM)
        --    CAGD 1 1984


uses    Standard, 
    	TColStd,
    	TColGeom, 
	TColgp,
	GeomAbs,
    	gp, 
    	Geom,
	Geom2d,
    	Convert, 
	AdvApp2Var
	    

is
 
  class BSplineCurveKnotSplitting;
        --- Purpose : This algorithm searches the knot values corresponding to the 
        --  splitting of a given B-spline curve into  several arcs with
        --  the same continuity. The continuity order is given at the
        --  construction time. It is possible to compute the curve arcs
        --  corresponding to this splitting with the method of package 
        --  SplitBSplineCurve.


  class BSplineSurfaceKnotSplitting;
        --- Purpose :
        --  This algorithm searches the knot values corresponding to the
        --  splitting of a given B-spline surface into several patches with
        --  the same continuity. The continuity order is given at the
        --  construction time. It is possible to compute the surface patches
        --  corresponding to the splitting with the method of package
        --  SplitBSplineSurface.


  class BSplineCurveToBezierCurve;
        --- Purpose : 
        --  This algorithm converts a B-spline curve from the package Geom
        --  into several Bezier curves.
        
  class CompCurveToBSplineCurve;
        --- Purpose : 
        --  This algorithm converts and concat sevral curve in a 
        --  B-spline curve.

  class BSplineSurfaceToBezierSurface;
        --- Purpose : 
        --  This algorithm converts a B-spline surface from the package Geom
        --  into several Bezier surfaces.  

 class CompBezierSurfacesToBSplineSurface;
    	---Purpose: Convert a grid of Bezier Surfaces
    	--          that are have continuity CM to an 
    	--          Bspline Surface that has continuity CM
    	   
 class  ApproxSurface;  
        ---Purpose: Convert a surface from Geom by an approximation method
            --          
 class  ApproxCurve;  
        ---Purpose: Convert a curve from Geom by an approximation method
            --
  SplitBSplineCurve (C               : BSplineCurve from Geom; 
                     FromK1, ToK2    : Integer;
                     SameOrientation : Boolean = Standard_True)
     returns mutable BSplineCurve from Geom
         --- Purpose : 
         --  This method computes the arc of B-spline curve between the two 
         --  knots FromK1 and ToK2.  If C is periodic the arc has the same
         --  orientation as C if SameOrientation = Standard_True.  
         --  If C is not periodic  SameOrientation is not used for the
         --  computation and C is oriented from the knot fromK1 to the knot toK2.  
         --  We just keep the local definition of C between the knots
         --  FromK1 and ToK2.  The returned B-spline curve has its first
         --  and last knots with a multiplicity equal to degree + 1, where
         --  degree is the polynomial degree of C.
         --  The indexes of the knots FromK1 and ToK2 doesn't include the
         --  repetition of multiple knots in their definition.
     raises  DomainError from Standard;
         --- Purpose :  Raised if FromK1 = ToK2
         --             Raised if FromK1 or ToK2 are out of the bounds 
         --             [FirstUKnotIndex, LastUKnotIndex]



  SplitBSplineCurve (C                   : BSplineCurve from Geom; 
                     FromU1, ToU2        : Real;
                     ParametricTolerance : Real;
                     SameOrientation     : Boolean = Standard_True)
     returns mutable BSplineCurve from Geom
        --- Purpose :
        --  This function computes the segment of B-spline curve between the 
        --  parametric values FromU1, ToU2.
        --  If C is periodic the arc has the same orientation as C if
        --  SameOrientation = True.  
        --  If C is not periodic SameOrientation is not used for the 
        --  computation and C is oriented fromU1 toU2. 
        --  If U1 and U2 and two parametric values we consider that 
        --  U1 = U2 if Abs (U1 - U2) <= ParametricTolerance and 
        --  ParametricTolerance must  be greater or equal to Resolution
        --  from package gp.
     raises DomainError from Standard;
        --- Purpose :
        --  Raised if FromU1 or ToU2 are out of the parametric bounds of the
        --  curve (The tolerance criterion is ParametricTolerance).
        --  Raised if Abs (FromU1 - ToU2) <= ParametricTolerance
        --  Raised if ParametricTolerance < Resolution from gp.



  SplitBSplineSurface (S : BSplineSurface from Geom; 
                       FromUK1, ToUK2, FromVK1, ToVK2 : Integer; 
                       SameUOrientation : Boolean = Standard_True;
                       SameVOrientation : Boolean = Standard_True)
     returns mutable BSplineSurface from Geom
        --- Purpose : 
        --  Computes the B-spline surface patche between the knots values
        --  FromUK1, ToUK2, FromVK1, ToVK2.
        --  If S is periodic in one direction the patche has the same 
        --  orientation as S in this direction if the flag is true in this
        --  direction (SameUOrientation, SameVOrientation).
        --  If S is not periodic SameUOrientation and SameVOrientation are not
        --  used for the computation and S is oriented FromUK1 ToUK2 and 
        --  FromVK1 ToVK2.
     raises DomainError from Standard;
        --- Purpose :  Raised if 
        --             FromUK1 = ToUK2 or FromVK1 = ToVK2
        --             FromUK1 or ToUK2 are out of the bounds 
        --             [FirstUKnotIndex, LastUKnotIndex]
        --             FromVK1 or ToVK2 are out of the bounds 
        --             [FirstVKnotIndex, LastVKnotIndex]



  SplitBSplineSurface (S : BSplineSurface from Geom; 
                       FromK1, ToK2    : Integer;
                       USplit          : Boolean;
                       SameOrientation : Boolean = Standard_True)
     returns mutable BSplineSurface from Geom
        --- Purpose : 
        --  This method splits a B-spline surface patche between the
        --  knots values FromK1, ToK2 in one direction.
        --  If USplit = True then the splitting direction is the U parametric
        --  direction else it is the V parametric direction.
        --  If S is periodic in the considered direction the patche has the
        --  same orientation as S in this direction if SameOrientation is True
        --  If S is not periodic in this direction SameOrientation is not used
        --  for the computation and S is oriented FromK1 ToK2.
     raises  DomainError from Standard;
        --- Purpose : Raised if FromK1 = ToK2 or if
        --            FromK1 or ToK2 are out of the bounds 
        --            [FirstUKnotIndex, LastUKnotIndex] in the 
        --            considered parametric direction.


  SplitBSplineSurface (S : BSplineSurface from Geom; 
                       FromU1, ToU2, FromV1, ToV2 : Real; 
                       ParametricTolerance        : Real;
                       SameUOrientation           : Boolean = Standard_True;
                       SameVOrientation           : Boolean = Standard_True)
     returns mutable BSplineSurface from Geom
        --- Purpose :
        --  This method computes the B-spline surface patche between the
        --  parametric values FromU1, ToU2, FromV1, ToV2.
        --  If S is periodic in one direction the patche has the same 
        --  orientation as S in this direction if the flag is True in this
        --  direction (SameUOrientation, SameVOrientation).
        --  If S is not periodic SameUOrientation and SameVOrientation are not
        --  used for the computation and S is oriented FromU1 ToU2 and 
        --  FromV1 ToV2.
        --  If U1 and U2 and two parametric values we consider that U1 = U2 if
        --  Abs (U1 - U2) <= ParametricTolerance and ParametricTolerance must
        --  be greater or equal to Resolution from package gp.
     raises DomainError from Standard;
        --- Purpose :
        --  Raised if FromU1 or ToU2 or FromV1 or ToU2 are out of the 
        --  parametric bounds of the surface (the tolerance criterion is
        --  ParametricTolerance).
        --  Raised if Abs (FromU1 - ToU2) <= ParametricTolerance or
        --  Abs (FromV1 - ToV2) <= ParametricTolerance.
        --  Raised if ParametricTolerance < Resolution.



  SplitBSplineSurface (S : BSplineSurface from Geom; 
                       FromParam1, ToParam2 : Real;
                       USplit               : Boolean; 
                       ParametricTolerance  : Real;
                       SameOrientation      : Boolean = Standard_True)
     returns mutable BSplineSurface from Geom
        --- Purpose : 
        --  This method splits the B-spline surface S in one direction
        --  between the parametric values FromParam1, ToParam2.
        --  If USplit = True then the Splitting direction is the U parametric
        --  direction else it is the V parametric direction.
        --  If S is periodic in the considered direction the patche has 
        --  the same orientation as S in this direction if SameOrientation 
        --  is true.
        --  If S is not periodic in the considered direction SameOrientation 
        --  is not used for the computation and S is oriented FromParam1 
        --  ToParam2.
        --  If U1 and U2 and two parametric values we consider that U1 = U2 
        --  if Abs (U1 - U2) <= ParametricTolerance and ParametricTolerance
        --  must be greater or equal to Resolution from package gp.
     raises DomainError from Standard;
        --- Purpose :
        --  Raises if FromParam1 or ToParam2 are out of the parametric bounds
        --  of the surface in the considered direction.
        --  Raises if Abs (FromParam1 - ToParam2) <= ParametricTolerance.


  CurveToBSplineCurve (C                : Curve from Geom ;
    	    	       Parameterisation : ParameterisationType from Convert 
    	    	       =  Convert_TgtThetaOver2)
     returns mutable BSplineCurve from Geom
        --- Purpose : This function converts a non infinite curve from
        --  Geom into a  B-spline curve.  C must be   an ellipse or  a
        --  circle  or a trimmed conic  or a trimmed  line or a Bezier
        --  curve or a trimmed  Bezier curve or a  BSpline curve or  a
        --  trimmed  BSpline curve or  an  OffsetCurve.  The returned  B-spline is
        --  not periodic except  if C is a Circle  or an  Ellipse.  If
        --   the  Parameterisation is  QuasiAngular than  the returned
        --   curve is NOT periodic  in case a  periodic Geom_Circle or
        --  Geom_Ellipse.  For TgtThetaOver2_1 and TgtThetaOver2_2 the
        --   method   raises  an exception  in    case  of a  periodic
        --  Geom_Circle or a Geom_Ellipse ParameterisationType applies
        --   only    if  the curve  is   a  Circle  or  an   ellipse :
        --  TgtThetaOver2,  -- TgtThetaOver2_1, -- TgtThetaOver2_2, --
        --  TgtThetaOver2_3, -- TgtThetaOver2_4,
    	--    
	-- Purpose: this is the classical rational parameterisation
	--                    2
	--               1 - t
	--  cos(theta) = ------
	--                    2
	--               1 + t
	--                   
	--                 2t
	--  sin(theta) = ------
	--                     2
	--                1 + t
	--                   
	--  t = tan (theta/2)        
	-- 
	--  with TgtThetaOver2  the routine will compute the number of spans
	--  using the rule num_spans = [ (ULast - UFirst) / 1.2 ] + 1 
	--  with TgtThetaOver2_N, N  spans will be forced: an error will 
	--  be raized if (ULast - UFirst) >= PI and N = 1,
	--  ULast - UFirst >= 2 PI and N = 2
	--   
	-- QuasiAngular,
	--  here t is a rational function that approximates  
	--  theta ----> tan(theta/2).
	--  Neverthless the composing with above function yields exact
	--  functions whose square sum up to 1
	-- RationalC1 ;
	--  t is replaced by a polynomial function of u so as to grant
	--  C1 contiuity across knots.
	-- Exceptions 
    	--        Standard_DomainError:
    	-- -   if the curve C is infinite, or
    	-- -   if C is a (complete) circle or ellipse, and Parameterisation is equal to
    	--   Convert_TgtThetaOver2_1 or Convert_TgtThetaOver2_2.
    	--   Standard_ConstructionError:
    	-- -   if C is a (complete) circle or ellipse, and if Parameterisation is not equal to
    	--   Convert_TgtThetaOver2, Convert_RationalC1,
    	--   Convert_QuasiAngular (the curve is converted
    	--   in these three cases) or to Convert_TgtThetaOver2_1 or
    	--   Convert_TgtThetaOver2_2 (another exception is raised in these two cases).
    	-- -   if C is a trimmed circle or ellipse, if Parameterisation is equal to
    	--   Convert_TgtThetaOver2_1 and if U2 - U1 > 0.9999 * Pi, where U1 and U2 are
    	--   respectively the first and the last parameters of the
    	--   trimmed curve (this method of parameterization
    	--   cannot be used to convert a half-circle or a half-ellipse, for example), or
    	-- -   if C is a trimmed circle or ellipse, if
    	--   Parameterisation is equal to Convert_TgtThetaOver2_2 and U2 - U1 >
    	--   1.9999 * Pi where U1 and U2 are
    	--   respectively the first and the last parameters of the
    	--   trimmed curve (this method of parameterization
    	--   cannot be used to convert a quasi-complete circle or ellipse). 
     raises DomainError,
      	    ConstructionError;
	
  SurfaceToBSplineSurface (S : Surface from Geom)
     returns mutable BSplineSurface from Geom
        --- Purpose : 
        --  This algorithm converts a non infinite surface from Geom
        --  into a B-spline surface.
        --  S must be a trimmed plane or a trimmed cylinder or a trimmed cone
        --  or a trimmed sphere or a trimmed torus or a sphere or a torus or
        --  a Bezier surface of a trimmed Bezier surface or a trimmed swept
        --  surface with a corresponding basis curve which can be turned into
        --  a B-spline curve   (see the method CurveToBSplineCurve).
    	--  Raises DomainError if the type of the surface is not previously defined.
     raises DomainError;
      
  ConcatG1(ArrayOfCurves  : in out Array1OfBSplineCurve from TColGeom;
    	   ArrayOfToler   : in           Array1OfReal   from TColStd;
    	   ArrayOfConcatenated    : out  HArray1OfBSplineCurve from TColGeom;
	   ClosedG1Flag           : in   Boolean                from Standard ;
	   ClosedTolerance        : in   Real                   from Standard) ;
    	   
    	--- Purpose : This Method concatenates G1 the ArrayOfCurves as far
    	--  as it  is possible.  
    	--  ArrayOfCurves[0..N-1]
    	--  ArrayOfToler contains the  biggest tolerance of the two
    	--               points shared by two consecutives curves.
    	--               Its dimension: [0..N-2]
    	--  ClosedG1     indicates if the ArrayOfCurves is closed.
    	--               In this case ClosedG1 contains the biggest tolerance
    	--               of the two points which are at the closure.
    	--               Otherwise its value is 0.0


  ConcatC1(ArrayOfCurves  : in out Array1OfBSplineCurve from TColGeom;
    	   ArrayOfToler   : in           Array1OfReal   from TColStd;
	   ArrayOfIndices : out        HArray1OfInteger from TColStd;
    	   ArrayOfConcatenated    : out  HArray1OfBSplineCurve from TColGeom;
	   ClosedG1Flag           : in   Boolean                 from Standard ;
	   ClosedTolerance        : in   Real                   from Standard) ;

    	--- Purpose : This Method concatenates C1 the ArrayOfCurves as far
    	--  as it is possible.
    	--  ArrayOfCurves[0..N-1]
    	--  ArrayOfToler contains the  biggest tolerance of the two
    	--               points shared by two consecutives curves.
    	--               Its dimension: [0..N-2]
    	--  ClosedG1     indicates if the ArrayOfCurves is closed.
    	--               In this case ClosedG1 contains the biggest tolerance
    	--               of the two points which are at the closure.
    	--               Otherwise its value is 0.0

   ConcatC1(ArrayOfCurves         : in out Array1OfBSplineCurve from TColGeom;
    	   ArrayOfToler           : in           Array1OfReal   from TColStd;
	   ArrayOfIndices         : out        HArray1OfInteger from TColStd;
    	   ArrayOfConcatenated    : out  HArray1OfBSplineCurve from TColGeom;
    	   ClosedG1Flag           : in   Boolean              from Standard ;
	   ClosedTolerance        : in   Real               from Standard ;
	   AngularTolerance       : in Real                  from Standard) ;
	   
    	--- Purpose : This Method concatenates C1 the ArrayOfCurves as far
    	--  as it is possible.
    	--  ArrayOfCurves[0..N-1]
    	--  ArrayOfToler contains the  biggest tolerance of the two
    	--               points shared by two consecutives curves.
    	--               Its dimension: [0..N-2]
    	--  ClosedG1     indicates if the ArrayOfCurves is closed.
    	--               In this case ClosedG1 contains the biggest tolerance
    	--               of the two points which are at the closure.
    	--               Otherwise its value is 0.0
    	-- 

  C0BSplineToC1BSplineCurve(BS              : in out BSplineCurve from Geom;
    	    	    	    tolerance       : in Real from Standard; 
                            AngularTolerance: in Real =  1.0e-7);
    	---Purpose : This  Method reduces as far as   it is possible the
    	--  multiplicities of  the  knots of  the BSpline BS.(keeping  the
    	--  geometry).  It returns a new BSpline which  could still be C0.
    	--  tolerance is a  geometrical tolerance.   
	--  The  Angular toleranceis in radians  and mesures  the angle of
    	--  the tangents  on  the left and on  the right  to decide if  the
    	-- curve is G1 or not at a given point


  C0BSplineToArrayOfC1BSplineCurve(BS        : in  BSplineCurve from Geom;
    	    	    	    	   tabBS     : out HArray1OfBSplineCurve from TColGeom;
				   tolerance : in Real from Standard);
    	--- Purpose : This Method   reduces as far  as  it is possible  the
    	--  multiplicities  of  the knots  of the BSpline  BS.(keeping the geometry).
    	--  It returns an array of BSpline C1. tolerance is a geometrical tolerance.
 
  C0BSplineToArrayOfC1BSplineCurve(BS               : in  BSplineCurve from Geom;
    	    	    	    	   tabBS            : out HArray1OfBSplineCurve from TColGeom;
				   AngularTolerance : in Real from Standard ;
				   tolerance        : in Real from Standard);
    	--- Purpose :This   Method reduces as far   as it is  possible the
    	--  multiplicities of  the  knots of  the  BSpline BS.(keeping the
    	--  geometry).  It returns an array of BSpline C1.  tolerance is a
    	--  geometrical tolerance : it  allows for the maximum deformation
    	--  The  Angular tolerance is in  radians and mesures the angle of
    	--  the tangents on the left and on the right to decide if the curve
    	--  is C1 or not at a given point

end GeomConvert;










