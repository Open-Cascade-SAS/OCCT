-- File:	IFSelect_AppliedModifiers.cdl
-- Created:	Mon May  2 18:34:11 1994
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1994


class AppliedModifiers  from IFSelect  inherits TShared

    ---Purpose : This class allows to memorize and access to the modifiers
    --           which are to be applied to a file. To each modifier, is bound
    --           a list of integers (optionnal) : if this list is absent, the
    --           modifier applies to all the file. Else, it applies to the
    --           entities designated by these numbers in the produced file.
    --           
    --           To record a modifier, and a possible list of entity numbers
    --           to be applied on :
    --             AddModif (amodifier);
    --             loop on  AddNum (anumber);
    --           
    --           To query it,  Count gives the count of recorded modifiers,
    --           then for each one :
    --             Item (numodif, amodifier, entcount);
    --             IsForAll ()  -> can be called, if True, applies on the whole file
    --             
    --             for (i = 1; i <= entcount; i ++)
    --               nument = ItemNum (i);  -> return an entity number

uses  GeneralModifier, SequenceOfGeneralModifier,
      HSequenceOfInteger from TColStd, IntList

is

    Create (nbmax,nbent : Integer) returns mutable AppliedModifiers;
    ---Purpose : Creates an AppliedModifiers, ready to record up to <nbmax>
    --           modifiers, on a model of <nbent> entities

    AddModif (me : mutable; modif : mutable GeneralModifier) returns Boolean;
    ---Purpose : Records a modifier. By default, it is to apply on all a
    --           produced file. Further calls to AddNum will restrict this.
    --           Returns True if done, False if too many modifiers are already
    --           recorded

    AddNum (me : mutable; nument : Integer) returns Boolean;
    ---Purpose : Adds a number of entity of the output file to be applied on.
    --           If a sequence of AddNum is called after AddModif, this
    --           Modifier will be applied on the list of designated entities.
    --           Else, it will be applied on all the file
    --           Returns True if done, False if no modifier has yet been added

    Count (me) returns Integer;
    ---Purpose : Returns the count of recorded modifiers

    Item (me : mutable; num : Integer;
    	  modif : out mutable GeneralModifier; entcount : out Integer)
	    returns Boolean;
    ---Purpose : Returns the description for applied modifier n0 <num> :
    --           the modifier itself, and the count of entities to be applied
    --           on. If no specific list of number has been defined, returns
    --           the total count of entities of the file
    --           If this count is zero, then the modifier applies to all
    --           the file (see below). Else, the numbers are then queried by
    --           calls to ItemNum between 1 and <entcount>
    --           Returns True if OK, False if <num> is out of range

    ItemNum (me; nument : Integer) returns Integer;
    ---Purpose : Returns a numero of entity to be applied on, given its rank
    --           in the list. If no list is defined (i.e. for all the file),
    --           returns <nument> itself, to give all the entities of the file
    --           Returns 0 if <nument> out of range

    ItemList (me) returns HSequenceOfInteger;
    ---Purpose : Returns the list of entities to be applied on (see Item)
    --           as a HSequence (IsForAll produces the complete list of all
    --           the entity numbers of the file

    IsForAll (me) returns Boolean;
    ---Purpose : Returns True if the applied modifier queried by last call to
    --           Item is to be applied to all the produced file.
    --           Else, <entcount> returned by Item gives the count of entity
    --           numbers, each one is queried by ItemNum

fields

    themodifs : SequenceOfGeneralModifier;
    thelists  : IntList;
    thenbent  : Integer;
    theentcnt : Integer;

end AppliedModifiers;
