-- Created on: 1991-06-18
-- Created by: Didier PIFFAULT
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class TangentZone from Intf

	---Purpose: Describes   a  zone  of  tangence  between  polygons  or
	--          polyhedra as a sequence of points of intersection.

uses    SectionPoint from Intf,
    	SeqOfSectionPoint from Intf


raises  OutOfRange from Standard


is

-- User Interface :

    NumberOfPoints (me)
    	    	    returns Integer is static;
    ---Purpose: Returns number of SectionPoint in this TangentZone.
    ---C++: inline

    GetPoint       (me;
    	    	    Index    : in Integer)
    	    	    returns SectionPoint from Intf
    	    	    raises OutOfRange from Standard
    	    	    is static;
    ---Purpose: Gives   the   SectionPoint   of  address  <Index>  in  the
    --          TangentZone.
    --          
    ---C++: return const &


    IsEqual        (me;
    	    	    Other    : in TangentZone from Intf)
    	    	    returns Boolean is static;
    ---Purpose: Compares two TangentZones.
    --          
    ---C++: alias operator ==


    Contains       (me;
    	    	    ThePI    : in SectionPoint from Intf)
    	    	    returns Boolean is static;
    ---Purpose: Checks if <ThePI> is in TangentZone.


    ParamOnFirst   (me;
    	    	    paraMin : in out Real from Standard;
    	    	    paraMax : in out Real from Standard) is static;
    ---C++: inline
    ---Purpose: Gives  the parameter range of the  TangentZone on the first
    --          argument of the Interference. (Usable only for polygon)


    ParamOnSecond  (me;
    	    	    paraMin : in out Real from Standard;
    	    	    paraMax : in out Real from Standard) is static;
    ---C++: inline
    ---Purpose: Gives the parameter range of the  TangentZone on the second
    --          argument of the Interference. (Usable only for polygon)


    InfoFirst      (me;
    	    	    segMin  : in out Integer from Standard;
    	    	    paraMin : in out Real from Standard;
    	    	    segMax  : in out Integer from Standard;
    	    	    paraMax : in out Real from Standard) is static;
    ---Purpose: Gives information  about  the    first argument   of   the
    --          Interference. (Usable only for polygon)

    InfoSecond     (me;
    	    	    segMin  : in out Integer from Standard;
    	    	    paraMin : in out Real from Standard;
    	    	    segMax  : in out Integer from Standard;
    	    	    paraMax : in out Real from Standard) is static;
    ---Purpose: Gives   informations  about  the  second   argument of  the
    --          Interference. (Usable only for polygon)


    RangeContains  (me;
    	    	    ThePI    : in SectionPoint from Intf)
    	    	    returns Boolean is static;
    ---Purpose: Returns True if  <ThePI>  is in the parameter  range of the
    --          TangentZone.

    HasCommonRange (me;
    	    	    Other    : in TangentZone from Intf)
    	    	    returns Boolean is static;
    ---Purpose: Returns True if the TangentZone  <Other> has  a common part
    --          with <me>.


-- Builder :

    Create          returns TangentZone;
    ---Purpose: Builds an empty tangent zone.

    Create         (Other : TangentZone)
            	    returns TangentZone;
    ---Purpose: Copies a Tangent zone.


    Append         (me       : in out;
    	    	    Pi       : SectionPoint from Intf)
    	    	    is static;
    ---Purpose: Adds a SectionPoint to the TangentZone.


    Append         (me       : in out;
    	    	    Tzi      : TangentZone from Intf)
    	    	    is static;
    ---Purpose: Adds the TangentZone <Tzi> to <me>.


    Insert         (me       : in out;
    	    	    Pi       : SectionPoint from Intf)
		    returns Boolean
    	    	    is static;
    ---Purpose: Inserts a SectionPoint in the TangentZone.


    PolygonInsert  (me       : in out;
    	    	    Pi       : SectionPoint from Intf)
    	    	    is static;
    ---Purpose: Inserts a point in the polygonal TangentZone.


    InsertBefore   (me       : in out;
    	    	    Index    : in Integer;
    	    	    Pi       : SectionPoint from Intf)
    	    	    is static;
    ---Purpose: Inserts a SectionPoint before <Index> in the TangentZone.

    InsertAfter    (me       : in out;
    	    	    Index    : in Integer;
    	    	    Pi       : SectionPoint from Intf)
    	    	    is static;
    ---Purpose: Inserts a SectionPoint after <Index> in the TangentZone.


    Dump           (me;
    	    	    Indent   : in Integer) is static;

fields

    Result            : SeqOfSectionPoint;
    ParamOnFirstMin   : Real from Standard;
    ParamOnFirstMax   : Real from Standard;
    ParamOnSecondMin  : Real from Standard;
    ParamOnSecondMax  : Real from Standard;


end TangentZone;
