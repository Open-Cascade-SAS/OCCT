-- File:	RWStepElement_RWCurve3dElementDescriptor.cdl
-- Created:	Thu Dec 12 17:28:59 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWCurve3dElementDescriptor from RWStepElement

    ---Purpose: Read & Write tool for Curve3dElementDescriptor

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    Curve3dElementDescriptor from StepElement

is
    Create returns RWCurve3dElementDescriptor from RWStepElement;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : Curve3dElementDescriptor from StepElement);
	---Purpose: Reads Curve3dElementDescriptor

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: Curve3dElementDescriptor from StepElement);
	---Purpose: Writes Curve3dElementDescriptor

    Share (me; ent : Curve3dElementDescriptor from StepElement;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWCurve3dElementDescriptor;
