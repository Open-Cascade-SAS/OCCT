-- Created on: 2007-12-04
-- Created by: Sergey ZARITCHNY
-- Copyright (c) 2007-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DeltaOnModificationOfExtStringArray from TDataStd inherits DeltaOnModification from TDF

	---Purpose: This class provides default services for an
	--          AttributeDelta on a MODIFICATION action.

uses
    Attribute               from TDF,
    HArray1OfExtendedString from TColStd,
    ExtStringArray          from TDataStd, 
    HArray1OfInteger        from TColStd 
    
is
    Create (Arr : ExtStringArray     from TDataStd)
    	returns mutable DeltaOnModificationOfExtStringArray from TDataStd;
	---Purpose: Initializes a TDF_DeltaOnModification.

    Apply (me : mutable)
    	is redefined virtual;
    	---Purpose: Applies the delta to the attribute.
fields
 myIndxes  :  HArray1OfInteger from TColStd; 
 myValues  :  HArray1OfExtendedString from TColStd; 
 myUp1     :  Integer          from Standard;
 myUp2     :  Integer          from Standard; 
 
end DeltaOnModificationOfExtStringArray;


