-- Created on: 1992-05-27
-- Created by: Remi LEQUETTE
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.





class TFace from PBRep inherits TFace from PTopoDS

	---Purpose: The Tface from PBRep  is  based  on the TFace  from
	--          TopoDS. The TFace contains :
	--          
	--          * A surface, a tolerance, a location
	--          
	--          * A NaturalRestriction flag,   when this  flag  is
	--          True the  boundary of the  face is known to be the
	--          parametric space (Umin, UMax, VMin, VMax).

uses
    Surface       from PGeom,
    Triangulation from PPoly,
    Location      from PTopLoc
    
is

    Create returns mutable TFace from PBRep;
	---Purpose: Creates an empty TFace.
    	---Level: Internal 
	
    
    Surface(me) returns Surface from PGeom
    is static;
    	---Level: Internal 

    Triangulation(me) returns any Triangulation from PPoly
    is static;
	---Level: Internal    

    Location(me) returns Location from PTopLoc
    is static;
    	---Level: Internal 
    	
    Tolerance(me) returns Real
    is static;
    	---Level: Internal 

    Surface(me : mutable; S : Surface from PGeom)
    is static;
    	---Level: Internal 

    Triangulation(me : mutable; T : Triangulation from PPoly)
    is static;
	---Level: Internal 
    	
    Location(me : mutable; L : Location from PTopLoc)
    is static;
    	---Level: Internal 
    	
    Tolerance(me : mutable; T : Real)
    is static;
    	---Level: Internal 

    NaturalRestriction(me) returns Boolean
    is static;
    	---Level: Internal 
    
    NaturalRestriction(me : mutable; N : Boolean)
    is static;
    	---Level: Internal 
    
fields

    mySurface            : Surface  from PGeom;
    myTriangulation      : Triangulation from PPoly;
    myLocation           : Location from PTopLoc;
    myTolerance          : Real;
    myNaturalRestriction : Boolean;

end TFace;

