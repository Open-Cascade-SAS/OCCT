-- Created on: 1993-02-25
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class BlockIterator from TopOpeBRepBuild 

---Purpose: Iterator on the elements of a block.

raises

    NoMoreObject from Standard

is

    Create returns BlockIterator from TopOpeBRepBuild;
    Create(Lower,Upper : Integer from Standard) 
    returns BlockIterator from TopOpeBRepBuild;
    
    Initialize(me : in out) is static;
    ---C++: inline
    More(me) returns Boolean from Standard is static;
    ---C++: inline
    Next(me : in out) raises NoMoreObject is static;
    ---C++: inline
    Value(me) returns Integer from Standard is static;
    ---C++: inline
    Extent(me) returns Integer from Standard is static;
    ---C++: inline

fields

    myLower : Integer from Standard;
    myUpper : Integer from Standard;
    myValue : Integer from Standard;

end BlockIterator from TopOpeBRepBuild;
