-- File:	StepToGeom_MakeLine2d.cdl
-- Created:	Wed Aug  4 10:53:16 1993
-- Author:	Martine LANGLOIS
---Copyright:	 Matra Datavision 1993

class MakeLine2d from StepToGeom

    ---Purpose: This class implements the mapping between classes 
    --          Line from StepGeom which describes a line from
    --          Prostep and Line from Geom2d.
  
uses 
     Line from Geom2d,
     Line from StepGeom
     
is 

    Convert ( myclass; SC : Line from StepGeom;
                       CC : out Line from Geom2d )
    returns Boolean from Standard;

end MakeLine2d;
