-- Created on: 1996-06-05
-- Created by: Mister rmi
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PolygonOnTriangulation from PPoly inherits Persistent from Standard

    	---Purpose: This class represents a 3d Polygon based on
    	--          indices of triangulation nodes.
    	--          
    	--          This polygon may also have a parametric
    	--          representation.


uses HArray1OfInteger  from PColStd,
     HArray1OfReal     from PColStd

raises NullObject from Standard

is

    Create returns mutable PolygonOnTriangulation from PPoly;
    
    Create(Nodes : HArray1OfInteger from PColStd;
    	   Defl  : Real             from Standard)
    returns mutable PolygonOnTriangulation from PPoly;
    	---Purpose: Defaults with allocation of nodes.
    
    Create(Nodes      : HArray1OfInteger from PColStd;
       	   Defl       : Real             from Standard;
           Parameters : HArray1OfReal    from PColStd) 
    returns mutable PolygonOnTriangulation from PPoly;
    	---Purpose: Defaults with allocation of nodes.
    
    Deflection(me) returns Real;
    
    Deflection(me : mutable; D : Real);


    NbNodes(me) returns Integer;
    
    Nodes(me) returns HArray1OfInteger from PColStd;
	---Purpose: Reference on the 3d nodes indices.

    Nodes(me : mutable; Nodes : HArray1OfInteger from PColStd);
    
    HasParameters(me) returns Boolean from Standard;
    
    Parameters(me) returns HArray1OfReal from PColStd;
	---Purpose: Returns the parameters values.

    Parameters(me : mutable; Param : HArray1OfReal from PColStd);
    
    
fields

    myDeflection    : Real             from Standard;
    myNodes         : HArray1OfInteger from PColStd;
    myParameters    : HArray1OfReal    from PColStd; 
    	 -- myParameters is Optional (pointer can be null)
    
end PolygonOnTriangulation;
