-- Created on: 1999-10-25
-- Created by: Sergey ZARITCHNY <szy@philipox.nnov.matra-dtv.fr>
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Loader from QANewBRepNaming 

    	---Purpose: 

uses MakeShape      from BRepBuilderAPI, 
     Shape          from TopoDS,  
     Edge           from TopoDS,
     ShapeEnum      from TopAbs, 
     Builder        from TNaming, 
     DataMapOfShapeShape from TopTools, 
     MapOfShape     from TopTools,
     Label          from TDF, 
     TagSource      from TDF

is 

    LoadGeneratedShapes (myclass; 
			 MakeShape          : in out MakeShape from BRepBuilderAPI;
    	    	    	 ShapeIn       : in     Shape     from TopoDS;
			 GeneratedFrom : in     ShapeEnum from TopAbs;
			 Buider        : in out Builder   from TNaming);
    	---Purpose :  Load in   the naming data-structure   the  shape
    	--          generated  from FACE,  EDGE, VERTEX,..., after the
    	--          MakeShape   operation.  <ShapeIn>  is  the initial
    	--          shape.   <GeneratedFrom>   defines  the   kind  of
    	--          shape generation    to    record  in   the  naming
    	--          data-structure. The <builder> is used to store the
    	--          set of evolutions in the data-framework of TDF.

			 
    LoadModifiedShapes (myclass; 
		        MakeShape          : in out MakeShape from BRepBuilderAPI; 
    	    	    	ShapeIn      : in     Shape     from TopoDS;
			ModifiedFrom : in     ShapeEnum from TopAbs;
			Buider       : in out Builder   from TNaming; 
    	    	    	theBool      : Boolean from Standard = Standard_False);
    	---Purpose  : Load in the naming data-structure the shape
    	--              modified from FACE, EDGE, VERTEX,...,
    	--              after the MakeShape operation.
    	--            <ShapeIn> is the initial shape.
    	--            <ModifiedFrom> defines the kind of shape modification
    	--              to record in the naming data-structure.
    	--            The <builder> is used to store the set of evolutions
    	--              in the data-framework of TDF.
	 
   LoadDeletedShapes (myclass; 
		      MakeShape          : in out MakeShape from BRepBuilderAPI; 
    	    	      ShapeIn            : in     Shape     from TopoDS;
		      KindOfDeletedShape : in     ShapeEnum from TopAbs;
		      Buider             : in out Builder   from TNaming);
    	---Purpose : Load in the naming data-structure the shape
    	--             deleted after the MakeShape operation.
    	--           <ShapeIn> is the initial shape.
    	--           <KindOfDeletedShape> defines the kind of
    	--             deletion to record in the naming data-structure.
    	--           The <builder> is used to store the set of evolutions
    	--             in the data-framework of TDF.		       
		      
    LoadAndOrientGeneratedShapes (myclass;
      MakeShape          : in out MakeShape from BRepBuilderAPI;
      ShapeIn            : in     Shape               from TopoDS;
      GeneratedFrom      : in     ShapeEnum           from TopAbs;
      Buider             : in out Builder             from TNaming;
      SubShapesOfResult  : in     DataMapOfShapeShape from TopTools);        
      ---Purpose  : The same as LoadGeneratedShapes plus performs orientation of
      --           loaded shapes according orientation of SubShapes


    LoadAndOrientModifiedShapes (myclass;
      MakeShape          : in out MakeShape from BRepBuilderAPI;
      ShapeIn            : in     Shape               from TopoDS;
      ModifiedFrom       : in     ShapeEnum           from TopAbs;
      Buider             : in out Builder             from TNaming;
      SubShapesOfResult  : in     DataMapOfShapeShape from TopTools);        
      ---Purpose  : The same as LoadModifiedShapes plus performs orientation of
      --            loaded shapes according orientation of SubShapes


    ModifyPart (myclass; 
    	    	PartShape  : in     Shape    from TopoDS;
    	    	Primitive  : in     Shape    from TopoDS;
       	    	Label      : in     Label    from TDF);
    	---Category: Tool
	---Level: Internal
    
    HasDangleShapes(myclass; ShapeIn : in Shape from TopoDS) 
    returns Boolean from Standard;

    LoadGeneratedDangleShapes(myclass;  
    	    	 	      ShapeIn       : in     Shape from TopoDS; 
		     	      GeneratedFrom : in     ShapeEnum from TopAbs; 
		     	      GenBuider     : in out Builder from TNaming);  

    LoadGeneratedDangleShapes(myclass;  
    	    	 	      ShapeIn       : in     Shape from TopoDS; 
		     	      GeneratedFrom : in     ShapeEnum from TopAbs;  
			      OnlyThese     : in     MapOfShape from TopTools;
		     	      GenBuider     : in out Builder from TNaming); 

    LoadModifiedDangleShapes(myclass;   
    	    	    	     MakeShape     : in out MakeShape from BRepBuilderAPI;
    	    	 	     ShapeIn       : in     Shape from TopoDS; 
		     	     GeneratedFrom : in     ShapeEnum from TopAbs; 
		     	     GenBuider     : in out Builder from TNaming); 

    LoadDeletedDangleShapes(myclass;  
    	    	    	    MakeShape     : in out MakeShape from BRepBuilderAPI;
    	    	 	    ShapeIn       : in     Shape from TopoDS; 
		     	    ShapeType     : in     ShapeEnum from TopAbs; 
		     	    DelBuider     : in out Builder from TNaming); 
    
    LoadDangleShapes(myclass;  
		     theShape : Shape from TopoDS;		     
		     theLabelGenerator : Label from TDF); 

    LoadDangleShapes(myclass;  
		     theShape : Shape from TopoDS;	
		     ignoredShape : Shape from TopoDS;	     
		     theLabelGenerator : Label from TDF); 

    GetDangleShapes(myclass;
    	    	    ShapeIn : Shape from TopoDS;
		    GeneratedFrom : ShapeEnum from TopAbs;
    	    	    Dangles : out DataMapOfShapeShape from TopTools)
    ---Purpose: Returns dangle sub shapes Generator - Dangle.
    returns Boolean from Standard;

    GetDangleShapes(myclass;
    	    	    ShapeIn : Shape from TopoDS;
		    GeneratedFrom : ShapeEnum from TopAbs;
    	    	    Dangles : out MapOfShape from TopTools)
    ---Purpose: Returns dangle sub shapes.
    returns Boolean from Standard;

    IsDangle(myclass;
    	     theDangle : Shape from TopoDS;
	     theShape : Shape from TopoDS)
    ---Warning!: Don't use this method inside an iteration process!
    returns Boolean from Standard;

end Loader;
