-- Created on: 1995-11-28
-- Created by: Jean-Pierre COMBE
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PerpenPresentation from DsgPrs

        ---Purpose: A framework to define display of perpendicular
    	-- constraints between shapes.
uses
    Presentation from Prs3d,
    Pnt from gp,
    Dir from gp,
    Drawer from Prs3d,
    ExtendedString from TCollection
    	
is  
    Add( myclass; aPresentation: Presentation from Prs3d;
    	    	  aDrawer: Drawer from Prs3d;
    	    	  pAx1:          Pnt from gp;
		  pAx2:          Pnt from gp;
                  pnt1:          Pnt from gp;
		  pnt2:          Pnt from gp;
		  OffsetPoint:   Pnt from gp;
    	    	  intOut1:       Boolean from Standard;
    	    	  intOut2:       Boolean from Standard);
	---Purpose: Defines the display of elements showing
    	-- perpendicular constraints between shapes.
    	-- These include the two axis points pAx1 and pAx2,
    	-- the two points pnt1 and pnt2, the offset point
    	-- OffsetPoint and the two Booleans intOut1} and intOut2{.
    	-- These arguments are added to the presentation
    	-- object aPresentation. Their display attributes are
    	-- defined by the attribute manager aDrawer.


end PerpenPresentation;
