-- Created on: 1993-01-22
-- Created by: Gilles DEBARBOUILLE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class DynamicClass from Dynamic

inherits

    TShared from MMgt 
	---Purpose: A  dynamic class  is  defined   as a  sequence  of
	--          parameters and   as a   sequence of   methods. The
	--          specifications  are similar   to C++  classes. The
	--          class  has  to  be   defined  in terms  of  fields
	--          (Parameters) and methods. An instance of the class
	--          must be   made to set  the  fields and to  use the
	--          functionalities.

    
uses

    OStream from Standard,
    CString from Standard,
    HAsciiString      from TCollection,
    DynamicInstance   from Dynamic,
    Parameter         from Dynamic,
    ParameterNode     from Dynamic,
    Method            from Dynamic,
    SequenceOfMethods from Dynamic

    
is

    Create(aname : CString from Standard) returns mutable DynamicClass from Dynamic;
    
    ---Level: Public 
    
    ---Purpose: Creates a new empty instance of DynamicClass.
    
    Parameter(me : mutable ; aparameter : Parameter from Dynamic)
    
    ---Level: Public 
    
    ---Purpose: Adds another parameter <aparameter> to the sequence of
    --          parameter definitions.
    
    is static;
    
    CompiledMethod(me : mutable ; amethod , anaddress : CString from Standard)
    
    ---Level: Public 
    
    ---Purpose: Adds another method to the sequence of methods. It has
    --          <amethod> as name  and <anaddress> as mangled  name of
    --          the corresponding C++ function which must be called.
    
    is static;
    
    InterpretedMethod(me : mutable ; amethod , afile : CString from Standard)
    
    ---Level: Public 
    
    ---Purpose: Adds  another method to the  sequence of methods.   It
    --          has <amethod> as name and <afile> as interpreted file.
    
    is static;
    
    Method(me ; amethod : CString from Standard) returns any Method from Dynamic
    
    ---Level: Public 
    
    ---Purpose: Returns a reference to the method object identified by
    --          the string <amethod>.
    
    is virtual;
    
    Instance(me) returns mutable DynamicInstance from Dynamic
    
    ---Level: Public 
    
    ---Purpose: Returns an instance object of this class.

    is virtual;

    Dump(me ; astream : in out OStream from Standard)
    
    ---Level: Internal 
    
    ---Purpose: useful for debugging.

    is virtual;
    
fields

    thename               : HAsciiString      from TCollection;
    thefirstparameternode : ParameterNode     from Dynamic;
    thesequenceofmethods  : SequenceOfMethods from Dynamic;

end ;
