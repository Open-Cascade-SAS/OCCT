-- Created on: 1998-04-17
-- Created by: Andre LIEUTIER
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class  HPG1Constraint  from  NLPlate  inherits  HGPPConstraint from  NLPlate 
---Purpose: define a PinPoint (no G0)  G1 Constraint used to load a Non
--  Linear Plate
uses
     XY from gp,
     D1  from  Plate
     
is
    Create(UV : XY; D1T : D1 from Plate) returns mutable HPG1Constraint;
    -- create a G1 Constraint
    -- 


    SetIncrementalLoadAllowed(me: mutable; ILA : Boolean) 
    is  redefined;
    -- If True, allow the Constraint to be loaded incrementally during optimization
    -- default is False
    -- 

    SetOrientation(me:  mutable; Orient  :  Integer  =  0) 
    is  redefined;
    --  set the orientation (meaningless for non G1 Constraints) 
    -- 	-1 means that the Surface Normal have to be -1*the Constraint Normal
    --  0  means that G1 constraint is up to a normal inversion (default value)
    --  1  means that the Surface Normal have to be equal to the Constraint Normal.
    --  remarks : within the current implementation, this is effective only in case of
    --  incremental loading computation


    IncrementalLoadAllowed(me)  returns  Boolean 
    is redefined;
    -- If True, allow the Constraint to be loaded incrementally during optimization
    -- default is False
    -- 

    ActiveOrder(me)  returns  Integer 
    is   redefined; 
    --  returns the constraint active  order, i.e. the maximum between
    --  -- the initial constraint i.e 1 (for G1 Constraints)
    --  
    -- 

    IsG0(me) returns Boolean 
    is  redefined;

    Orientation(me:  mutable)  returns  Integer
    is  redefined;
    --  set the orientation (meaningless for  non G1 Constraints)
    -- 	-1 means that the Surface Normal have to be -1*the Constraint Normal
    --  0  means that G1 constraint is up to a normal inversion (default value)
    --  1  means that the Surface Normal have to be equal to the Constraint Normal.
    --  remarks : within the current implementation, this is effective only in case of
    --  incremental loading computation
    -- 

    G1Target(me) returns D1  from  Plate 
    ---C++: return const &
    is   redefined; 

fields
    IncrementalLoadingAllowed : Boolean;
    myG1Target : D1 from Plate; 
    myOrientation  :  Integer;
end;
