-- Created on: 1993-01-11
-- Created by: SIVA
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package IGESSolid


        ---Purpose : This package consists of B-Rep and CSG Solid entities

uses

        Standard,
        TCollection,
	TColStd,
	TColgp,
        gp,
	Message,
        Interface,
        IGESData,
        IGESBasic,
        IGESGeom

is

        class Block;

        class RightAngularWedge;

        class Cylinder;

        class ConeFrustum;

        class Sphere;

        class Torus;

        class SolidOfRevolution;

        class SolidOfLinearExtrusion;

        class Ellipsoid;

        class BooleanTree;

        class SelectedComponent;

        class SolidAssembly;

        class ManifoldSolid;

        class PlaneSurface;

        class CylindricalSurface;

        class ConicalSurface;

        class SphericalSurface;

        class ToroidalSurface;

        class SolidInstance;

        class VertexList;

        class EdgeList;

        class Loop;

        class Face;

        class Shell;

    	--    Tool for Entities    --

        class ToolBlock;
        class ToolRightAngularWedge;
        class ToolCylinder;
        class ToolConeFrustum;
        class ToolSphere;
        class ToolTorus;
        class ToolSolidOfRevolution;
        class ToolSolidOfLinearExtrusion;
        class ToolEllipsoid;
        class ToolBooleanTree;
        class ToolSelectedComponent;
        class ToolSolidAssembly;
        class ToolManifoldSolid;
        class ToolPlaneSurface;
        class ToolCylindricalSurface;
        class ToolConicalSurface;
        class ToolSphericalSurface;
        class ToolToroidalSurface;
        class ToolSolidInstance;
        class ToolVertexList;
        class ToolEdgeList;
        class ToolLoop;
        class ToolFace;
        class ToolShell;

    -- Definition and Exploitation of Entities defined in this Package

    class Protocol;
    class ReadWriteModule;
    class GeneralModule;
    class SpecificModule;

    class TopoBuilder;

    -- Instantiations

    class  Array1OfLoop       instantiates  Array1 from TCollection (Loop);
    class  Array1OfFace       instantiates  Array1 from TCollection (Face);
    class  Array1OfShell      instantiates  Array1 from TCollection (Shell);
    class  Array1OfVertexList instantiates  Array1 from TCollection (VertexList);
    class HArray1OfLoop       instantiates HArray1 from TCollection (Loop,Array1OfLoop);
    class HArray1OfFace       instantiates HArray1 from TCollection (Face,Array1OfFace);
    class HArray1OfShell      instantiates HArray1 from TCollection (Shell,Array1OfShell);
    class HArray1OfVertexList instantiates HArray1 from TCollection (VertexList,Array1OfVertexList);

    --  Package methods

    Init;
    ---Purpose : Prepares dynamic data (Protocol, Modules) for this package

    Protocol  returns Protocol from IGESSolid;
    ---Purpose : Returns the Protocol for this Package

end IGESSolid;
