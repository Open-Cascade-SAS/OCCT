-- File:        CameraUsage.cdl
-- Created:     Mon Dec  4 12:02:24 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWCameraUsage from RWStepVisual

	---Purpose : Read & Write Module for CameraUsage

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     CameraUsage from StepVisual,
     EntityIterator from Interface

is

	Create returns RWCameraUsage;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable CameraUsage from StepVisual);

	WriteStep (me; SW : in out StepWriter; ent : CameraUsage from StepVisual);

	Share(me; ent : CameraUsage from StepVisual; iter : in out EntityIterator);

end RWCameraUsage;
