-- Created on: 1993-01-09
-- Created by: CKY / Contract Toubro-Larsen ( Deepak PRABHU )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package IGESDefs

        ---Purpose : To embody general definitions of Entities
        --           (Parameters, Tables ...)

uses

        Standard,
        TCollection,
	TColStd,
	Message,
        Interface,
        IGESData,
        IGESBasic,
        IGESGraph

is

        class   AssociativityDef;

        class   MacroDef;

        class   UnitsData;

        class   AttributeDef;

        class   TabularData;

        class   GenericData;

        class   AttributeTable;

    	--    Tools for Entities    --

        class ToolAssociativityDef;
        class ToolMacroDef;
        class ToolUnitsData;
        class ToolAttributeDef;
        class ToolTabularData;
        class ToolGenericData;
        class ToolAttributeTable;

	-- Definition and Exploitation of Entities defined in this Package

        class Protocol;
	class ReadWriteModule;
	class GeneralModule;
	class SpecificModule;

        -- Instantiations

     class  Array1OfTabularData instantiates  Array1 from TCollection(TabularData);

     class HArray1OfTabularData instantiates HArray1 from TCollection
    	(TabularData,Array1OfTabularData);
     class HArray1OfHArray1OfTextDisplayTemplate instantiates
    --	HArray1 (HArray1OfTextDisplayTemplate,Array1OfHArray1OfTextDisplayTemplate);
      JaggedArray from Interface (HArray1OfTextDisplayTemplate from IGESGraph);

        -- Package Methods

    Init;
    ---Purpose : Prepares dynamic data (Protocol, Modules) for this package

    Protocol  returns Protocol from IGESDefs;
    ---Purpose : Returns the Protocol for this Package

end IGESDefs;
