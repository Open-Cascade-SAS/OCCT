-- File:	Materials_MaterialsDictionary.cdl
-- Created:	Mon Jan 18 10:55:43 1993
-- Author:	Gilles DEBARBOUILLE
--		<gde@bravox>
---Copyright:	 Matra Datavision 1993


class MaterialsDictionary from Materials 

	---Purpose: This class creates  a dictionary of materials.

inherits

    Transient
    
uses
    OStream           from  Standard,
    HAsciiString      from TCollection,
    MaterialsSequence from Materials,
    Material          from Materials

raises

    NoSuchObject from Standard

is

    Create returns mutable MaterialsDictionary from Materials;
    ---Level: Internal    
    ---Purpose: Returns a  MaterialsDictionary  object which  contains
    --          the sequence of all the   materials the user wants  to
    --          consider.
    
    Material(me ; amaterial : CString from Standard) returns Material from Materials    
    raises NoSuchObject from Standard   
    ---Level: Internal   
    ---Purpose: Retrieves from the dictionary the object material with
    --          <amaterial> as name.  If <amaterial> does not exist in
    --          the dictionary an exeption is raised.
    is static;
    
    ExistMaterial(me ; aName : CString from Standard) returns Boolean from Standard;
    ---Purpose: True if the materialofname aName exists ...
    
    NumberOfMaterials(me) returns Integer from Standard  
    ---Level: Internal 
    ---Purpose: Returns  the number of  materials previously stored in
    --          the dictionary.
    is static;
    
    Material(me ; anindex : Integer from Standard) returns Material from Materials
    ---Level: Internal
    ---Purpose: This method used  with  the  previous one, allow   the
    --          exploration  of   all  the  dictionary.  It  returns a
    --          Material instance.
    is static;
    
    UpToDate(me) returns Boolean from Standard
    ---Level: Internal
    ---Purpose: Returns true if there has been no  modification of the
    --          file Materials.dat  since the   creation of the dictionary
    --          object, false otherwise.  
    is static;
    
    Dump(me ; astream : in out OStream from Standard )
    ---Level: Internal
    ---Purpose: Useful for debugging.
    is static;
    
fields

    thefilename          : HAsciiString from TCollection;
    thetime              : Integer from Standard;
    thematerialssequence : MaterialsSequence from Materials;

end MaterialsDictionary;
