-- Created on: 1992-11-19
-- Created by: Remi LEQUETTE
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Intersector from BRepClass 
inherits IntConicCurveOfGInter from Geom2dInt

	---Purpose: Intersect an Edge  with a segment.
	--          Implement the Intersector2d required by the classifier.

uses
    Lin2d from gp,
    Dir2d from gp,
    Edge  from BRepClass

is
    Create returns Intersector from BRepClass;
    
    Perform(me : in out; 
    	    L : Lin2d from gp; P : Real; Tol : Real; 
    	    E : Edge from BRepClass)
	---Purpose: Intersect the line segment and the edge.
    is static;

    LocalGeometry(me; E : Edge from BRepClass;
    	    	      U : Real; 
    	    	      T : out Dir2d from gp; 
    	    	      N : out Dir2d from gp; 
    	    	      C : out Real)
	---Purpose: Returns in <T>,  <N> and <C>  the tangent,  normal
	--          and  curvature of the edge  <E> at parameter value
	--          <U>.
    is static;

end Intersector;
