-- Created on: 1993-06-14
-- Created by: Martine LANGLOIS
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MakeDirection from GeomToStep inherits Root from GeomToStep

    ---Purpose: This class implements the mapping between classes 
    --          Direction from Geom, Geom2d and Dir, Dir2d from gp, and the
    --          class Direction from StepGeom which describes a direction
    --          from Prostep. 
  
uses Dir from gp,
     Dir2d from gp,
     Direction from Geom,
     Direction from Geom2d,
     Direction from StepGeom
     
raises NotDone from StdFail
     
is 

Create ( D : Dir from gp ) returns MakeDirection;

Create ( D : Dir2d from gp ) returns MakeDirection;

Create ( D : Direction from Geom ) returns MakeDirection;

Create ( D : Direction from Geom2d ) returns MakeDirection;

Value (me) returns Direction from StepGeom
    raises NotDone
    is static;
    ---C++: return const&
    
fields

    theDirection : Direction from StepGeom;
    	-- The solution from StepGeom
    	
end MakeDirection;


