-- File:	IGESAppli_ToolFlowLineSpec.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolFlowLineSpec  from IGESAppli

    ---Purpose : Tool to work on a FlowLineSpec. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses FlowLineSpec from IGESAppli,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolFlowLineSpec;
    ---Purpose : Returns a ToolFlowLineSpec, ready to work


    ReadOwnParams (me; ent : mutable FlowLineSpec;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : FlowLineSpec;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : FlowLineSpec;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a FlowLineSpec <ent>, from
    --           its specific (own) parameters

    DirChecker (me; ent : FlowLineSpec) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : FlowLineSpec;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : FlowLineSpec; entto : mutable FlowLineSpec;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : FlowLineSpec;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolFlowLineSpec;
