-- Created on: 1993-02-22
-- Created by: Philippe DAUTRY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Axis2Placement from PGeom inherits AxisPlacement from PGeom

	---Purpose : This class describes an  axis two placement built
	--         with a point and two directions.
	--          
	---See Also : Axis2Placement from Geom.

uses Ax1      from gp,
     Dir      from gp

is


  Create returns Axis2Placement from PGeom;
        ---Purpose : Returns an Axis2Placement with default values.
    	---Level: Internal 


  Create (aAxis : Ax1 from gp; aXDirection: Dir from gp)
    returns Axis2Placement from PGeom;
        ---Purpose : Creates an Axis2Placement with <A2>.
    	---Level: Internal 


  XDirection (me : mutable; aXDirection : Dir from gp);
        ---Purpose : Set the value of the field xDirection with <aXDirection>.
    	---Level: Internal 


  XDirection (me) returns Dir from gp;
   	---Purpose : Returns the "XDirection". This is a unit vector.
    	---Level: Internal 


fields

  xDirection : Dir from gp;

end;
