-- File:	StepAP203_CcDesignApproval.cdl
-- Created:	Fri Nov 26 16:26:31 1999 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0
-- Copyright:	Matra Datavision 1999

class CcDesignApproval from StepAP203
inherits ApprovalAssignment from StepBasic

    ---Purpose: Representation of STEP entity CcDesignApproval

uses
    Approval from StepBasic,
    HArray1OfApprovedItem from StepAP203

is
    Create returns CcDesignApproval from StepAP203;
	---Purpose: Empty constructor

    Init (me: mutable; aApprovalAssignment_AssignedApproval: Approval from StepBasic;
                       aItems: HArray1OfApprovedItem from StepAP203);
	---Purpose: Initialize all fields (own and inherited)

    Items (me) returns HArray1OfApprovedItem from StepAP203;
	---Purpose: Returns field Items
    SetItems (me: mutable; Items: HArray1OfApprovedItem from StepAP203);
	---Purpose: Set field Items

fields
    theItems: HArray1OfApprovedItem from StepAP203;

end CcDesignApproval;
