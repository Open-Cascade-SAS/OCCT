-- Created on: 1993-11-10
-- Created by: Laurent BOURESCHE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class StripeMap from ChFiDS 

	---Purpose: 

uses 
     IndexedDataMapOfVertexListOfStripe from ChFiDS,
     Vertex from TopoDS,
     ListOfStripe from ChFiDS,
     Stripe from ChFiDS
is

    Create returns StripeMap from ChFiDS;

    Add(me : in out; V : Vertex from TopoDS; F : Stripe from ChFiDS) 
    is static;
    
    
    Extent(me) returns Integer
    ---C++: inline
    is static;
    
    FindFromKey(me; V: Vertex from TopoDS) 
    returns ListOfStripe from ChFiDS 
    ---C++: alias operator()
    ---C++: return const &
    is static;
    
    FindFromIndex(me; I : Integer from Standard) 
    returns ListOfStripe from ChFiDS
    ---C++: alias operator()
    ---C++: return const &
    is static;


    FindKey(me; I : Integer from Standard) returns Vertex  from TopoDS
    ---C++: inline
    ---C++: return const &
    is static;


    Clear(me : in out) is static;


fields

 mymap : IndexedDataMapOfVertexListOfStripe from ChFiDS;

end StripeMap;
