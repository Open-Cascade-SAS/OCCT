-- Created on: 1993-08-24
-- Created by: Bruno DUMORTIER
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Torus from ProjLib inherits Projector from ProjLib

	---Purpose: Projects elementary curves on a torus.

uses
    CurveType  from GeomAbs,
    Torus      from gp,
    Lin        	   from gp,
    Circ       	   from gp,
    Elips      	   from gp,
    Parab      	   from gp,
    Hypr       	   from gp,
    Lin2d      from gp,
    Circ2d     from gp,
    Elips2d    from gp,
    Parab2d    from gp,
    Hypr2d     from gp

raises
    NoSuchObject from Standard

is

    Create returns Torus from ProjLib;
	---Purpose: Undefined projection.

    Create(To : Torus from gp) returns Torus from ProjLib;
	---Purpose: Projection on the torus <To>.

    Create(To : Torus  from gp;
           C  : Circ from gp) returns Torus from ProjLib;
	---Purpose: Projection of the circle <C> on the torus <To>.



    Init(me : in out;
    	 To : Torus from gp)
    is static;
	 
     Project(me : in out;
     	     L  : Lin from gp)
     is redefined;
 
    Project(me : in out;
    	    C  : Circ from gp)
    is redefined;

     Project(me : in out;
     	     E  : Elips from gp)
     is redefined;
 
     Project(me : in out;
     	     P  : Parab from gp)
     is redefined;
 
     Project(me : in out;
     	     H  : Hypr from gp)
     is redefined;
	     

fields

    myTorus : Torus from gp;

end Torus;
