-- Created on: 1999-07-19
-- Created by: Denis PASCAL
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



deferred class Driver from TFunction inherits TShared from MMgt 

    ---Purpose: This  driver  class provide  services  around function
    --          execution.   One instance of  this class is  built for
    --          the whole  session.    The driver  is bound   to   the
    --          DriverGUID in the DriverTable class.
    --          It allows you to create classes which inherit from
    --          this abstract class.
    --          These subclasses identify the various algorithms
    --          which can be applied to the data contained in the
    --          attributes of sub-labels of a model.
    --          A single instance of this class and each of its
    --          subclasses is built for the whole session.
uses 
  
     Logbook   from TFunction,  
     Label     from TDF,
     LabelList from TDF
      
is 
 
    Initialize returns mutable Driver from TFunction; 


    ---Purpose: initialisation of the driver
    --          ============================

    Init(me : mutable; L : Label from TDF);
    	---Purpose: Initializes the label L for this function prior to its  execution.
     
    Label(me) returns Label from TDF;  
        ---C++: inline
        ---Purpose: Returns the label of the driver for this function.

    Validate(me; log : in out Logbook from TFunction)
    is virtual;
    	---Purpose: Validates labels of a function  in <log>. 
    	-- This function is the one initialized in this function driver.
    	-- Warning
    	-- In regeneration mode, the solver must call this
    	-- method even if the function is not executed. 
     
     
    ---Purpose: execution of function
    --          =====================

    MustExecute (me; log : Logbook from TFunction)
    	---Purpose: Analyzes the labels in the logbook log.
    	-- Returns true if attributes have been modified.
    	-- If the function label itself has been modified, the function must be executed.
    returns Boolean from Standard
    is virtual;

    Execute (me; log : in out Logbook from TFunction)
    	---Purpose: Executes the function in this function driver and
    	-- puts the impacted labels in the logbook log.
    returns Integer from Standard
    is deferred;
 
 
    ---Purpose: arguments & results of functions
    --          ================================
 
    Arguments (me; args : out LabelList from TDF)
    ---Purpose: The method fills-in the list by labels, 
    --          where the arguments of the function are located.
    is virtual;
 
    Results (me; res : out LabelList from TDF)
    ---Purpose: The method fills-in the list by labels,
    --          where the results of the function are located.
    is virtual;
 
fields 
 
    myLabel : Label from TDF;

end Driver;    
