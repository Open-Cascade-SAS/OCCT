-- Created on: 1991-01-10
-- Created by: Arnaud BOUZY
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


deferred class NamedExpression from Expr
    
inherits GeneralExpression from Expr  

    ---Purpose: Describe an expression used  by its name (as constants 
    --          or variables). A single reference is made to a 
    --          NamedExpression in every Expression (i.e. a 
    --          NamedExpression is shared).

uses AsciiString from TCollection


is

    GetName(me)
    returns AsciiString
    ---C++: return const &
    ---Level: Advanced
    is static;

    SetName(me : mutable; name : AsciiString)
    ---Level: Internal
    is static;

    IsShareable(me)
    ---Purpose: Tests if <me> can be shared by one or more expressions 
    --          or must be copied. This method redefines to a True 
    --          value the GeneralExpression method.
    returns Boolean
    is redefined;
    
    IsIdentical(me; Other : GeneralExpression)
    ---Purpose: Tests if <me> and <Other> define the same expression.
    --          This method does not include any simplification before
    --          testing.
    returns Boolean;

    String(me)
    ---Purpose: returns a string representing <me> in a readable way.
    returns AsciiString from TCollection;

fields

    myName : AsciiString;

end NamedExpression;
