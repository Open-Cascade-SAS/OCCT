-- Created on: 1994-03-03
-- Created by: Jean Louis FRENKEL
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package TColQuantity 

---Purpose: the  classes of this package should be used
--          when exporting arrays of real representing lengths, 
--          for having benefit of the unit conversion.
uses

    TCollection,
    Quantity
    
is
    class Array1OfLength instantiates Array1 from TCollection (Length from Quantity);
    class Array2OfLength instantiates Array2 from TCollection (Length from Quantity);
    class HArray1OfLength        instantiates 
    	HArray1 from TCollection  (Length from Quantity, Array1OfLength from TColQuantity); 
    class HArray2OfLength        instantiates 
    	HArray2 from TCollection  (Length from Quantity, Array2OfLength from TColQuantity); 
end TColQuantity;
