-- Created on: 1997-02-18
-- Created by: Alexander BRIVIN
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package VrmlConverter 

        ---Purpose:
        -- Computes different kinds of presentation and converts CasCade objects 
        -- ( points, curves, surfaces, shapes ... ) into nodes of VRML format 
        -- ( package Vrml ), into specific geometry shapes ( AsciiText, Cone, 
        -- IndexedFaceSet, IndexedLineSet, .... ) for requested (or default) properties 
        -- of the geometry and its appearance ( Material, Normal, Texture2, ... ) 
        -- and requested (or default)  properties of cameras and lights ( OrthograpicCamera, 
        -- PerspectiveCamera, DirectionalLight, SpotLight ).

        -- All requested properties of a current representation are specified
        -- in aDrawer of Drawer class, which qualifies how the presentation 
        -- algorithms compute the presentation of a specific kind of object. 
        -- This includes for example color, maximal chordial deviation, etc... with default values.

        -- In the result the  classes of this package Add a corresponding VRML 
        -- description to anOStream.

uses
 
        Vrml,
        Aspect, 
	Poly, 
        TColgp, 
    	MMgt,
	Adaptor3d,
        BRepAdaptor,
	TopoDS,
        HLRAlgo,
        Quantity, 
	TopTools

is
 
       	---Category: Aspect classes.
	-- The aspect classes qualifies how to represent
	-- a given kind of object.

 
    class  Drawer;
	---Purpose: qualifies the aspect properties for  
	--          the VRML conversation of a specific kind of object. 
	--          This includes for example color,  maximal chordial deviation, etc...

    class  ShadingAspect; 
	---Purpose: qualifies the aspect properties for  
	--          the VRML conversation of  a ShadedShape. 

    class  LineAspect; 
	---Purpose: qualifies the aspect properties for  
	--          the VRML conversation of a Curve and  a  DeflectionCurve . 

    class  IsoAspect; 
	---Purpose: qualifies the aspect properties for  
	--          the VRML conversation of iso curves . 

    class  PointAspect; 
	---Purpose: qualifies the aspect properties for  
	--          the VRML conversation of a Point Set . 
      


       	---Category: Presentation classes.
       	---Purpose:  To compute different kinds of presentation, to convert 
       	--           CasCade objects into VRML objects for requested aspect 
       	--           properties  and to add the  results to the stream. 


   class ShadedShape; 
    	---Purpose:  computes  the  shading presentation of shapes
    	--           by triangulation algorithms. 
 
  
   class Curve;
   	---Purpose: computes the presentation of objects to be
	--          seen as curves. The computation will be made
	--          whith a constant number of points.

   class DeflectionCurve;		      
	---Purpose: computes the presentation of objects to be seen as
	--          curves. The  computation will be made  according to
	--          a maximal chordial deviation.

	     
   class WFRestrictedFace; 
	---Purpose: computes the wireframe presentation of faces with
	--          restrictions by displaying a given number of U and/or
	--          V isoparametric curves. The isoparametric curves are
	--          drawn with a fixed number of points.


   class WFDeflectionRestrictedFace;
	---Purpose: computes the wireframe presentation of faces with
	--          restrictions by displaying a given number of U and/or
	--          V isoparametric curves. The isoparametric curves are
	--          drawn with respect to a maximal chordial deviation.


   class WFShape;  
   	---Purpose: computes the wireframe presentation of compound set 
   	--          of  faces,  edges  and vertices by displaying a given  
   	--          number of U and/or V isoparametric curves.
  

   class WFDeflectionShape;  
    	---Purpose: computes the wireframe presentation of compound 
    	--          set  of faces,  edges and vertices by displaying 
    	--          a given number of U and/or V isoparametric  curves.
      

   class HLRShape;
        ---Purpose: computes the presentation of objects with
	--          removal of their hidden lines for a specific
	--          projector.
	
   class Projector;
	---Purpose: defines the projection parameters for the hidden
	--          lines removal algorithm  and calculates properties of cameras  
    	--          and lights from Vrml ( OrthograpicCamera, PerspectiveCamera,  
    	--          DirectionalLight, PointLight, SpotLight )  
    	--          to display all shapes of scene with  arbitrary locations 
	--          for requested the Projection Vector .

 
    -- Enumeration for cameras  and  lights  from  Vrml 

   enumeration TypeOfCamera  
     is  	  
         NoCamera,
         PerspectiveCamera,
         OrthographicCamera
     end TypeOfCamera;

   enumeration TypeOfLight 
     is  	  
         NoLight,
         DirectionLight,
         PointLight,
         SpotLight
     end TypeOfLight;
       
end VrmlConverter;
