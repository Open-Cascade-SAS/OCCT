-- Created on: 1997-12-09
-- Created by: Jean-Louis Frenkel
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


private deferred class ReadWriter from PCDM inherits Transient from Standard

uses
    ExtendedString from TCollection,  
    AsciiString from TCollection, 
    Data from Storage, 
    Document from CDM, 
    MessageDriver from CDM,
    SequenceOfExtendedString from TColStd,  
    BaseDriver from Storage,  
    OpenMode from Storage, 
    SequenceOfReference from PCDM

is

    
    Version(me) returns AsciiString from TCollection
    is deferred;
    ---Purpose: returns PCDM_ReadWriter_1.
    
    WriteReferenceCounter(me; aData: mutable Data from Storage; aDocument: Document from CDM)
    is deferred;
    
    WriteReferences(me; aData: mutable Data from Storage; aDocument: Document from CDM; theReferencerFileName: ExtendedString from TCollection)
    is deferred;

    
    WriteExtensions(me; aData: mutable Data from Storage; aDocument: Document from CDM)
    is deferred;

    
    WriteVersion(me; aData: mutable Data from Storage; aDocument: Document from CDM)
    is deferred;

    
    ReadReferenceCounter(me; theFileName: ExtendedString from TCollection;   
			     theMsgDriver: MessageDriver from CDM)
    returns Integer from Standard
    is deferred;

    ReadReferences(me; aFileName: ExtendedString from TCollection; theReferences: in out  SequenceOfReference from PCDM; theMsgDriver: MessageDriver from CDM)
    is deferred;

    ReadExtensions(me; aFileName: ExtendedString from TCollection; theExtensions: in out  SequenceOfExtendedString from TColStd; theMsgDriver: MessageDriver from CDM)
    is deferred;
    
    ReadDocumentVersion(me; aFileName: ExtendedString from TCollection; theMsgDriver: MessageDriver from CDM)
    returns Integer from Standard
    is deferred;

---Category: commom methods


    Open(myclass; aDriver: in out BaseDriver from Storage; aFileName: ExtendedString from TCollection; anOpenMode: OpenMode from  Storage);
    
    Reader(myclass; aFileName: ExtendedString from TCollection)
    returns ReadWriter from PCDM;
    ---Purpose: returns the convenient Reader for a File.
    --          
    
    Writer(myclass)
    returns ReadWriter from PCDM;
    

    WriteFileFormat(myclass; aData: mutable Data from Storage; aDocument: Document from CDM);
    
    FileFormat(myclass; aFileName: ExtendedString from TCollection)
    returns ExtendedString from TCollection;
    ---Purpose: tries  to get a format  in the  file.  returns an empty
    --          string if the file could not be read or does not have 
    --          a FileFormat information.
end ReadWriter from PCDM;
