-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SurfaceCurve from StepGeom 

inherits Curve from StepGeom 

uses

	HArray1OfPcurveOrSurface from StepGeom, 
	PreferredSurfaceCurveRepresentation from StepGeom, 
	PcurveOrSurface from StepGeom, 
	HAsciiString from TCollection
is

	Create returns mutable SurfaceCurve;
	---Purpose: Returns a SurfaceCurve


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aCurve3d : mutable Curve from StepGeom;
	      aAssociatedGeometry : mutable HArray1OfPcurveOrSurface from StepGeom;
	      aMasterRepresentation : PreferredSurfaceCurveRepresentation from StepGeom) is virtual;

	-- Specific Methods for Field Data Access --

	SetCurve3d(me : mutable; aCurve3d : mutable Curve);
	Curve3d (me) returns mutable Curve;
	SetAssociatedGeometry(me : mutable; aAssociatedGeometry : mutable HArray1OfPcurveOrSurface);
	AssociatedGeometry (me) returns mutable HArray1OfPcurveOrSurface;
	AssociatedGeometryValue (me; num : Integer) returns PcurveOrSurface;
	NbAssociatedGeometry (me) returns Integer;
	SetMasterRepresentation(me : mutable; aMasterRepresentation : PreferredSurfaceCurveRepresentation);
	MasterRepresentation (me) returns PreferredSurfaceCurveRepresentation;

fields

	curve3d : Curve from StepGeom;
	associatedGeometry : HArray1OfPcurveOrSurface from StepGeom; -- a SelectType
	masterRepresentation : PreferredSurfaceCurveRepresentation from StepGeom; -- an Enumeration

end SurfaceCurve;
