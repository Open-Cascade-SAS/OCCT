-- Created on: 1996-09-17
-- Created by: Odile Olivier
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ShapeTypeFilter from StdSelect inherits Filter from SelectMgr

	--- Purpose: A filter framework which allows you to define a filter
    	-- for a specific shape type. The types available include:
    	-- -   compound
    	-- -   compsolid
    	-- -   solid
    	-- -   shell
	-- -   face
    	-- -   wire
    	-- -   edge
    	-- -   vertex.

uses
    Shape from TopoDS,
    EntityOwner from SelectMgr,
    ShapeEnum from TopAbs
is

    Create (aType: ShapeEnum from TopAbs)
    returns ShapeTypeFilter from StdSelect;
    	---Purpose: Constructs a filter object defined by the shape type aType.
    
    IsOk (me;anobj : EntityOwner from SelectMgr) 
    returns Boolean from Standard is redefined virtual;

    Type(me) returns ShapeEnum from TopAbs;
    	---Purpose: Returns the type of shape selected by the filter.
    	---C++: inline

    ActsOn(me; aStandardMode : ShapeEnum from TopAbs)
    returns Boolean from Standard is redefined virtual;

fields

    myType : ShapeEnum from TopAbs;

end ShapeTypeFilter;
