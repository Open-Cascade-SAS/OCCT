-- Created on: 2002-12-12
-- Created by: data exchange team
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class AnalysisItemWithinRepresentation from StepElement
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity AnalysisItemWithinRepresentation

uses
    HAsciiString from TCollection,
    RepresentationItem from StepRepr,
    Representation from StepRepr

is
    Create returns AnalysisItemWithinRepresentation from StepElement;
	---Purpose: Empty constructor

    Init (me: mutable; aName: HAsciiString from TCollection;
                       aDescription: HAsciiString from TCollection;
                       aItem: RepresentationItem from StepRepr;
                       aRep: Representation from StepRepr);
	---Purpose: Initialize all fields (own and inherited)

    Name (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Name
    SetName (me: mutable; Name: HAsciiString from TCollection);
	---Purpose: Set field Name

    Description (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Description
    SetDescription (me: mutable; Description: HAsciiString from TCollection);
	---Purpose: Set field Description

    Item (me) returns RepresentationItem from StepRepr;
	---Purpose: Returns field Item
    SetItem (me: mutable; Item: RepresentationItem from StepRepr);
	---Purpose: Set field Item

    Rep (me) returns Representation from StepRepr;
	---Purpose: Returns field Rep
    SetRep (me: mutable; Rep: Representation from StepRepr);
	---Purpose: Set field Rep

fields
    theName: HAsciiString from TCollection;
    theDescription: HAsciiString from TCollection;
    theItem: RepresentationItem from StepRepr;
    theRep: Representation from StepRepr;

end AnalysisItemWithinRepresentation;
