-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PresentationStyleSelect from StepVisual inherits SelectType from StepData

	-- <PresentationStyleSelect> is an EXPRESS Select Type construct translation.
	-- it gathers : PointStyle, CurveStyle, SurfaceStyleUsage, SymbolStyle, FillAreaStyle, TextStyle
	-- Rev4 : only remain PointStyle, CurveStyle, SurfaceStyleUsage

uses

	PointStyle,
	CurveStyle,
	SurfaceStyleUsage
--	SymbolStyle,
--	FillAreaStyle,
--	TextStyle
is

	Create returns PresentationStyleSelect;
	---Purpose : Returns a PresentationStyleSelect SelectType

	CaseNum (me; ent : Transient) returns Integer;
	---Purpose: Recognizes a PresentationStyleSelect Kind Entity that is :
	--        1 -> PointStyle
	--        2 -> CurveStyle
	--        3 -> SurfaceStyleUsage
	--        4 -> SymbolStyle
	--        5 -> FillAreaStyle
	--        6 -> TextStyle
	--        0 else

	PointStyle (me) returns any PointStyle;
	---Purpose : returns Value as a PointStyle (Null if another type)

	CurveStyle (me) returns any CurveStyle;
	---Purpose : returns Value as a CurveStyle (Null if another type)

	SurfaceStyleUsage (me) returns any SurfaceStyleUsage;
	---Purpose : returns Value as a SurfaceStyleUsage (Null if another type)

end PresentationStyleSelect;

