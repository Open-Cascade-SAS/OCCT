-- Created on: 2003-08-22
-- Created by: Sergey KUUL
-- Copyright (c) 2003-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class GeoTolAndGeoTolWthDatRefAndModGeoTolAndPosTol from StepDimTol
    	    	    	inherits GeometricTolerance from StepDimTol
			
uses
    HAsciiString from TCollection,
    MeasureWithUnit from StepBasic,
    ShapeAspect from StepRepr,
    GeometricToleranceWithDatumReference from StepDimTol,
    ModifiedGeometricTolerance from StepDimTol,
    PositionTolerance from StepDimTol
    
is

    Create returns mutable GeoTolAndGeoTolWthDatRefAndModGeoTolAndPosTol;
    
    Init (me: mutable; aName: HAsciiString from TCollection;
    		       aDescription: HAsciiString from TCollection;
		       aMagnitude: MeasureWithUnit from StepBasic;
		       aTolerancedShapeAspect: ShapeAspect from StepRepr;
		       aGTWDR : GeometricToleranceWithDatumReference;
		       aMGT : ModifiedGeometricTolerance);


    SetGeometricToleranceWithDatumReference(me: mutable; aGTWDR : GeometricToleranceWithDatumReference);
    
    GetGeometricToleranceWithDatumReference(me) returns mutable GeometricToleranceWithDatumReference;
    
    SetModifiedGeometricTolerance(me: mutable; aMGT : ModifiedGeometricTolerance);
    
    GetModifiedGeometricTolerance(me) returns mutable ModifiedGeometricTolerance;
    
    SetPositionTolerance(me: mutable; aPT : PositionTolerance);
    
    GetPositionTolerance(me) returns mutable PositionTolerance;
    
fields

    myGeometricToleranceWithDatumReference : GeometricToleranceWithDatumReference;
    myModifiedGeometricTolerance : ModifiedGeometricTolerance;
    myPositionTolerance : PositionTolerance;
    
end GeoTolAndGeoTolWthDatRefAndModGeoTolAndPosTol;
