-- Created on: 1995-10-20
-- Created by: Yves FRICAUD
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Interval from BRepOffset 

	---Purpose: 

uses
    Type from BRepOffset
    
is

    Create;
    
    Create (U1,U2 : Real from Standard;
    	    Type  : Type from BRepOffset)
    returns Interval from BRepOffset;
    
    First (me : in out; U : Real from Standard)
    	---C++: inline
    is static;
    
    Last  (me : in out; U : Real from Standard)
        ---C++: inline
    is static;    
    
    Type  (me : in out; T : Type from BRepOffset)
       ---C++: inline
    is static;
    
    First (me) returns Real from Standard
       ---C++: inline
    is static;    
    
    Last  (me) returns Real from Standard
       ---C++: inline
    is static;
    
    Type  (me) returns Type from BRepOffset
       ---C++: inline
    is static;    
    

fields

    f,l  : Real from Standard;
    type : Type from BRepOffset;
    
end Interval;
