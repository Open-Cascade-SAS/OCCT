-- Created by: DAUTRY Philippe
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

--      	-----------------------------

---Version:	0.0
--Version	Date		Purpose
--		0.0	Oct 10 1997	Creation


class DefaultDeltaOnRemoval from TDF
    inherits DeltaOnRemoval from TDF

	---Purpose: This class provides a default implementation of a
	--          TDF_DeltaOnRemoval.

uses

    Label     from TDF,
    Attribute from TDF
    
-- raises

is

    Create(anAttribute : Attribute from TDF);
	---Purpose: Creates a TDF_DefaultDeltaOnRemoval.

    Apply (me : mutable)
    	is redefined virtual;
    	---Purpose: Applies the delta to the attribute.

end DefaultDeltaOnRemoval;
