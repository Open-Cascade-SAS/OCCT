-- Created by: Peter KURNEV
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Tools from BOPAlgo 

---Purpose: 

uses  
    BaseAllocator from BOPCol, 
    IndexedDataMapOfIntegerListOfInteger from BOPCol,  
    DataMapOfIntegerListOfInteger from BOPCol, 
    PDS from BOPDS, 
    PaveBlock from BOPDS,  
    IndexedDataMapOfPaveBlockListOfInteger from BOPDS, 
    IndexedDataMapOfPaveBlockListOfPaveBlock from BOPDS, 
    DataMapOfIntegerListOfPaveBlock from BOPDS
--raises

is
    --- 
    --- static methods 
    --- 
    MakeBlocksCnx(myclass; 
        theMILI     :IndexedDataMapOfIntegerListOfInteger from BOPCol; 
        theMBlocks  :out DataMapOfIntegerListOfInteger from BOPCol; 
        theAllocator:out BaseAllocator from BOPCol);  

    MakeBlocks(myclass; 
        theMILI     :IndexedDataMapOfPaveBlockListOfPaveBlock from BOPDS; 
        theMBlocks  :out DataMapOfIntegerListOfPaveBlock from BOPDS; 
        theAllocator:out BaseAllocator from BOPCol); 
 
    PerformCommonBlocks(myclass; 
        theMBlocks  :out IndexedDataMapOfPaveBlockListOfPaveBlock from BOPDS; 
        theAllocator:out BaseAllocator from BOPCol; 
        pDS: out PDS from BOPDS);
    
    FillMap(myclass; 
        tneN1:Integer from Standard; 
        tneN2:Integer from Standard; 
        theMILI : out IndexedDataMapOfIntegerListOfInteger from BOPCol; 
        theAllocator: out BaseAllocator from BOPCol); 
    
     
    FillMap(myclass; 
        tnePB1:PaveBlock from BOPDS; 
        tnePB2:PaveBlock from BOPDS; 
        theMILI : out IndexedDataMapOfPaveBlockListOfPaveBlock from BOPDS; 
        theAllocator: out BaseAllocator from BOPCol);
 
    FillMap(myclass; 
        tnePB1:PaveBlock from BOPDS; 
        tneF:Integer from Standard;  
        theMILI : out IndexedDataMapOfPaveBlockListOfInteger from BOPDS; 
        theAllocator: out BaseAllocator from BOPCol); 
 
    PerformCommonBlocks(myclass; 
        theMBlocks  :IndexedDataMapOfPaveBlockListOfInteger from BOPDS; 
        theAllocator:out BaseAllocator from BOPCol; 
        pDS: out PDS from BOPDS);
--fields

end Tools;
