-- Created on: 1997-10-07
-- Created by: Laurent BUCHARD
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Tool from BRepTopAdaptor 

uses 
    Face       from TopoDS,
    TopolTool  from BRepTopAdaptor,
    HSurface   from Adaptor3d


is 

  Create
     returns Tool from BRepTopAdaptor;

  Create(F     : Face from TopoDS;
    	 Tol2d : Real from Standard)
     returns Tool from BRepTopAdaptor;
     
  Create(Surface: HSurface from Adaptor3d;
         Tol2d  : Real from Standard)
     returns Tool from BRepTopAdaptor;
 
 
  Init(me    : in out;
       F     : Face from TopoDS;
       Tol2d : Real from Standard);
       
  Init(me     : in out;
       Surface: HSurface from Adaptor3d;
       Tol2d  : Real from Standard);       
	  
  ---- 

  GetTopolTool(me: in out) 
     returns TopolTool from BRepTopAdaptor;
     
  SetTopolTool(me: in out ; 
               TT: TopolTool from BRepTopAdaptor);
	
  GetSurface(me: in out)
    returns HSurface from Adaptor3d;
    
	
  ---
	
  Destroy(me: in out) ;
    ---C++: alias ~
    
fields

  myloaded    : Boolean   from Standard;
  myTopolTool : TopolTool from BRepTopAdaptor; 
  myHSurface  : HSurface  from Adaptor3d;

end Tool;
