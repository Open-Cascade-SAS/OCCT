-- Created on: 1995-08-07
-- Created by: Modelistation
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class WFDeflectionRestrictedFace from StdPrs
	  
inherits Root from Prs3d
	 

	---Purpose: A framework to provide display of U and V
    	-- isoparameters of faces, while allowing you to impose
    	-- a deflection on them.

uses
    HSurface             from BRepAdaptor,
    Presentation         from Prs3d,
    Drawer               from Prs3d,
    Length               from Quantity, 
    NListOfSequenceOfPnt from Prs3d

    
is
    Add(myclass; aPresentation: Presentation from Prs3d; 
        	 aFace        : HSurface     from BRepAdaptor;
    	    	 aDrawer      : Drawer       from Prs3d);
	---Purpose: Defines a display featuring U and V isoparameters.
    	-- Adds the surface aFace to the
    	-- StdPrs_WFRestrictedFace algorithm. This face is
    	-- found in a shape in the presentation object
    	-- aPresentation, and its display attributes - in
    	-- particular, the number of U and V isoparameters - are
    	-- set in the attribute manager aDrawer.
    	-- aFace is BRepAdaptor_HSurface surface created
    	-- from a face in a topological shape.   which is passed
    	-- as an argument through the
    	-- BRepAdaptor_HSurface surface created from it.
    	-- This is what allows the topological face to be treated
    	-- as a geometric surface.	 
    
    AddUIso(myclass; aPresentation: Presentation from Prs3d; 
        	     aFace        : HSurface     from BRepAdaptor;
    	    	     aDrawer      : Drawer       from Prs3d);
    	---Purpose:	Defines a display featuring U isoparameters
    	-- respectively. Add the surface aFace to the
    	-- StdPrs_WFRestrictedFace algorithm. This face
    	-- is found in a shape in the presentation object
    	-- aPresentation, and its display attributes - in
    	-- particular, the number of U isoparameters -
    	-- are set in the attribute manager aDrawer.
    	-- aFace is BRepAdaptor_HSurface surface
    	-- created from a face in a topological shape.   which
    	-- is passed to the function as an argument through
    	-- the BRepAdaptor_HSurface surface created from
    	-- it. This is what allows the topological face to be
    	-- treated as a geometric surface.
        
    AddVIso(myclass; aPresentation: Presentation from Prs3d; 
        	     aFace        : HSurface     from BRepAdaptor;
    	    	     aDrawer      : Drawer       from Prs3d);
    	---Purpose:	Defines a display featuring V isoparameters
    	-- respectively. Add the surface aFace to the
    	-- StdPrs_WFRestrictedFace algorithm. This face
    	-- is found in a shape in the presentation object
    	-- aPresentation, and its display attributes - in
    	-- particular, the number of V isoparameters -
    	-- are set in the attribute manager aDrawer.
    	-- aFace is BRepAdaptor_HSurface surface
    	-- created from a face in a topological shape.   which
    	-- is passed to the function as an argument through
    	-- the BRepAdaptor_HSurface surface created from
    	-- it. This is what allows the topological face to be
    	-- treated as a geometric surface.
    
    Add(myclass;  aPresentation: Presentation from Prs3d; 
    	          aFace        : HSurface     from BRepAdaptor;
		  DrawUIso, DrawVIso: Boolean from Standard;
		  Deflection   : Length       from Quantity;
		  NBUiso,NBViso: Integer      from Standard;
		  aDrawer      : Drawer       from Prs3d; 
    	    	  Curves       : out NListOfSequenceOfPnt from Prs3d);
	---Purpose: Defines a display of a delection-specified face. The
    	-- display will feature U and V isoparameters.
    	-- Adds the topology aShape to the
    	-- StdPrs_WFRestrictedFace algorithm. This shape is
    	-- found in the presentation object aPresentation, and
    	-- its display attributes - except the number of U and V
    	-- isoparameters - are set in the attribute manager aDrawer.
    	-- The function sets the number of U and V
    	-- isoparameters, NBUiso and NBViso, in the shape. To
    	-- do this, the arguments DrawUIso and DrawVIso must be true.
    	-- aFace is BRepAdaptor_HSurface surface created
    	-- from a face in a topological shape.   which is passed
    	-- as an argument through the
    	-- BRepAdaptor_HSurface surface created from it.
    	-- This is what allows the topological face to be treated
    	-- as a geometric surface.  
	-- Curves give a sequence of face curves, it is used if the PrimitiveArray  
        -- visualization approach is activated (it is activated by default).
        
    Match(myclass; X,Y,Z    : Length   from Quantity;
                   aDistance: Length   from Quantity;
        	   aFace    : HSurface from BRepAdaptor;
    	    	   aDrawer  : Drawer   from Prs3d)
    returns Boolean from Standard;
		 
    MatchUIso(myclass; X,Y,Z    : Length   from Quantity;
                       aDistance: Length   from Quantity;
        	       aFace    : HSurface from BRepAdaptor;
    	    	       aDrawer  : Drawer   from Prs3d)
    returns Boolean from Standard;
		 
    MatchVIso(myclass; X,Y,Z    : Length   from Quantity;
                       aDistance: Length   from Quantity;
         	       aFace    : HSurface from BRepAdaptor;
    	    	       aDrawer  : Drawer   from Prs3d)
    returns Boolean from Standard;
		 

    Match(myclass;X,Y,Z        : Length       from Quantity;
                  aDistance    : Length       from Quantity;
    	          aFace        : HSurface     from BRepAdaptor; 
    	    	  aDrawer      : Drawer       from Prs3d;
		  DrawUIso, DrawVIso: Boolean from Standard;
		  aDeflection  : Length       from Quantity;
		  NBUiso,NBViso: Integer      from Standard)

    returns Boolean from Standard;	  
		   
end WFDeflectionRestrictedFace;

