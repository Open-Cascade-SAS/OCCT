-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ContextDependentInvisibility from StepVisual 

inherits Invisibility from StepVisual 

uses

	InvisibilityContext from StepVisual, 
	HArray1OfInvisibleItem from StepVisual
is

	Create returns mutable ContextDependentInvisibility;
	---Purpose: Returns a ContextDependentInvisibility


	Init (me : mutable;
	      aInvisibleItems : mutable HArray1OfInvisibleItem from StepVisual) is redefined;

	Init (me : mutable;
	      aInvisibleItems : mutable HArray1OfInvisibleItem from StepVisual;
	      aPresentationContext : InvisibilityContext from StepVisual) is virtual;

	-- Specific Methods for Field Data Access --

	SetPresentationContext(me : mutable; aPresentationContext : InvisibilityContext);
	PresentationContext (me) returns InvisibilityContext;

fields

	presentationContext : InvisibilityContext from StepVisual; -- a SelectType

end ContextDependentInvisibility;
