-- Created on: 2003-01-28
-- Created by: data exchange team
-- Copyright (c) 2003-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class ProductOrFormationOrDefinition from StepBasic
inherits SelectType from StepData

    ---Purpose: Representation of STEP SELECT type ProductOrFormationOrDefinition

uses
    Product from StepBasic,
    ProductDefinitionFormation from StepBasic,
    ProductDefinition from StepBasic

is
    Create returns ProductOrFormationOrDefinition from StepBasic;
	---Purpose: Empty constructor

    CaseNum (me; ent: Transient) returns Integer;
	---Purpose: Recognizes a kind of ProductOrFormationOrDefinition select type
	--          1 -> Product from StepBasic
	--          2 -> ProductDefinitionFormation from StepBasic
	--          3 -> ProductDefinition from StepBasic
	--          0 else

    Product (me) returns Product from StepBasic;
	---Purpose: Returns Value as Product (or Null if another type)

    ProductDefinitionFormation (me) returns ProductDefinitionFormation from StepBasic;
	---Purpose: Returns Value as ProductDefinitionFormation (or Null if another type)

    ProductDefinition (me) returns ProductDefinition from StepBasic;
	---Purpose: Returns Value as ProductDefinition (or Null if another type)

end ProductOrFormationOrDefinition;
