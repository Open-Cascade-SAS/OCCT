-- Created on: 1997-02-06
-- Created by: Kernel
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

private class InternalData from Storage

inherits TShared from MMgt

uses BucketOfPersistent from Storage,
     HPArray from Storage,
     MapOfCallBack from Storage         
is
    Create returns InternalData from Storage;
    
    Clear(me : mutable);
    
    fields
    
      myPtoA               : BucketOfPersistent from Storage;
      myObjId              : Integer from Standard;
      myTypeId             : Integer from Standard;
      myReadArray          : HPArray from Storage;
      myTypeBinding        : MapOfCallBack from Storage;      
      
    friends class Schema from Storage   
    
end;
