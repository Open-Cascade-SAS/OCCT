--
-- File:        AlienImage_SGIRGBAlienData.cdl
-- Created:     23/03/93
-- Author:      BBL
--
---Copyright:   Matravision 1993
--

class SGIRGBAlienData from AlienImage inherits AlienImageData from AlienImage

        ---Version: 0.0

        ---Purpose: This class defines a SGI .rgb Alien image.
        ---Keywords:
        ---Warning:
        ---References:

uses
        File                    from OSD,
        AsciiString             from TCollection,
        ColorImage              from Image,
        PseudoColorImage        from Image,
        Image                   from Image,
        X11XColor               from AlienImage,
        SGIRGBFileHeader        from AlienImage

raises
        OutOfRange      from Standard,
        TypeMismatch    from Standard

is
        Create returns mutable SGIRGBAlienData from AlienImage ;

        Clear( me : in out mutable ) ;
        ---Level: Public
        ---Purpose: Frees memory allocated by SGIRGBAlienData
        ---C++: alias ~

        Read ( me : in out mutable ; afile : in out File from OSD )
          returns Boolean from Standard ;
        ---Level: Public
          ---Purpose: Read content of a  SGIRGBAlienData object from a file .
          --          Returns True if file is a SGI .rgb file .

        Write( me : in immutable; afile : in out File from OSD )
          returns Boolean from Standard ;
        ---Level: Public
          ---Purpose: Write content of a  SGIRGBAlienData object to a file .

        SetName( me : in out mutable ;
                 aName : in AsciiString from TCollection)
        is redefined;
        ---Level: Public
          ---Purpose: Set Image name .

        Name( me : in immutable ) returns AsciiString from TCollection
        is redefined;
          ---C++: return const &
        ---Level: Public
          ---Purpose: Get Image name .

        ToImage( me : in  immutable) 
          returns mutable Image from Image 
          raises TypeMismatch from Standard ;
        ---Level: Public
          ---Purpose : convert a SGIRGBAlienData object to a Image object.

        FromImage( me : in out mutable ; anImage : in Image from Image )
          raises TypeMismatch from Standard ;
        ---Level: Public
          ---Purpose : convert a Image object to a SGIRGBAlienData object.

        --
        --                      Private Method
        --

        ToPseudoColorImage( me : in immutable) 
          returns PseudoColorImage from Image is private ;
        ---Level: Internal
          ---Purpose : convert a AlienImage object to a Image object.

        ToColorImage( me : in immutable) 
          returns ColorImage from Image is private ;
        ---Level: Internal
          ---Purpose : convert a AlienImage object to a Image object.

fields

        myHeader : SGIRGBFileHeader from AlienImage is protected ;
        myRedData, myGreenData, myBlueData : Address from Standard is protected;
                -- ( unsigned short * )

end ;
 
