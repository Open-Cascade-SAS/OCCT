-- Created on: 1999-08-02
-- Created by: Denis PASCAL
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Current from TDataStd inherits Attribute from TDF

	---Purpose: this attribute,  located at root label,  manage an
	--          access to a current label.

uses Attribute       from TDF,
     Label           from TDF,
     GUID            from Standard,
     DataSet         from TDF,
     RelocationTable from TDF

is

    ---Purpose: class methods
    --          =============


    GetID (myclass)   
    	---C++: return const &  
    returns GUID from Standard;


    Set (myclass; L : Label from TDF);   
    ---Purpose: Set <L> as current of <L> Framework.


    Get (myclass; acces : Label from TDF)    
    ---Purpose: returns current of <acces> Framework. raise if (!Has)
    returns Label from TDF;    


    Has (myclass; acces : Label from TDF)
    ---Purpose: returns True if a  current label is managed in <acces>
    --          Framework.
    returns Boolean from Standard;
    
    ---Purpose: class methods
    --          =============    

    Create
    returns Current from TDataStd;    

    SetLabel (me : mutable; current : Label from TDF);
    
    GetLabel (me)
    returns Label from TDF;

    	---Category: TDF_Attribute methods
    	--           =====================
    
    ID (me)
    	---C++: return const & 
    returns GUID from Standard;

    Restore (me: mutable; With : Attribute from TDF);

    NewEmpty (me)
    returns Attribute from TDF;

    Paste (me; Into : Attribute from TDF;
	       RT   : RelocationTable from TDF);    

    Dump(me; anOS : in out OStream from Standard)
    returns OStream from Standard
    is redefined;
    ---C++: return &


fields

    myLabel : Label from TDF;

end Current;
