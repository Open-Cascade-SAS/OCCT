-- Created on: 1991-12-13
-- Created by: Christophe MARION
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Intervals from Intrv
	---Purpose: The class  Intervals is a  sorted  sequence of non
	--          overlapping  Real Intervals.

uses
    Integer            from Standard,
    Interval           from Intrv,
    SequenceOfInterval from Intrv

raises
    OutOfRange

is
    Create returns Intervals from Intrv;
	---Purpose: Creates a void sequence of intervals.

    Create(Int : Interval from Intrv) returns Intervals from Intrv;
	---Purpose: Creates a sequence of one interval.
	
    Create(Int : Intervals from Intrv) returns Intervals from Intrv;
	---Purpose: Creates   by   copying  an   existing  sequence of
	--          intervals.
	
    Intersect(me : in out; Tool : Interval from Intrv)
	---Purpose: Intersects the intervals with the interval <Tool>.
    is static;

    Intersect(me : in out; Tool : Intervals from Intrv)
	---Purpose: Intersects the intervals with the intervals in the
	--          sequence  <Tool>.
    is static;

    Subtract(me : in out; Tool : Interval from Intrv)
    is static;

    Subtract(me : in out; Tool : Intervals from Intrv)
    is static;

    Unite(me : in out; Tool : Interval from Intrv)
    is static;

    Unite(me : in out; Tool : Intervals from Intrv)
    is static;

    XUnite(me : in out; Tool : Interval from Intrv)
    is static;

    XUnite(me : in out; Tool : Intervals from Intrv)
    is static;

    NbIntervals(me) returns Integer from Standard
    	---C++: inline
    is static;

    Value(me; Index : Integer from Standard) 
    returns Interval from Intrv
    	---C++: inline
    	---C++: return const &
    raises OutOfRange from Standard
    is static;
    
fields
    myInter : SequenceOfInterval from Intrv;

end Intervals;
