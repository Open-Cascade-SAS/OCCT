-- Created on: 1993-04-06
-- Created by: Philippe DAUTRY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Hyperbola from PGeom2d inherits Conic from PGeom2d

        ---Purpose :Defines the main branch of an hyperbola.
        --         
	---See Also : Hyperbola from Geom2d.

uses Ax22d from gp

is


  Create returns mutable Hyperbola from PGeom2d;
        ---Purpose :Creates an Hyperbola with default values.
	---Level: Internal 


  Create (aPosition : Ax22d from gp;
    	  aMajorRadius, aMinorRadius : Real from Standard)
     returns mutable Hyperbola from PGeom2d;
	---Purpose :  Creates an   Hyperbola    with      <aPosition>,
	--         <aMajorRadius> and  <aMinorRadius> as field values.
	--         The major  radius of the hyperbola is  on the XAxis
	--         and   the minor  radius is  on    the YAxis of  the
	--         hyperbola.
	---Level: Internal 


  MajorRadius (me : mutable; aMajorRadius : Real from Standard);
	---Purpose: Set the value of the field majorRadius with <aMajorRadius>.
	---Level: Internal 


  MajorRadius (me)  returns Real from Standard;
	---Purpose: Returns the value of the field majorRadius.
	---Level: Internal 


  MinorRadius (me : mutable; aMinorRadius : Real from Standard);
	---Purpose: Set the value of the field minorRadius with <aMinorRadius>.
	---Level: Internal 


  MinorRadius (me)  returns Real from Standard;
	---Purpose: Returns the value of the field minorRadius.
	---Level: Internal 


fields

     majorRadius : Real from Standard;
     minorRadius : Real from Standard;

end;

