-- File:	Extrema_FuncExtCS.cdl
-- Created:	Mon Jan 22 17:06:01 1996
-- Author:	Laurent PAINNOT
--		<lpa@nonox>
---Copyright:	 Matra Datavision 1996


private class FuncExtCS from Extrema

 inherits FunctionSetWithDerivatives from math
    ---Purpose: Fonction permettant de rechercher les extrema de la 
    --          distance entre une courbe et une surface.

uses    POnSurf           from Extrema,
    	POnCurv           from Extrema,
	SequenceOfPOnSurf from Extrema,
	SequenceOfPOnCurv from Extrema,
	SequenceOfReal    from TColStd,
	Pnt               from gp,
	Vector            from math,
	Matrix            from math,
	Curve             from Adaptor3d,
    	CurvePtr          from Adaptor3d,
	Surface           from Adaptor3d,
    	SurfacePtr        from Adaptor3d

raises  OutOfRange from Standard

is
    Create returns FuncExtCS;

    Create (C: Curve from Adaptor3d; S: Surface from Adaptor3d) returns FuncExtCS;
    	---Purpose:

    Initialize(me: in out; C: Curve from Adaptor3d; S: Surface from Adaptor3d)
    	---Purpose: sets the field mysurf of the function.
    is static;
    
    ------------------------------------------------------------
    -- In all next methods, an exception is raised if the fields 
    -- were not initialized.

    NbVariables (me) returns Integer;

    NbEquations (me) returns Integer;

    Value (me: in out; UV: Vector; F: out Vector) returns Boolean;
    	---Purpose: Calcul de Fi(U,V).

    Derivatives (me: in out; UV: Vector; DF: out Matrix)
    	returns Boolean;
    	---Purpose: Calcul de Fi'(U,V).

    Values (me: in out; UV: Vector; F: out Vector; DF: out Matrix)
    	returns Boolean;
    	---Purpose: Calcul de Fi(U,V) et Fi'(U,V).

    GetStateNumber (me: in out) returns Integer
    	---Purpose: Memorise l'extremum trouve.
    	is redefined;

    NbExt (me) returns Integer;
    	---Purpose: Renvoie le nombre d'extrema trouves.

    SquareDistance (me; N: Integer) returns Real
    	---Purpose: Renvoie la valeur de la Nieme distance.
    	raises  OutOfRange;
	    	-- si N < 1 ou N > NbExt(me).

    PointOnCurve (me; N: Integer) returns POnCurv
    	---Purpose: Renvoie le Nieme extremum sur C.
    	---C++: return const&
    	raises  OutOfRange;
	    	-- si N < 1 ou N > NbExt(me).

    PointOnSurface (me; N: Integer) returns POnSurf
    	---Purpose: Renvoie le Nieme extremum sur S.
    	---C++: return const&
    	raises  OutOfRange;
	    	-- si N < 1 ou N > NbExt(me).

    Bidon1(me) returns SurfacePtr from Adaptor3d
    is static private;

    Bidon2(me) returns CurvePtr from Adaptor3d
    is static private;


fields
    myC    : CurvePtr from Adaptor3d;
    myS    : SurfacePtr from Adaptor3d;
    
    myP1   : Pnt from gp;
    myP2   : Pnt from gp;

    myt    : Real;          -- valeur courante de U sur C
    myU    : Real;          -- valeur courante de U sur S
    myV    : Real;          -- valeur courante de V sur S

    mySqDist:  SequenceOfReal    from TColStd;
    myPoint1: SequenceOfPOnCurv from Extrema;
    myPoint2: SequenceOfPOnSurf from Extrema;
    
    myCinit: Boolean;
    mySinit: Boolean;

end FuncExtCS;
