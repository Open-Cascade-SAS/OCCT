-- Created on: 1994-08-30
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ShapeShapeInterference from TopOpeBRepDS 
    inherits Interference from TopOpeBRepDS

	---Purpose: Interference

uses

    Transition from TopOpeBRepDS,
    Kind       from TopOpeBRepDS,
    Config     from TopOpeBRepDS,
    OStream    from Standard    

is

    Create(T  : Transition from TopOpeBRepDS;
	   ST : Kind from TopOpeBRepDS;
	   S  : Integer from Standard;
	   GT : Kind from TopOpeBRepDS;
	   G  : Integer from Standard;
    	   GBound : Boolean from Standard;
    	   C  : Config from TopOpeBRepDS)
    
    ---Purpose: a shape interfers on shape <G> with shape <S>.
    -- examples : 
    -- create a ShapeShapeInterference describing :
    -- vertex V of edge E1 found on edge E2 :
    -- ST,S,GT,G = TopOpeBRepDS_EDGE,E2,TopOpeBRepDS_VERTEX,V
    -- 
    -- create a ShapeShapeInterference describing
    -- vertex V of edge E found on face F :
    -- ST,S,GT,G = TopOpeBRepDS_FACE,F,TopOpeBRepDS_VERTEX,V
    --
    -- <GBound> indicates if shape <G> is a bound of shape <S>.
    --     
    -- <SCC> : 
    -- UNSH_GEOMETRY : 
    -- 	 <S> and <Ancestor> have any types, 
    -- 	 <S> and <Ancestor> don't share the same geometry 
    -- SAME_ORIENTED : 
    -- 	 <S> and <Ancestor> have identical types, 
    -- 	 <S> and <Ancestor> orientations are IDENTICAL.
    -- DIFF_ORIENTED : 
    -- 	 <S> and <Ancestor> have identical types, 
    -- 	 <S> and <Ancestor> orientations are DIFFERENT.
    -- 
    returns ShapeShapeInterference from TopOpeBRepDS; 
	    
    
    Config(me) returns Config from TopOpeBRepDS
    is static;

    GBound(me) returns Boolean from Standard
    is static;

    SetGBound(me : mutable; b : Boolean from Standard)
    is static;    
        
    Dump(me; OS : in out OStream from Standard) returns OStream
    is redefined;
    ---C++: return &


fields

    myGBound : Boolean from Standard;
    myC      : Config from TopOpeBRepDS;
    
end ShapeShapeInterference from TopOpeBRepDS;
