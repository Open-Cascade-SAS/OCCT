-- Created on: 1992-05-22
-- Created by: Jean Claude VAUTHIER
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class BSplineSurface  from DrawTrSurf 

inherits Surface from DrawTrSurf

        --- Purpose :
        --  This class defines a drawable BSplineSurface. 
        --  With this class you can draw the control points and the knots 
        --  of the surface.
        --  You can use the general class Surface from DrawTrSurf too,
        --  if you just want to sea boundaries and isoparametric curves.

uses BSplineSurface from Geom,
     Color from Draw,
     MarkerShape from Draw,
     Display from Draw,
     Drawable3D from Draw

is



  Create (S : BSplineSurface from Geom)
     returns mutable BSplineSurface from DrawTrSurf;
        --- Purpose : default drawing mode.
        --  The isoparametric curves corresponding to the knots values are 
        --  drawn.
        --  The control points and the knots points are drawn.
        --  The boundaries are yellow, the isoparametric curves are blues.
        --  For the discretisation 50 points are computed in each parametric
        --  direction.


  Create (S : BSplineSurface from Geom;
          BoundsColor, IsosColor, PolesColor, KnotsColor : Color from Draw;
          KnotsShape : MarkerShape from Draw; KnotsSize : Integer;
          ShowPoles, ShowKnots : Boolean; Discret : Integer; Deflection : Real;
          DrawMode : Integer)
     returns mutable BSplineSurface from DrawTrSurf;
        --- Purpose :
        --  The isoparametric curves corresponding to the knots values are 
        --  drawn.



  Create (S : BSplineSurface from Geom;
          NbUIsos, NbVIsos : Integer;
          BoundsColor, IsosColor, PolesColor, KnotsColor : Color from Draw;
          KnotsShape : MarkerShape from Draw; KnotsSize : Integer;
          ShowPoles, ShowKnots : Boolean; Discret : Integer; Deflection : Real;
          DrawMode : Integer)
     returns mutable BSplineSurface from DrawTrSurf;
	--- Purpose : Parametric equidistant iso curves are drawn.


  DrawOn (me; dis : in out Display from Draw)
     is redefined static;


  ShowPoles  (me : mutable)
     is static;


  ShowKnots  (me : mutable)
     is static;


  ShowIsos (me : mutable; Nu, Nv : Integer)
        --- Purpose : change the number of isoparametric curves to be drawn.
     is redefined;


  ShowKnotsIsos (me : mutable)
        --- Purpose : change the number of isoparametric curves to be drawn.
     is static;


  ClearIsos (me : mutable)
        --- Purpose : rub out all the isoparametric curves.
     is redefined;
     

  ClearPoles (me : mutable)
     is static;
  

  ClearKnots (me : mutable)
     is static;


  FindPole(me; X,Y : Real; D : Display from Draw; Prec : Real; 
            UIndex, VIndex : in out Integer)
  is static;
  

  FindUKnot(me; X,Y : Real; D : Display from Draw; Prec : Real; 
            UIndex : in out Integer)
  is static;


  FindVKnot(me; X,Y : Real; D : Display from Draw; Prec : Real; 
            VIndex : in out Integer)
  is static;


  SetPolesColor (me : mutable; aColor : Color from Draw)
        ---C++: inline
     is static;


  SetKnotsColor (me : mutable; aColor : Color from Draw)
        ---C++: inline
     is static;


  SetKnotsShape (me : mutable; Shape : MarkerShape from Draw)
        ---C++: inline
     is static;


  KnotsShape (me)  returns MarkerShape from Draw
        ---C++: inline
     is static;
  

  KnotsColor (me)  returns Color from Draw
        ---C++: inline
     is static;
  

  PolesColor (me)  returns Color from Draw
        ---C++: inline
     is static;
    
  Copy(me) returns mutable Drawable3D from Draw
	---Purpose: For variable copy.
  is redefined;
	

fields

  drawPoles   : Boolean;
  drawKnots   : Boolean;
  knotsIsos   : Boolean;
  knotsForm   : MarkerShape from Draw;
  knotsLook   : Color from Draw;
  knotsDim    : Integer;
  polesLook   : Color from Draw;

end BSplineSurface;
