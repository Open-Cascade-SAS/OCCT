-- Created on: 1993-01-22
-- Created by: Gilles DEBARBOUILLE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class FuzzyDefinition from Dynamic
inherits

    FuzzyClass from Dynamic
    
	---Purpose: It  is the class  useful for  setting a particular
	--          definition   of  an   object.  This  definition is
	--          caracterized by  a  collection of parameters. Each
	--          parameter  is identified by its  name, the type of
	--          its referenced   value and if  necessary a default
	--          value.

uses

    OStream from Standard,
    CString from Standard,
    HAsciiString from TCollection,
    AsciiString  from TCollection


is

    Create(aname : CString from Standard) returns mutable FuzzyDefinition from Dynamic;
    
    ---Level: Public 
    
    ---Purpose: Creates a FuzzyDefinition with <aname> as type.
    
    Type(me) returns AsciiString from TCollection
    
    ---Level: Public 
    
    ---Purpose: Returns the type of object.
    
    is redefined;
    
    Dump(me ; astream : in out OStream from Standard)
    
    ---Level: Internal 
    
    ---Purpose: Useful for debugging.

    is redefined;
    
fields

    thename : HAsciiString from TCollection;

end FuzzyDefinition;
