-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SurfaceSideStyle from StepVisual 

inherits TShared from MMgt

uses

	HAsciiString from TCollection, 
	HArray1OfSurfaceStyleElementSelect from StepVisual, 
	SurfaceStyleElementSelect from StepVisual
is

	Create returns mutable SurfaceSideStyle;
	---Purpose: Returns a SurfaceSideStyle

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aStyles : mutable HArray1OfSurfaceStyleElementSelect from StepVisual) is virtual;

	-- Specific Methods for Field Data Access --

	SetName(me : mutable; aName : mutable HAsciiString);
	Name (me) returns mutable HAsciiString;
	SetStyles(me : mutable; aStyles : mutable HArray1OfSurfaceStyleElementSelect);
	Styles (me) returns mutable HArray1OfSurfaceStyleElementSelect;
	StylesValue (me; num : Integer) returns SurfaceStyleElementSelect;
	NbStyles (me) returns Integer;

fields

	name : HAsciiString from TCollection;
	styles : HArray1OfSurfaceStyleElementSelect from StepVisual; -- a SelectType

end SurfaceSideStyle;
