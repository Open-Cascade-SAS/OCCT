-- Created on: 1995-03-22
-- Created by: Jean-Louis  Frenkel
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

private class StoreList from CDF inherits Transient from Standard

uses
    Document from CDM,
    ListOfDocument from CDM,
    MapOfDocument from CDM,
    MapIteratorOfMapOfDocument from CDM,
    MetaData from CDM,
    ExtendedString from TCollection,
    StoreStatus from PCDM

raises NoSuchObject from Standard
is

    Create(aDocument: Document from CDM)
    returns StoreList from CDF;
    
    IsConsistent(me) returns Boolean from Standard;

    
    Store(me: mutable; aMetaData: out MetaData from CDM;
		       aStatusAssociatedText: out ExtendedString from TCollection)
    returns StoreStatus from PCDM
    ---Purpose: stores each object of the storelist in the reverse
    --          order of which they had been added.
    raises NoSuchObject from Standard;
    ---Warning: if the active dbunit cannot be found


     ---Category: Private methods.


    Add(me: mutable; aDocument: Document from CDM)
    is private;

 ---Category: iteration methods
    Init(me: mutable);
    More(me) returns Boolean from Standard;
    Next(me: mutable);
    Value(me) returns Document from CDM;
    
    
fields

    myItems: MapOfDocument from CDM;
    myStack: ListOfDocument from CDM;
    myIterator: MapIteratorOfMapOfDocument from CDM;
    myMainDocument: Document from CDM;
end StoreList from CDF;
