-- Created on: 1992-01-21
-- Created by: GG
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Update:	             		


class PerspectiveView from V3d

    	---Purpose : Creates and modifies a perspective
	--           See the methods of the class View	



inherits View from V3d


uses

	Viewer from V3d,
	OrthographicView from V3d,
	PlaneAngle from Quantity

raises

        BadValue from V3d
	
is

    	Create ( VM : mutable Viewer ) returns mutable PerspectiveView;
	---Level: Public
	---Purpose: Defines a perspective view in a viewer VM.
	--          The default angle of opening is given
	--          by the viewer.
     

    	Create ( VM : mutable Viewer ; V : OrthographicView )
					returns mutable PerspectiveView;  
	---Level: Public
	---Purpose: Creates a perspective view from the parameters 
	--	    of an orthographic view.
        --          The parameters of the original view are duplicated
        --          in the resulting view (Projection,Mapping,Context) .
        --          The view thus created must be activated in a new window.
	--          The default angle of opening is given
	--          by the viewer.



    	Create ( VM : mutable Viewer ; V : PerspectiveView ) 
					returns mutable PerspectiveView ; 
	---Level: Public
	---Purpose: Creates one perspective view from another.
        --          The parameters of the original view are duplicated
        --          in the resulting view (Projection,Mapping,Context) .
        --          The view thus created must be activated in a new window.

        Copy ( me ) returns mutable PerspectiveView from V3d is static;
	---Level: Public
	
        --------------------------------------------------------
        ---Category: Methods to modify the status of the view
        --------------------------------------------------------

    	SetAngle ( me : mutable ; Angle : PlaneAngle ) 
	---Level: Public
	---Purpose: Modifies the angle of opening of the perspective in RADIANS.
	--	    The projection window is resized according to the
	--	    formula :
	--	    TAN(Angle/2) = Size/Length       
	--	    	Size expresses the smallest dimension of the window.
    	--	        Length expresses the focal length.
	raises BadValue from V3d
	---Purpose:  Warning! raises BadValue from V3d
	--	    if the opening angle is <= 0 or >= PI 
        is static;
	
    	Angle ( me ) returns PlaneAngle  is static; 
	---Level: Public
	---Purpose: Returns the value of the angle of opening.

    	SetPerspective ( me : mutable ; Angle : PlaneAngle; 
		                 UVRatio, ZNear, ZFar : Real ) 
	---Level: Public
	---Purpose: Modifies the viewing perspective volume by given
	--		angle of opening of the perspective in RADIANS,
	--      aspect ratio of window width to its height and 
	--      near and far clipping planes
	raises BadValue from V3d
	--	    if the opening angle is <= 0 or >= PI or
    --      the ZNear<0, ZFar<0 or ZNear>=Zfar.
        is static;
	
end PerspectiveView;
