-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class Torus   from gp   inherits Storable

        --- Purpose :
        --  Describes a torus.
        -- A torus is defined by its major and minor radii and
        -- positioned in space with a coordinate system (a gp_Ax3
        -- object) as follows:
        -- -   The origin of the coordinate system is the center of the torus;
        -- -   The surface is obtained by rotating a circle of radius
        --   equal to the minor radius of the torus about the "main
        --   Direction" of the coordinate system. This circle is
        --   located in the plane defined by the origin, the "X
        --   Direction" and the "main Direction" of the coordinate
        --   system. It is centered on the "X Axis" of this coordinate
        --   system, and located at a distance, from the origin of
        --   this coordinate system, equal to the major radius of the   torus;
        -- -   The "X Direction" and "Y Direction" define the
        --   reference plane of the torus.
        -- The coordinate system described above is the "local
        -- coordinate system" of the torus.
        -- Note: when a gp_Torus torus is converted into a
        -- Geom_ToroidalSurface torus, some implicit properties
        -- of its local coordinate system are used explicitly:
        -- -   its origin, "X Direction", "Y Direction" and "main
        --   Direction" are used directly to define the parametric
        --   directions on the torus and the origin of the parameters,
        -- -   its implicit orientation (right-handed or left-handed)
        --   gives the orientation (direct, indirect) to the
        --   Geom_ToroidalSurface torus.
        -- See Also
        -- gce_MakeTorus which provides functions for more
        -- complex torus constructions
        -- Geom_ToroidalSurface which provides additional
        -- functions for constructing tori and works, in particular,
        -- with the parametric equations of tori.




uses Array1OfReal from TColStd, 
     Ax1          from gp,
     Ax2          from gp,
     Ax3          from gp,
     Dir          from gp,
     Pnt          from gp,
     Trsf         from gp,
     Vec          from gp

raises ConstructionError from Standard,
       DimensionError    from Standard

is


  Create  returns Torus;
        ---C++: inline
        --- Purpose : creates an indefinite Torus.

  Create (A3 : Ax3; MajorRadius, MinorRadius : Real)   returns Torus
        ---C++: inline
        --- Purpose :
        -- a torus centered on the origin of coordinate system
        --   A3, with major radius MajorRadius and minor radius
        --   MinorRadius, and with the reference plane defined
        --   by the origin, the "X Direction" and the "Y Direction" of A3.
        --  Warnings :
        --  It is not forbidden to create a torus with
        --  MajorRadius = MinorRadius = 0.0 
        -- Raises ConstructionError if MinorRadius < 0.0 or if MajorRadius < 0.0
     raises ConstructionError;
    

  SetAxis (me : in out; A1 : Ax1)
        ---C++: inline
        --- Purpose : Modifies this torus, by redefining its local coordinate
        -- system so that:
        -- -   its origin and "main Direction" become those of the
        -- axis A1 (the "X Direction" and "Y Direction" are then recomputed).
        -- Raises ConstructionError if the direction of A1 is parallel to the "XDirection"
        --  of the coordinate system of the toroidal surface.
     raises ConstructionError
       
     is static;

  SetLocation (me : in out; Loc : Pnt)   is static;
        ---C++:inline
        --- Purpose : Changes the location of the torus.

  SetMajorRadius (me : in out; MajorRadius : Real)
        ---C++: inline
        --- Purpose : Assigns value to the major radius  of this torus. 
        -- Raises ConstructionError if MajorRadius - MinorRadius <= Resolution()
     raises ConstructionError
     
     is static;

  SetMinorRadius (me : in out; MinorRadius : Real)
        ---C++: inline
        --- Purpose : Assigns value to the  minor radius of this torus.
        -- Raises ConstructionError if MinorRadius < 0.0 or if
        --  MajorRadius - MinorRadius <= Resolution from gp.
     raises ConstructionError
       
     is static;

  SetPosition (me : in out; A3 : Ax3)   is static;
        ---C++: inline
        --- Purpose : Changes the local coordinate system of the surface.

  Area (me)  returns Real  is static;
        ---C++: inline
        --- Purpose : Computes the area of the torus.

  UReverse (me : in out)
        ---C++: inline
	---Purpose: Reverses the   U   parametrization of   the  torus
	--          reversing the YAxis.
  is static;

  VReverse (me : in out)
	---Purpose: Reverses the   V   parametrization of   the  torus
	--          reversing the ZAxis.
  is static;

  Direct (me) returns Boolean from Standard
        ---C++:inline
        ---Purpose: returns true if the Ax3, the local coordinate system of this torus, is right handed.
  is static;

  Axis (me)   returns Ax1  is static;
        ---C++:inline
        --- Purpose : returns the symmetry axis of the torus.
    	---C++: return const&

  Coefficients (me; Coef : out Array1OfReal from TColStd)
        --- Purpose :
        --  Computes the coefficients of the implicit equation of the surface
        --  in the absolute cartesian coordinate system :
        -- Coef(1) * X**4 + Coef(2) * Y**4 + Coef(3) * Z**4 +
        -- Coef(4) * X**3 * Y + Coef(5) * X**3 * Z + Coef(6) * Y**3 * X +
        -- Coef(7) * Y**3 * Z + Coef(8) * Z**3 * X + Coef(9) * Z**3 * Y +
        -- Coef(10) * X**2 * Y**2 + Coef(11) * X**2 * Z**2 +
        -- Coef(12) * Y**2 * Z**2 + Coef(13) * X**3 + Coef(14) * Y**3 +
        -- Coef(15) * Z**3 + Coef(16) * X**2 * Y + Coef(17) * X**2 * Z +
        -- Coef(18) * Y**2 * X + Coef(19) * Y**2 * Z + Coef(20) * Z**2 * X +
        -- Coef(21) * Z**2 * Y + Coef(22) * X**2 + Coef(23) * Y**2 +
        -- Coef(24) * Z**2 + Coef(25) * X * Y + Coef(26) * X * Z +
        -- Coef(27) * Y * Z + Coef(28) * X + Coef(29) * Y + Coef(30) *  Z + 
        -- Coef(31) = 0.0
        -- Raises DimensionError if the length of Coef is lower than 31.
     raises DimensionError
    
     is static;

  Location (me)  returns Pnt  is static;
        ---C++:inline
        --- Purpose : Returns the Torus's location.
    	---C++: return const&

  Position (me)  returns Ax3  is static;
        --- Purpose : Returns the local coordinates system of the torus.
        ---C++: inline
    	---C++: return const&

  MajorRadius (me) returns Real   is static;
        --- Purpose : returns the major radius of the torus.
        ---C++: inline

  MinorRadius (me) returns Real   is static;
        --- Purpose : returns the minor radius of the torus.
        ---C++: inline

  Volume (me)  returns Real  is static;
        --- Purpose : Computes the volume of the torus.
        ---C++: inline

  XAxis (me)  returns Ax1   is static;
        ---C++:inline
        --- Purpose : returns the axis X of the torus.

  YAxis (me)  returns Ax1  is static;
        ---C++:inline
        --- Purpose : returns the axis Y of the torus.

       
  Mirror (me : in out; P : Pnt)   
       is static;

  Mirrored (me; P : Pnt)  returns Torus  is static;
 --- Purpose :
        --  Performs the symmetrical transformation of a torus 
        --  with respect to the point P which is the center of the 
        --  symmetry.

                    
   
  Mirror (me : in out; A1 : Ax1)    
       is static;

  Mirrored (me; A1 : Ax1)   returns Torus  is static;
        --- Purpose :
        --  Performs the symmetrical transformation of a torus with
        --  respect to an axis placement which is the axis of the
        --  symmetry.



     
  Mirror (me : in out; A2 : Ax2)    
        is static;

  Mirrored (me; A2 : Ax2)    returns Torus  is static;
        --- Purpose :
        --  Performs the symmetrical transformation of a torus with respect 
        --  to a plane. The axis placement A2 locates the plane of the
        --  of the symmetry : (Location, XDirection, YDirection).


  Rotate (me : in out; A1 : Ax1; Ang : Real)
        ---C++:inline
        is static;

  Rotated (me; A1 : Ax1; Ang : Real) returns Torus  is static;
        ---C++:inline

        --- Purpose :
        --  Rotates a torus. A1 is the axis of the rotation.
        --  Ang is the angular value of the rotation in radians.



  Scale (me : in out; P : Pnt; S : Real)         is static;
        ---C++:inline

  Scaled (me; P : Pnt; S : Real)  returns Torus  is static;
        ---C++:inline


        --- Purpose : 
        --  Scales a torus. S is the scaling value.
        --  The absolute value of S is used to scale the torus



  Transform (me : in out; T : Trsf)              is static;
        ---C++:inline

  Transformed (me; T : Trsf)     returns Torus   is static;
        ---C++:inline

        --- Purpose :
        --  Transforms a torus with the transformation T from class Trsf.

      
       

  Translate (me : in out; V : Vec) 
        ---C++:inline
        is static;

  Translated (me; V : Vec)  returns Torus  is static;
        ---C++:inline
        --- Purpose :
        --  Translates a torus in the direction of the vector V.
        --  The magnitude of the translation is the vector's magnitude.

     
  Translate (me : in out; P1, P2 : Pnt)         is static;   
        ---C++:inline

  Translated (me; P1, P2 : Pnt)  returns Torus  is static;
        ---C++:inline
        --- Purpose :
        --  Translates a torus from the point P1 to the point P2.



fields

  pos         : Ax3;
  majorRadius : Real;
  minorRadius : Real;

end;


