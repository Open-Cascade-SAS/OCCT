-- Created on: 1998-07-22
-- Created by: Christian CAILLET
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Vars  from XSControl    inherits TShared  from MMgt

    ---Purpose : Defines a receptacle for externally defined variables, each
    --           one has a name
    --           
    --           I.E. a WorkSession for XSTEP is generally used inside a
    --           context, which brings variables, especially shapes and
    --           geometries. For instance DRAW or an application engine
    --           
    --           This class provides a common form for this. It also provides
    --           a default implementation (locally recorded variables in a
    --           dictionary), but which is aimed to be redefined

uses CString, Transient, DictionaryOfTransient,
     Pnt from gp, Pnt2d from gp,
     Geometry from Geom, Curve from Geom, Curve from Geom2d, Surface from Geom,
     Shape from TopoDS

is

    Create returns Vars;

    Set (me : mutable; name : CString; val : Transient)  is virtual;

    Get (me; name : in out CString) returns Transient  is virtual;


    GetGeom (me; name : in out CString) returns Geometry  is virtual;

    GetCurve2d (me; name : in out CString) returns Curve from Geom2d  is virtual;

    GetCurve   (me; name : in out CString) returns Curve from Geom  is virtual;

    GetSurface (me; name : in out CString) returns Surface from Geom  is virtual;

    SetPoint   (me : mutable; name : CString; val : Pnt   from gp)  is virtual;

    SetPoint2d (me : mutable; name : CString; val : Pnt2d from gp)  is virtual;

    GetPoint   (me; name : in out CString; pnt : out Pnt   from gp) returns Boolean  is virtual;

    GetPoint2d (me; name : in out CString; pnt : out Pnt2d from gp) returns Boolean  is virtual;


    SetShape   (me : mutable; name : CString; val : Shape from TopoDS)  is virtual;

    GetShape   (me; name : in out CString) returns Shape from TopoDS  is virtual;

fields

    thevars : DictionaryOfTransient;

end Vars;
