-- Created on: 1993-03-10
-- Created by: JCV
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



deferred class Point from Geom inherits Geometry from Geom



    	---Purpose : The abstract class Point describes the common
    	-- behavior of geometric points in 3D space.
    	-- The Geom package also provides the concrete class
    	-- Geom_CartesianPoint.

uses Pnt from gp

is


  Coord (me; X, Y, Z : out Real) 
        ---Purpose : returns the Coordinates of <me>.
     is deferred;


  Pnt (me)  returns Pnt
        ---Purpose : returns a non transient copy of <me>
     is deferred;


  X (me)  returns Real
        ---Purpose : returns the X coordinate of <me>.
     is deferred;


  Y (me)  returns Real
        ---Purpose : returns  the Y coordinate of <me>.
     is deferred;


  Z (me)   returns Real
        ---Purpose : returns the Z coordinate of <me>.
     is deferred;


  Distance (me; Other : Point)  returns Real;
        ---Purpose : Computes the distance between <me> and <Other>.

  
  SquareDistance (me; Other : Point)  returns Real;
        ---Purpose : Computes the square distance between <me> and <Other>.

end;

