-- Created on: 2000-07-10
-- Created by: Vincent DELOS
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class AncestorsAndSuccessors from BooleanOperations 

	---Purpose:   provides all the ancestors   and successors of a
	--          given  shape. Exemple : for  an edge the ancestors
	--          are the wires that hold it  and the successors are
	--          its vertices.

uses
    Orientation from TopAbs,
    SequenceOfInteger from TColStd,
    AncestorsSeqAndSuccessorsSeq from BooleanOperations
    
is

    Create returns AncestorsAndSuccessors from BooleanOperations;
      
    Create (AncSuccessors: AncestorsSeqAndSuccessorsSeq; shift: Integer) returns AncestorsAndSuccessors from BooleanOperations;
    ---Purpose: allocates space and fills it with the data of AncSuccessors.
    
    Destroy(me:in out);
    ---C++: alias ~
	
    
    Dump (me);
    ---Purpose: to display the fields.

    
    --------------------
    -- INLINE METHODS --
    --------------------

    GetAncestor (me; AncestorIndex: Integer) returns Integer;
    ---C++: inline    
    SetAncestor (me:in out; AncestorIndex,AncestorNumber: Integer);
    ---C++: inline
    GetAncestors(me; theArrayOfAncestors:out Address;AncestorsNumber:out Integer);
    ---C++: inline    
    
    GetSuccessor (me; SuccessorIndex: Integer) returns Integer;
    ---C++: inline    
    SetSuccessor (me:in out; SuccessorIndex,SuccessorNumber: Integer);
    ---C++: inline
    GetSuccessors(me; theArrayOfSuccessors:out Address; SuccessorsNumber:out Integer);
    ---C++: inline    

    GetOrientation (me; OrientationIndex: Integer) returns Orientation;
    ---C++: inline    
    SetOrientation (me:in out; OrientationIndex: Integer; anOrientation: Orientation from TopAbs);
    ---C++: inline
    GetOrientations(me; theArrayOfOrientations:out Address;OrientationsNumber:out Integer);
    ---C++: inline    

    NumberOfAncestors  (me) returns Integer;
    ---C++: inline
    NumberOfSuccessors (me) returns Integer;
    ---C++: inline


fields

myAncestors: Address;
---Purpose: the array containing all the ancestors of our given shape.

mySuccessors: Address;
---Purpose: the array containing all the successors.

myOrientations: Address;
---Purpose: the array containing all the orientation of the successors.

myAncestorsSize : Integer;
---Purpose: the number of ancestors.

mySuccessorsSize: Integer;
---Purpose: the number of successors.

end AncestorsAndSuccessors;
