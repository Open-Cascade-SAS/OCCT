-- Created on: 1999-04-06
-- Created by: Fabrice SERVANT
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

--  modified by Edward AGAPOV (eap) Thu Feb 14 2002 (occ139)
--  Add Prepend(), replace array with sequence

class SectionLine from IntPolyh

uses
    
    SeqOfStartPoints from IntPolyh,
    StartPoint from IntPolyh


is


    Create;
    
    Create(nn : Integer from Standard) ; 
    
    Init(me: in out; nn: Integer from Standard) 
    is static;

    Value(me; nn: Integer from Standard)
    	---C++: alias operator [] 
    	---C++: return const &
    returns StartPoint from IntPolyh    
    is static;
    
    ChangeValue(me: in out;  nn: Integer from Standard)
    	---C++: alias operator [] 
    	---C++: return &
    returns StartPoint from IntPolyh    
    is static;
    
    Copy(me: in out; Other : SectionLine from IntPolyh)
    	---C++: alias operator =
    	---C++: return &
    returns SectionLine from IntPolyh
    is static;
    
    GetN(me)
    returns Integer from Standard
    is static;
    
    NbStartPoints(me)
    returns Integer from Standard
    is static;
    
    IncrementNbStartPoints(me: in out)
    is static;
    
    Destroy(me: in out)
    	---C++: alias ~
    is static;
    
    Dump(me) 
    is static;
    
    Prepend(me:in out; SP: StartPoint from IntPolyh)
    is static;
     	
fields

--    n,nbstartpoints : Integer from Standard;
--    ptr :Address from Standard;
    mySeqOfSPoints : SeqOfStartPoints from IntPolyh;
    
end SectionLine from IntPolyh;
