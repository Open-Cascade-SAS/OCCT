-- File:	RWStepDimTol_RWFlatnessTolerance.cdl
-- Created:	Wed Jun  4 13:34:34 2003 
-- Author:	Galina KULIKOVA
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWFlatnessTolerance from RWStepDimTol

    ---Purpose: Read & Write tool for FlatnessTolerance

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    FlatnessTolerance from StepDimTol

is
    Create returns RWFlatnessTolerance from RWStepDimTol;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : FlatnessTolerance from StepDimTol);
	---Purpose: Reads FlatnessTolerance

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: FlatnessTolerance from StepDimTol);
	---Purpose: Writes FlatnessTolerance

    Share (me; ent : FlatnessTolerance from StepDimTol;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWFlatnessTolerance;
