-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class BoxDomain from StepShape 

inherits TShared from MMgt

uses

	CartesianPoint from StepGeom, 
	Real from Standard
is

	Create returns mutable BoxDomain;
	---Purpose: Returns a BoxDomain

	Init (me : mutable;
	      aCorner : mutable CartesianPoint from StepGeom;
	      aXlength : Real from Standard;
	      aYlength : Real from Standard;
	      aZlength : Real from Standard) is virtual;

	-- Specific Methods for Field Data Access --

	SetCorner(me : mutable; aCorner : mutable CartesianPoint);
	Corner (me) returns mutable CartesianPoint;
	SetXlength(me : mutable; aXlength : Real);
	Xlength (me) returns Real;
	SetYlength(me : mutable; aYlength : Real);
	Ylength (me) returns Real;
	SetZlength(me : mutable; aZlength : Real);
	Zlength (me) returns Real;

fields

	corner : CartesianPoint from StepGeom;
	xlength : Real from Standard;
	ylength : Real from Standard;
	zlength : Real from Standard;

end BoxDomain;
