-- Created on: 1992-08-26
-- Created by: Jean Louis FRENKEL
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package StdPrs
    	---Purpose: The StdPrs package provides standard display tools
	-- for specific geometries and topologies whereas
	-- Prs3d provides those for generic objects. Among
	-- these classes are definitions of the display of the
	-- specific geometry or topology in various display
	-- modes such as wireframe, shading or hidden line removal mode.
    	       
uses
  Prs3d,
	Geom,
	Geom2d,
	Adaptor3d,
	Adaptor2d,
  GeomAdaptor,
	Geom2dAdaptor,
  BRepAdaptor,
	TopTools,
	TopoDS,
	TopExp,
  TopAbs,
	BRepTools,
	Bnd,
  TColStd,
  HLRAlgo,
  HLRBRep,
  Quantity,
	BRepMesh,
	gp,
	TColgp,
	Poly,
	TopLoc, 
	Graphic3d

is
   class ToolPoint;
   class ToolVertex;
   class ToolRFace;
   class HLRToolShape;
   class ToolShadedShape;
   class ShadedShape;
    
   class PoleCurve;
	---Purpose: computes the presentation of curves by drawing
	--          a broken line linking the poles of the curve.

   class Plane;
   	---Purpose: computes the presentation of a infinite plane.

   class WFPoleSurface;
   	---Purpose: computes the presentation of surfaces by drawing a
	--          double network of lines linking the poles of the surface
	--          in the two parametric direction.
	

   class DeflectionCurve;		      
	---Purpose: computes the presentation of objects to be
	--          seen as curves. The computation will be made
	--          according to a maximal chordial deviation.
	          
	---Category: Wireframe algorithms
   
   class WFDeflectionSurface;
	---Purpose: computes the wireframe presentation of surfaces 
	--          by displaying a given number of U and/or V isoparametric
	---         curves. The isoparametric curves are drawn with respect
	--          to a given maximal chordial deviation.

   class ShadedSurface;
   	---Purpose: computes the shading presentation of surfaces.

   -----------------------------------------------
   --- deflection drawing classes :
   -----------------------------------------------

   class WFDeflectionRestrictedFace;
	  ---Purpose: computes the wireframe presentation of faces with
	--          restrictions by displaying a given number of U and/or
	--          V isoparametric curves. The isoparametric curves are
	--          drawn with respect to a maximal chordial deviation.
	--          The presentation includes the restriction curves.
		      
   class Curve;
   	---Purpose: computes the presentation of objects to be
	--          seen as curves. The computation will be made
	--          whith a constant number of points.


   class WFSurface;
   	---Purpose: computes the wireframe presentation of surfaces 
	--          by displaying a given number of U and/or V isoparametric
	---         curves. The isoparametric curves are drawn with respect
	--          to a given number of points.
			
   
   ---Category: Hidden lines removal algorithms.
   
   class HLRPolyShape; 
    ---Purpose: computes the presentation of objects with
	--          removal of their hidden lines for a specific
	--          projector. The polygonal algorithm is used.
  
   imported HLRShape;
   ---Purpose: computes the presentation of objects with
	--          removal of their hidden lines for a specific
	--          projector. The exact algorithm is used.
     
   imported NListOfSequenceOfPnt from Prs3d; 
   imported NListIteratorOfListOfSequenceOfPnt from Prs3d;
   
   imported WFShape;
   imported WFDeflectionShape;
   ---Purpose: computes the wireframe presentation of surfaces 
	--          by displaying planar sections.
   imported Vertex;
   imported Point;
   ---Purpose: computes the presentation of objects to be
	--          seen as points.
   imported WFRestrictedFace;
   ---Purpose:  Computes the wireframe presentation of faces with
  --           restrictions by displaying a given number of U and/or
  --           V isoparametric curves. The isoparametric curves are
  --           drawn with a fixed number of points.
  --           The presentation includes the restriction curves.
			
end StdPrs;



