-- Created on: 1996-02-01
-- Created by: Philippe MANGIN
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



private class EnergyOfBatten from FairCurve inherits Energy from FairCurve

	---Purpose: Energy Criterium to minimize in Batten.
	---Category: Private use

uses BattenLaw from FairCurve,  
     DistributionOfTension from FairCurve, 
     DistributionOfSagging from FairCurve,
     AnalysisCode from FairCurve,
     Vector  from  math,
     Matrix  from math,
     HArray1OfPnt2d from TColgp,
     Array1OfXY  from TColgp,
     Pnt2d from gp,
     HArray1OfReal from TColStd


is
    Create( BSplOrder     : Integer;
            FlatKnots     : HArray1OfReal;
	    Poles         : HArray1OfPnt2d;
    	    ContrOrder1   : Integer;
	    ContrOrder2   : Integer;
	    Law           : BattenLaw;
	    LengthSliding : Real;
	    FreeSliding   : Boolean = Standard_True;
            Angle1        : Real = 0;
            Angle2        : Real = 0 ) returns  EnergyOfBatten;
	    ---Purpose: Angles corresspond to the Ox axis

    
    LengthSliding(me)
    ---Purpose: return  the  lengthSliding = P1P2 + Sliding
    ---C++: inline
    returns  Real;
 
     
    Status(me) 
    ---Purpose: return  the status 
    ---C++: inline
    returns  AnalysisCode;
    
    
    ComputePoles(me: in out; X: Vector)
    ---Purpose: compute  the  poles wich correspond with the variable X
    is redefined protected; 
    
    Variable(me; X: out Vector)
    ---Purpose: compute the variables <X> wich correspond with the field <MyPoles>
    returns Boolean
    is redefined;  
	
    Compute(me:in out; DerivativeOrder : Integer; Result : out Vector)
        ---Purpose: compute the energy in intermediat format
    returns Boolean 
    is redefined protected;
    
fields
    MyLengthSliding : Real;
    OriginalSliding : Real;
    MyFreeSliding   : Boolean;
    MyBattenLaw     : BattenLaw;
    MyTension       : DistributionOfTension;
    MySagging       : DistributionOfSagging;
    MyStatus        : AnalysisCode;
    
end EnergyOfBatten;
