-- Created on: 1999-11-11
-- Created by: Vladislav ROMASHKO
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class BooleanOperation from QANewBRepNaming inherits TopNaming from QANewBRepNaming

    ---Purpose: To load the BooleanOperation results
	
uses 
 
--modified by NIZNHY-PKV Wed Jun 19 09:06:12 2002  f  
    BooleanOperation from BRepAlgo,
    --BooleanOperation from BRepAlgoAPI, 
--modified by NIZNHY-PKV Wed Jun 19 09:06:16 2002  t    
    Shape            from TopoDS,
    Label            from TDF,
    ListOfShape      from TopTools

is
 
    Create returns BooleanOperation from QANewBRepNaming;

    Create(ResultLabel : Label from TDF) 
    returns BooleanOperation from QANewBRepNaming;

    Init(me : in out; ResultLabel :  Label from TDF);
	 
--modified by NIZNHY-PKV Wed Jun 19 09:06:46 2002  f	
    Load (me; mkBoolOp : in out BooleanOperation from BRepAlgo);
--    Load (me; mkBoolOp : in out BooleanOperation from BRepAlgoAPI); 
--modified by NIZNHY-PKV Wed Jun 19 09:06:53 2002  t 

    ---Purpose : Load the boolean operation.
    --           Makes a new part attached to the ResultLabel.

    FirstModified (me)
    ---Purpose: Returns the label of the modified faces
    --          of the first shape (S1).
    returns Label from TDF;  
    
    FirstDeleted (me)
    ---Purpose: Returns the label of the deleted faces
    --          of the first shape (S1).
    returns Label from TDF; 

    SecondModified (me)
    ---Purpose: Returns the label of the modified faces
    --          of the second shape (S2).
    returns Label from TDF;  
    
    SecondDeleted (me)
    ---Purpose: Returns the label of the deleted faces
    --          of the second shape (S2).
    returns Label from TDF; 
          
    Intersections (me)
    ---Purpose: Returns the label of intersections
    returns Label from TDF; 
     
end BooleanOperation;
