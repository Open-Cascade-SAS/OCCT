-- Created on: 1997-04-11
-- Created by: VAUTHIER Jean-Claude
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class NamedShape from PNaming inherits Attribute from PDF

	---Purpose: This is the persistent attribute of the
	--          topological naming.

uses

    HArray1OfShape1 from PTopoDS,
    HArray1OfInteger from PColStd


is


    Create returns mutable NamedShape from PNaming;
	---Purpose: Creates a mutable NamedShape from PNaming.

    
    NbShapes(me) returns Integer;
	---Purpose: Returns the number of shapes.


    OldShapes(me : mutable; theShapes : HArray1OfShape1 from PTopoDS);
	---Purpose: Sets the field <myOldShapes>.
    
    OldShapes(me) returns HArray1OfShape1 from PTopoDS;
	---Purpose: Returns the field <myOldShapes>.
    

    NewShapes(me : mutable; theShapes : HArray1OfShape1 from PTopoDS);
	---Purpose: Sets the field <myNewShapes>.
    
    NewShapes(me) returns HArray1OfShape1 from PTopoDS;
	---Purpose: Returns the field <myNewShapes>.
    

    ShapeStatus(me : mutable; theShapeStatus : Integer from Standard);
	---Purpose: Sets the field <myShapeStatus>.
    
    ShapeStatus(me) returns Integer from Standard;
	---Purpose: Returns the field <myShapeStatus>.
    
    Version (me : mutable; theVersion : Integer from Standard);
    	---Purpose: Sets the field <myVersion>.
    
    Version (me) returns Integer from Standard;
        ---Purpose: Returns the field <myVersion>.
	    
fields

    myOldShapes    : HArray1OfShape1 from PTopoDS;
    myNewShapes    : HArray1OfShape1 from PTopoDS;
    myShapeStatus  : Integer         from Standard;
    myVersion      : Integer         from Standard;

end NamedShape;
