-- Created on: 1998-07-14
-- Created by: data exchange team
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package ShapeConstruct 

	---Purpose: This package provides new algorithms for constructing
-- new geometrical objects and topological shapes. It
-- complements and extends algorithms available in Open
-- CASCADE topological and geometrical toolkist.
-- The functionality provided by this package are the
-- following: 
  --    projecting curves on surface, 
--      adjusting curve to have given start and end points. P
uses
    gp,
    Geom,
    GeomAbs,
    Geom2d,
    TColgp,
    TColStd,
    ShapeExtend,
    ShapeAnalysis,
    Convert,
    BRepBuilderAPI,
    TopoDS,
    TopAbs,
    TopTools

is

    class Curve;

    class ProjectCurveOnSurface;

    ---WARNING: The following two classes are just a copy of those from GEOMLITE
    --          They must be removed as soon as bug in them is fixed	

    class CompBezierCurvesToBSplineCurve;

    class CompBezierCurves2dToBSplineCurve2d;

    class MakeTriangulation;
    	---Purpose: Tool for wire triangulation

    ConvertCurveToBSpline(C3D        : Curve from Geom;
    	    	    	  First      : Real;
			  Last       : Real;
    	    	    	  Tol3d      : Real; -- this and following parameters are used only if approximator have to be used.
			  Continuity : Shape from GeomAbs; 
    	    	    	  MaxSegments: Integer;
			  MaxDegree  : Integer)
    returns BSplineCurve from Geom;
    
    ConvertCurveToBSpline(C2D        : Curve from Geom2d;
    	    	    	  First      : Real;
			  Last       : Real;
    	    	    	  Tol2d      : Real; -- this and following parameters are used only if approximator have to be used.
			  Continuity : Shape from GeomAbs; 
    	    	    	  MaxSegments: Integer;
			  MaxDegree  : Integer)
    returns BSplineCurve from Geom2d;
    
    ConvertSurfaceToBSpline(surf       : Surface from Geom;
    			   UF,UL,VF,VL: Real;
			   Tol3d      : Real; -- this and following parameters are used only if approximator have to be used.
			   Continuity : Shape from GeomAbs; 
    	    	    	   MaxSegments: Integer;
			   MaxDegree  : Integer)
    returns BSplineSurface from Geom;
        
    JoinPCurves(theEdges : HSequenceOfShape from TopTools;
    	    	theFace  : Face from TopoDS;
    	    	theEdge : in out Edge from TopoDS)
    returns Boolean from Standard;
    	---Purpose: join pcurves of the <theEdge> on the <theFace>
	--    	    try to use pcurves from originas edges <theEdges>
    	--          Returns false if cannot join pcurves
	
    JoinCurves(c3d1,ac3d2 : Curve from Geom; 
    	    	Orient1, Orient2 : Orientation from TopAbs;
		first1,last1,first2,last2 : in out Real;
		c3dOut : out Curve from Geom;
		isRev1,isRev2 : out Boolean) returns Boolean;
		
    --- Purpose:Method for joininig curves 3D. 
    --          Parameters : c3d1,ac3d2 - initial curves
    --	                     Orient1, Orient2 - initial edges orientations.
    --                       first1,last1,first2,last2 - parameters for trimming curves 
    --	    	             (re-calculate with account of orientation edges)
    --                       c3dOut - result curve
    --                       isRev1,isRev2 - out parameters indicative on possible errors.
    --          Return value : True - if curves were joined successfully,
    --                               else - False.
    
    JoinCurves(c2d1,ac2d2 : Curve from Geom2d; 
    	    	Orient1, Orient2 : Orientation from TopAbs;
		first1,last1,first2,last2 : in out Real;
		c2dOut : out Curve from Geom2d;
		isRev1,isRev2 : out Boolean;
                isError : Boolean = Standard_False) returns Boolean;
		
    --- Purpose:Method for joininig curves 3D. 
    --          Parameters : c3d1,ac3d2 - initial curves
    --	                     Orient1, Orient2 - initial edges orientations.
    --                       first1,last1,first2,last2 - parameters for trimming curves 
    --	    	             (re-calculate with account of orientation edges)
    --                       c3dOut - result curve
    --                       isRev1,isRev2 - out parameters indicative on possible errors.
    --                       isError - input parameter indicative possible errors due to that one from edges have one vertex
    --         Return value : True - if curves were joined successfully,
    --                               else - False.
end ShapeConstruct;
