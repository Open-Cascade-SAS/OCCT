-- File:	BRepGProp_Face.cdl
-- Created:	Wed Apr 14 18:04:46 1993
-- Author:	Isabelle GRIGNON
--		<isg@sdsun2>
---Copyright:	 Matra Datavision 1993

class Face  from BRepGProp  

uses Pnt2d         from gp,
     Vec2d         from gp,
     Pnt           from gp,
     Vec           from gp,
     Edge          from TopoDS,
     Face          from TopoDS,
     Surface       from BRepAdaptor,
     Curve         from Geom2dAdaptor,
     Array1OfReal  from TColStd, 
     HArray1OfReal from TColStd, 
     IsoType       from GeomAbs
     
is 

  Create (IsUseSpan: Boolean from Standard = Standard_False) 
        ---Purpose: Constructor. Initializes the object with a flag IsUseSpan 
        --          that says if it is necessary to define spans on a face. 
        --          This option has an effect only for BSpline faces. Spans 
        --          are returned by the methods GetUKnots and GetTKnots.
	---C++: inline
  returns Face from BRepGProp;

  Create(F        : Face    from TopoDS; 
         IsUseSpan: Boolean from Standard = Standard_False) 
        ---Purpose: Constructor. Initializes the object with the face and the 
        --          flag IsUseSpan that says if it is necessary to define 
        --          spans on a face. This option has an effect only for 
        --          BSpline faces. Spans are returned by the methods GetUKnots 
        --          and GetTKnots.
	---C++: inline
  returns Face from BRepGProp;

  Load(me : in out; F : Face from TopoDS) 
  is static;

  VIntegrationOrder (me) returns Integer
  is static;
 
  NaturalRestriction(me) returns Boolean
    	---Purpose: Returns Standard_True if the face is not trimmed.
	---C++: inline
  is static;

  Value2d (me; U :Real) returns Pnt2d from gp 
        ---Purpose: Returns the value of the boundary curve of the face.
	---C++: inline
  is static;
  
  SIntOrder (me; Eps :Real) returns Integer
  is static;
  SVIntSubs (me) returns Integer
  is static;
  SUIntSubs (me) returns Integer
  is static;
  UKnots(me; Knots : out Array1OfReal from TColStd)
  is static;
  VKnots(me; Knots : out Array1OfReal from TColStd)
  is static;
  LIntOrder (me; Eps :Real) returns Integer
  is static;
  LIntSubs (me) returns Integer
  is static;
  LKnots(me; Knots : out Array1OfReal from TColStd)
  is static;
 
  --
  --   Methods required by GProp
  --   
    
  UIntegrationOrder (me) returns Integer
        ---Purpose: Returns the number of points required to do the 
        --          integration in the U parametric direction with 
        --          a good accuracy.
  is static;

  Bounds(me; U1,U2,V1,V2 : out Real)
        ---Purpose: Returns the parametric bounds of the Face.
  is static;
  
  Normal (me;  U, V : Real; P : out Pnt; VNor: out Vec)
	---Purpose: Computes the point of parameter U, V on the Face <S> and 
	--          the normal to the face at this point.
  is static;
 
  Load(me : in out; E : Edge from TopoDS) 
        ---Purpose: Loading the boundary arc.
  is static;

  FirstParameter (me) returns Real 
        ---Purpose: Returns the parametric value of the start point of
        --          the current arc of curve. 
	---C++: inline
  is static;

  LastParameter (me) returns Real 
        ---Purpose: Returns the parametric value of the end point of
        --          the current arc of curve. 
	---C++: inline
  is static;

  IntegrationOrder (me) returns Integer
        ---Purpose: Returns the number of points required to do the 
        --          integration along the parameter of curve.
  is static;

  D12d (me; U : Real ;P  : out Pnt2d from gp ;
                      V1 : out Vec2d from gp)
    	---Purpose: Returns the point of parameter U and the first derivative 
    	--          at this point of a boundary curve.
	---C++: inline
  is static;

-- Modified by skv - Fri Dec  9 16:44:00 2005 Begin 
  Load(me : in out; IsFirstParam: Boolean from Standard; 
                    theIsoType  : IsoType from GeomAbs);
        ---Purpose: Loading the boundary arc. This arc is either a top, bottom, 
        --          left or right bound of a UV rectangle in which the 
        --          parameters of surface are defined. 
	--          If IsFirstParam is equal to Standard_True, the face is 
        --          initialized by either left of bottom bound. Otherwise it is 
        --          initialized by the top or right one. 
	--          If theIsoType is equal to GeomAbs_IsoU, the face is 
        --          initialized with either left or right bound. Otherwise - 
        --          with either top or bottom one.

  GetUKnots(me; theUMin  :        Real          from Standard; 
                theUMax  :        Real          from Standard; 
		theUKnots: in out HArray1OfReal from TColStd);
	---Purpose: Returns an array of U knots of the face. The first and last 
        --          elements of the array will be theUMin and theUMax. The 
        --          middle elements will be the U Knots of the face greater 
        --          then theUMin and lower then theUMax in increasing order. 
	--          If the face is not a BSpline, the array initialized with 
        --          theUMin and theUMax only.

  GetTKnots(me; theTMin  :        Real          from Standard; 
                theTMax  :        Real          from Standard; 
		theTKnots: in out HArray1OfReal from TColStd);
	---Purpose: Returns an array of combination of T knots of the arc and 
        --          V knots of the face. The first and last elements of the 
        --          array will be theTMin and theTMax. The middle elements will 
        --          be the Knots of the arc and the values of parameters of 
        --          arc on which the value points have V coordinates close to V 
        --          knots of face. All the parameter will be greater then 
        --          theTMin and lower then theTMax in increasing order.
	--          If the face is not a BSpline, the array initialized with 
        --          theTMin and theTMax only.

-- Modified by skv - Fri Dec  9 16:44:00 2005 End

fields

    mySurface  : Surface from BRepAdaptor;
    myCurve    : Curve   from Geom2dAdaptor;
    mySReverse : Boolean from Standard;
    myIsUseSpan: Boolean from Standard;

end Face;
