-- Created on: 1993-03-26
-- Created by: Laurent BUCHARD
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


generic class MultiLineTool from ApproxInt (TheMultiLine   as any;
    	    	    	                    TheMultiMPoint as any)


uses 
      Status           from Approx,
      Array1OfPnt      from TColgp,
      Array1OfPnt2d    from TColgp,
      Array1OfVec      from TColgp,
      Array1OfVec2d    from TColgp
    
is
    
    
    FirstPoint(myclass; ML: TheMultiLine) returns Integer;
    	---C++:inline
    	---Purpose: Returns the number of multipoints of the TheMultiLine.

    LastPoint(myclass; ML: TheMultiLine) returns Integer;
    	---C++:inline
    	---Purpose: Returns the number of multipoints of the TheMultiLine.

    NbP2d(myclass; ML: TheMultiLine) returns Integer;
    	---C++:inline
    	---Purpose: Returns the number of 2d points of a TheMultiLine.


    NbP3d(myclass; ML: TheMultiLine) returns Integer; 
    	---C++:inline
   	---Purpose: Returns the number of 3d points of a TheMultiLine.


    Value(myclass; ML:  TheMultiLine; MPointIndex: Integer; tabPt: out Array1OfPnt);
    	---C++:inline
    	---Purpose: returns the 3d points of the multipoint <MPointIndex>
    	--          when only 3d points exist.


    Value(myclass; ML:  TheMultiLine; MPointIndex: Integer; 
          tabPt2d: out Array1OfPnt2d from TColgp);
    	---C++:inline
    	---Purpose: returns the 2d points of the multipoint <MPointIndex>
    	--          when only 2d points exist.


    Value(myclass; ML:  TheMultiLine; MPointIndex: Integer; 
          tabPt: out Array1OfPnt from TColgp; tabPt2d: out Array1OfPnt2d);
    	---C++:inline
    	---Purpose: returns the 3d and 2d points of the multipoint 
    	--          <MPointIndex>.

    Tangency(myclass; ML:  TheMultiLine; MPointIndex: Integer; tabV: out Array1OfVec from TColgp)
    returns Boolean;
    	---C++:inline
    	---Purpose: returns the 3d points of the multipoint <MPointIndex>
    	--          when only 3d points exist.


    Tangency(myclass; ML:  TheMultiLine; MPointIndex: Integer; 
          tabV2d: out Array1OfVec2d from TColgp)
    returns Boolean;
    	---C++:inline
    	---Purpose: returns the 2d tangency points of the multipoint 
    	--          <MPointIndex> only when 2d points exist.


    Tangency(myclass; ML:  TheMultiLine; MPointIndex: Integer; 
             tabV: out Array1OfVec from TColgp; tabV2d: out Array1OfVec2d from TColgp)
    returns Boolean;
    	---C++:inline
    	---Purpose: returns the 3d and 2d points of the multipoint 
    	--          <MPointIndex>.


--- methods not used but necessary


    Curvature(myclass; ML:  TheMultiLine; MPointIndex: Integer; 
             tabV: out Array1OfVec from TColgp)
    returns Boolean;
    	---C++:inline
    	---Purpose: returns the 3d curvature of the multipoint <MPointIndex>
    	--          when only 3d points exist.


    Curvature(myclass; ML:  TheMultiLine; MPointIndex: Integer; 
          tabV2d: out Array1OfVec2d from TColgp)
    returns Boolean;
    	---C++:inline
    	---Purpose: returns the 2d curvature points of the multipoint 
    	--          <MPointIndex> only when 2d points exist.


    Curvature(myclass; ML:  TheMultiLine; MPointIndex: Integer; 
             tabV: out Array1OfVec from TColgp; 
             tabV2d: out Array1OfVec2d from TColgp)
    returns Boolean;
    	---C++:inline
    	---Purpose: returns the 3d and 2d curvature of the multipoint 
    	--          <MPointIndex>.

    
     
    MakeMLBetween(myclass; ML:  TheMultiLine; I1, I2: Integer;
                  NbPMin: Integer) 
    returns TheMultiLine;
    	---C++:inline
    	---Purpose: Is called if WhatStatus returned "PointsAdded".
   
    WhatStatus(myclass; ML:  TheMultiLine; I1, I2: Integer) 
    	---C++:inline
    returns Status from Approx;
    
end MultiLineTool;    

