-- Created on: 1992-06-22
-- Created by: Gilles DEBARBOUILLE
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Quantity from Units 

inherits

    TShared from MMgt 


	---Purpose: This  class stores  in its  field all the possible
	--          units of all the unit systems for a given physical
	--          quantity. Each unit's  value  is  expressed in the
	--          S.I. unit system.

uses

    UnitsSequence from Units,
    Dimensions    from Units,
    HAsciiString  from TCollection,
    AsciiString   from TCollection

is

    Create(aname          : CString ;
           adimensions    : Dimensions    from Units ;
           aunitssequence : UnitsSequence from Units)
    
    ---Level: Internal 
    
    ---C++: inline
    
    ---Purpose: Creates  a new Quantity  object with <aname> which  is
    --          the name of the physical quantity, <adimensions> which
    --          is the physical dimensions, and <aunitssequence> which
    --          describes all the units known for this quantity.
    
    returns Quantity from Units;
    
    Name(me) returns AsciiString from TCollection
    
    ---Level: Internal 
    
    ---C++: inline
    
    ---Purpose: Returns in a AsciiString from TCollection the name of the quantity.
    
    is static;
    
    Dimensions(me) returns any Dimensions from Units
    
    ---Level: Internal 
    
    ---C++: inline
    
    ---Purpose: Returns the physical dimensions of the quantity.
    
    is static;
    
    Sequence(me) returns any UnitsSequence from Units
    
    ---Level: Internal 
    
    ---C++: inline
    
    ---Purpose: Returns <theunitssequence>, which  is the  sequence of
    --          all the units stored for this physical quantity.
    
    is static;
    
    IsEqual(me ; astring : CString) returns Boolean
    
    ---Level: Internal 
    
--    ---C++: alias "friend Standard_EXPORT Standard_Boolean operator ==(const Handle(Units_Quantity)&,const Standard_CString);"
    
    ---Purpose: Returns True if the name of the Quantity <me> is equal 
    --          to <astring>, False otherwise.
    
    is static;
    
    Dump(me ; ashift , alevel : Integer)
    
    ---Level: Internal 
    
    ---Purpose: Useful for debugging.
    
    is static;

fields

    thename          : HAsciiString  from TCollection;
    thedimensions    : Dimensions    from Units;
    theunitssequence : UnitsSequence from Units;

end Quantity;
