-- Created on: 1993-06-24
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class CurveTool from TopOpeBRepTool

uses

    Shape from TopoDS,
    Curve from Geom,
    Curve from Geom2d,
    Array1OfPnt from TColgp,
    Array1OfPnt2d from TColgp,
    GeomTool from TopOpeBRepTool,
    OutCurveType from TopOpeBRepTool
    
is

    Create returns CurveTool from TopOpeBRepTool;

    Create (OCT:OutCurveType from TopOpeBRepTool)
    returns CurveTool from TopOpeBRepTool;

    Create(GT:GeomTool from TopOpeBRepTool)
    returns CurveTool from TopOpeBRepTool;

    ChangeGeomTool(me:in out) returns GeomTool from TopOpeBRepTool is static;
    ---C++: return &
    GetGeomTool(me) returns GeomTool from TopOpeBRepTool is static;
    ---C++: return const &
    SetGeomTool(me:in out; GT:GeomTool from TopOpeBRepTool) is static;

    MakeCurves(me; 
    	       min,max:Real from Standard;
    	       C3D:Curve from Geom;
    	       PC1,PC2:Curve from Geom2d;
    	       S1,S2:Shape from TopoDS;
	       C3DN:out Curve from Geom;
    	       PC1N,PC2N:out Curve from Geom2d;
    	       Tol3d,Tol2d:out Real from Standard)
    returns Boolean from Standard is static;
    ---Purpose: Approximates curves.
    --          Returns False in the case of failure

    -- class methods

    MakeBSpline1fromPnt(myclass;P:Array1OfPnt from TColgp)
    returns Curve from Geom;  

    MakeBSpline1fromPnt2d(myclass;P:Array1OfPnt2d from TColgp)
    returns Curve from Geom2d;

    IsProjectable(myclass;S:Shape from TopoDS;C:Curve from Geom)
    returns Boolean;

    MakePCurveOnFace(myclass;
    	    	     S:Shape from TopoDS;
    	    	     C:Curve from Geom;
    	    	     TolReached2d : out Real from Standard;
		     first: Real from Standard = 0.0;
		     last: Real from Standard = 0.0)
    returns Curve from Geom2d;

fields 

    myGeomTool : GeomTool from TopOpeBRepTool is protected;

end CurveTool;
