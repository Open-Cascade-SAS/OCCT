-- Created on: 1995-09-21
-- Created by: Philippe GIRODENGO
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MeshExplorer from StlMesh 

	---Purpose: Provides  facilities to explore  the triangles  of
	--          each mesh domain.
	--          
uses  

    Mesh                   from StlMesh,
    SequenceOfMeshTriangle from StlMesh,
    SequenceOfXYZ          from TColgp

raises 

    OutOfRange   from Standard,
    NoMoreObject from Standard,
    NoSuchObject from Standard

is

    Create (M : Mesh)  returns MeshExplorer;
    

    Deflection (me) returns Real is static;
    	---Purpose: Returns the mesh deflection of the current domain.

    InitTriangle (me : in out; DomainIndex : Integer = 1)
    	---Purpose: Initializes the exploration  of the  triangles  of
    	--          the mesh domain of range <DomainIndex>.
    raises OutOfRange
    	---Purpose: Raised if <DomainIndex> is lower than 1 or greater
    	--          than the number of domains.
    is static;


    MoreTriangle (me) returns Boolean is static;
    	---C++: inline


    NextTriangle (me : in out) 
    raises NoMoreObject
    	---Purpose: Raised if there is no more triangle in the current
    	--          domain.
    is static;


    TriangleVertices (me; X1, Y1, Z1, X2, Y2, Z2, X3, Y3, Z3 : in out Real)
    raises NoSuchObject
    	---Purpose: Raised if there is no more triangle in the current
    	--          domain.
    is static;

   
    TriangleOrientation (me; Xn, Yn, Zn : in out Real)
    raises NoSuchObject
    	---Purpose: Raised if there is no more triangle in the current
    	--          domain.
    is static;



fields

    mesh            : Mesh;
    xn, yn, zn      : Real;
    v1, v2, v3      : Integer;
    domainIndex     : Integer;
    nbTriangles     : Integer;
    triangleIndex   : Integer;
    trianglesVertex : SequenceOfXYZ;
    trianglesdef    : SequenceOfMeshTriangle;

end MeshExplorer;







