-- Created on: 1993-02-22
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class LineOn2S from IntSurf 

	---Purpose: 

inherits TShared from MMgt


uses Allocator         from IntSurf,
     PntOn2S           from IntSurf,
     SequenceOfPntOn2S from IntSurf

raises OutOfRange from Standard

is

    Create (theAllocator: Allocator from IntSurf = 0)
    
    	returns mutable LineOn2S from IntSurf;
	

    Add(me: mutable; P: PntOn2S from IntSurf)
    
	---Purpose: Adds a point in the line.

	---C++: inline

    	is static;


    NbPoints(me)
    
	---Purpose: Returns the number of points in the line.

    	returns Integer from Standard
	---C++: inline
	
	is static;


    Value(me; Index: Integer from Standard)
    
	---Purpose: Returns the point of range Index in the line.
    
    	returns PntOn2S from IntSurf
	---C++: inline
	---C++: return const&
	
	raises OutOfRange from Standard
	--- The exception OutOfRange is raised when Index <= 0 or
	--  Index > NbPoints.
	
	is static;


    Reverse(me: mutable)
    
	---Purpose: Reverses the order of points of the line.

	---C++: inline

    	is static;



    Split(me: mutable;Index: Integer from Standard)

	---Purpose: Keeps in <me> the points 1 to Index-1, and returns
	--          the items Index to the end.

    	returns mutable LineOn2S from IntSurf

    	raises OutOfRange from Standard
	--- The exception OutOfRange is raised when Index <= 0 or
	--  Index > NbPoints.

	is static;


    Value(me: mutable; Index: Integer from Standard; P: PntOn2S from IntSurf)
    
	---Purpose: Replaces the point of range Index in the line.
    
	raises OutOfRange from Standard
	--- The exception OutOfRange is raised when Index <= 0 or
	--  Index > NbPoints.
	
	---C++: inline
        
	is static;
	
	
    SetUV(me: mutable; Index: Integer from Standard;
    	               OnFirst: Boolean from Standard;
		       U,V: Real from Standard)
    
	---Purpose: Sets the parametric coordinates on one of the surfaces
	--          of the point of range Index in the line.
    
	---C++: inline
        
	raises OutOfRange from Standard
	--- The exception OutOfRange is raised when Index <= 0 or
	--  Index > NbPoints.
	
	is static;
	
	
    Clear(me: mutable)
    
	---C++: inline
        
    	is static;


    InsertBefore(me:mutable; I: Integer from Standard; P: PntOn2S from IntSurf) 
    
    	is static;

    RemovePoint(me:mutable; I: Integer from Standard)
    
    	is static;


fields

    mySeq: SequenceOfPntOn2S from IntSurf;

end LineOn2S;
