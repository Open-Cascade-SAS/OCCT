-- Created on: 1996-09-25
-- Created by: Christian CAILLET
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SelectSignedSharing  from IFSelect  inherits SelectExplore

    ---Purpose : In the graph, explore the sharings of the input entities,
    --           until it encounters some which match a given Signature
    --           (for a limited level, filters the returned list)
    --           By default, fitted for any level

uses AsciiString, Transient,  Graph, EntityIterator, Signature

is

    Create (matcher : Signature;
            signtext : CString;
            exact : Boolean = Standard_True;
   	    level : Integer = 0)  returns mutable SelectSignedSharing;
    ---Purpose : Creates a SelectSignedSharing, defaulted for any level
    --           with a given Signature and text to match

    Signature (me) returns mutable Signature;
    ---Purpose : Returns the used Signature, then it is possible to access it,
    --           modify it as required

    SignatureText (me) returns AsciiString from TCollection;
    ---Purpose : Returns Text used to Sort Entity on its Signature
    ---C++ : return const &

    IsExact (me) returns Boolean;
    ---Purpose : Returns True if match must be exact

    Explore (me; level : Integer; ent : Transient; G : Graph;
    	     explored : in out EntityIterator)
    	returns Boolean;
    ---Purpose : Explores an entity : its sharing entities
    --           <ent> to take if it matches the Signature
    --           At level max, filters the result. Else gives all sharings


    ExploreLabel (me) returns AsciiString from TCollection;
    ---Purpose : Returns a text defining the criterium.
    --           (it refers to the text and exact flag to be matched, and is
    --           qualified by the Name provided by the Signature)

fields
 
    thematcher  : Signature;
    thesigntext : AsciiString from TCollection;
    theexact    : Boolean;

end SelectSignedSharing;
