-- Created on: 1999-03-09
-- Created by: data exchange team
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class DateItem from StepAP214 inherits ApprovalItem from StepAP214


uses
    	ApprovalPersonOrganization from StepBasic,
	AppliedPersonAndOrganizationAssignment from StepAP214,
    	AppliedOrganizationAssignment from StepAP214,
    	Effectivity from StepBasic

is
    Create returns DateItem;
	---Purpose : Returns a DateItem SelectType
	
	CaseNum (me; ent : Transient) returns Integer is redefined;
	---Purpose: Recognizes a DateItem Kind Entity that is :
	--        1 -> ApprovalPersonOrganization
	--        2 -> AppliedDateAndPersonAssignment
    	--        3 -> AppliedOrganizationAssignment
    	--        4 -> AssemblyComponentUsageSubstitute
	--        5 -> DocumentFile
	--        6 -> Effectivity
    	--        7 -> MaterialDesignation
    	--        8 -> MechanicalDesignGeometricPresentationRepresentation
	--        9 -> PresentationArea
    	--        10 -> Product
	--        11 -> ProductDefinition
    	--        12 -> ProductDefinitionFormation
	--        13 -> ProductDefinitionRelationship
    	--    	  14 -> PropertyDefinition
    	--        15 -> ShapeRepresentation
	--        0 else

	ApprovalPersonOrganization (me) returns any ApprovalPersonOrganization ;
	---Purpose : returns Value as a ApprovalPersonOrganization (Null if another type)

	AppliedPersonAndOrganizationAssignment (me) returns any AppliedPersonAndOrganizationAssignment ; 
	---Purpose : returns Value as a AppliedDateAndPersonAssignment (Null if another type)

    	AppliedOrganizationAssignment (me) returns any AppliedOrganizationAssignment ;
    	---Purpose : returns Value as a AppliedOrganizationAssignment (Null if another type)

	Effectivity (me) returns any Effectivity ;
	---Purpose : returns Value as a Effectivity (Null if another type)
	

end DateItem;
