-- File:	MakeCylindricalSurface.cdl
-- Created:	Mon Sep 28 11:51:29 1992
-- Author:	Remi GILET
--		<reg@sdsun2>
---Copyright:	 Matra Datavision 1992

class MakeCylindricalSurface from GC inherits Root from GC

    ---Purpose : This class implements the following algorithms used 
    --           to create a CylindricalSurface from Geom.
    --           * Create a CylindricalSurface parallel to another and 
    --           passing through a point.
    --           * Create a CylindricalSurface parallel to another at a 
    --           distance
    --             <Dist>.
    --           * Create a CylindricalSurface passing through 3 points.
    --           * Create a CylindricalSurface by its axis and radius.
    --           * Create a cylindricalSurface by its circular base.
    --  The local coordinate system of the CylindricalSurface is defined
    --  with an axis placement (see class ElementarySurface).
    --  
    --  The "ZAxis" is the symmetry axis of the CylindricalSurface, 
    --  it gives the direction of increasing parametric value V.
    --  
    --  The parametrization range is :
    --       U [0, 2*PI],  V ]- infinite, + infinite[
    --       
    --  The "XAxis" and the "YAxis" define the placement plane of the 
    --  surface (Z = 0, and parametric value V = 0)  perpendicular to 
    --  the symmetry axis. The "XAxis" defines the origin of the 
    --  parameter U = 0.  The trigonometric sense gives the positive 
    --  orientation for the parameter U.

uses Pnt                from gp,
     Ax1                from gp,
     Ax2                from gp,
     Circ               from gp,
     Cylinder           from gp,
     CylindricalSurface from Geom,
     Real               from Standard

raises NotDone from StdFail

is

Create (A2 : Ax2; Radius : Real) returns MakeCylindricalSurface;
    --- Purpose :
    --  A2 defines the local coordinate system of the cylindrical surface.
    --  The "ZDirection" of A2 defines the direction of the surface's
    --  axis of symmetry.
    --  At the creation the parametrization of the surface is defined
    --  such that the normal Vector (N = D1U ^ D1V) is oriented towards
    --  the "outside region" of the surface.
    -- Warnings :
    --  It is not forbidden to create a cylindrical surface with 
    --  Radius = 0.0
    --- Status is "NegativeRadius" if Radius < 0.0

Create (C : Cylinder from gp)  returns MakeCylindricalSurface;
    --- Purpose :
    --  Creates a CylindricalSurface from a non persistent Cylinder
    --  from package gp.

Create(Cyl   : Cylinder from gp;
       Point : Pnt      from gp) returns MakeCylindricalSurface;
    ---Purpose : Make a CylindricalSurface from Geom <TheCylinder> 
    --           parallel to another 
    --           CylindricalSurface <Cylinder> and passing through a 
    --           Pnt <Point>.

Create(Cyl  : Cylinder  from gp      ;
       Dist : Real      from Standard) returns MakeCylindricalSurface;
    ---Purpose : Make a CylindricalSurface from Geom <TheCylinder> 
    --           parallel to another 
    --           CylindricalSurface <Cylinder> at the distance <Dist> 
    --           which can be greater or lower than zero.
    --           The radius of the result is the absolute value of the
    --           radius of <Cyl> plus <Dist>

Create(P1     :     Pnt from gp;
       P2     :     Pnt from gp;
       P3     :     Pnt from gp) returns MakeCylindricalSurface;
    ---Purpose : Make a CylindricalSurface from Geom <TheCylinder> 
    --           passing through 3 Pnt <P1>,<P2>,<P3>.
    --           Its axis is <P1P2> and its radius is the distance 
    --           between <P3> and <P1P2>

Create(Axis   : Ax1  from gp      ;
       Radius : Real from Standard) returns MakeCylindricalSurface;
    ---Purpose: Make a CylindricalSurface by its axis <Axis> and radius 
    --          <Radius>.

Create(Circ   : Circ from gp) returns MakeCylindricalSurface;
    ---Purpose: Make a CylindricalSurface by its circular base.

Value(me) returns CylindricalSurface from Geom
    raises NotDone
    is static;
    ---Purpose: Returns the constructed cylinder.
    -- Exceptions StdFail_NotDone if no cylinder is constructed.
    ---C++: return const&

Operator(me) returns CylindricalSurface from Geom
    is static;
    ---C++: return const&
    ---C++: alias "Standard_EXPORT operator Handle_Geom_CylindricalSurface() const;"

fields

    TheCylinder : CylindricalSurface from Geom;
    --The solution from Geom.
    
end MakeCylindricalSurface;




