-- Created on: 1995-01-09
-- Created by: Modelistation
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Wedge from BRepPrim inherits GWedge from BRepPrim

	---Purpose: Provides constructors without Builders.

uses
    Ax2 from gp,
    Pnt from gp

raises
    DomainError

is

    Create(Axes : Ax2 from gp; dx, dy, dz : Real)
    returns Wedge from BRepPrim
	---Purpose: Creates a  Wedge  algorithm.   <Axes> is  the axis
	--          system for the primitive.
	--          
	--          XMin, YMin, ZMin are set to 0
	--          XMax, YMax, ZMax are set to dx, dy, dz
	--          Z2Min = ZMin
	--          Z2Max = ZMax
	--          X2Min = XMin
	--          X2Max = XMax
	--          The result is a box
	--          dx,dy,dz should be positive
	raises DomainError;

    Create(Axes : Ax2 from gp; dx, dy, dz, ltx : Real)
    returns Wedge from BRepPrim
	---Purpose: Creates  a Wedge  primitive. <Axes> is   the  axis
	--          system for the primitive.
	--          
	--          XMin, YMin, ZMin are set to 0
	--          XMax, YMax, ZMax are set to dx, dy, dz
	--          Z2Min = ZMin
	--          Z2Max = ZMax
	--          X2Min = ltx
	--          X2Max = ltx
	--          The result is a STEP right angular wedge
	--          dx,dy,dz should be positive
	--          ltx should not be negative
	raises DomainError;

    Create(Axes : Ax2 from gp; xmin, ymin, zmin, z2min, x2min,
                                   xmax, ymax, zmax, z2max, x2max : Real)
    returns Wedge from BRepPrim
	---Purpose: Create  a Wedge primitive.   <Axes>  is  the  axis
	--          system for the primitive.
	--          
	--          all the fields are set to the corresponding value
	--          XYZMax - XYZMin should be positive
	--          ZX2Max - ZX2Min should not be negative 
	raises DomainError;

end Wedge;
