-- File:	IGESDimen_SpecificModule.cdl
-- Created:	Tue Sep  7 11:14:37 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class SpecificModule  from IGESDimen  inherits  SpecificModule from IGESData

    ---Purpose : Defines Services attached to IGES Entities :
    --           Dump & OwnCorrect, for IGESDimen

uses Messenger from Message, IGESEntity, IGESDumper

is

    Create returns mutable SpecificModule from IGESDimen;
    ---Purpose : Creates a SpecificModule from IGESDimen & puts it into SpecificLib

    OwnDump (me; CN : Integer; ent : IGESEntity;
    	      dumper : IGESDumper;  S : Messenger from Message; own : Integer);
    ---Purpose : Specific Dump (own parameters) for IGESDimen

    OwnCorrect (me; CN : Integer; ent : mutable IGESEntity)
    	returns Boolean  is redefined;
    ---Purpose : Performs non-ambiguous Corrections on Entities which support
    --           them (BasicDimension,CenterLine,DimensionDisplayData,
    --           DimensionTolerance,DimensionUnits,DimensionedGeometry,
    --           NewDimensionedGeometry,Section,WitnessLine)

end SpecificModule;
