-- File:	StepAP203_StartRequest.cdl
-- Created:	Fri Nov 26 16:26:40 1999 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0
-- Copyright:	Matra Datavision 1999

class StartRequest from StepAP203
inherits ActionRequestAssignment from StepBasic

    ---Purpose: Representation of STEP entity StartRequest

uses
    VersionedActionRequest from StepBasic,
    HArray1OfStartRequestItem from StepAP203

is
    Create returns StartRequest from StepAP203;
	---Purpose: Empty constructor

    Init (me: mutable; aActionRequestAssignment_AssignedActionRequest: VersionedActionRequest from StepBasic;
                       aItems: HArray1OfStartRequestItem from StepAP203);
	---Purpose: Initialize all fields (own and inherited)

    Items (me) returns HArray1OfStartRequestItem from StepAP203;
	---Purpose: Returns field Items
    SetItems (me: mutable; Items: HArray1OfStartRequestItem from StepAP203);
	---Purpose: Set field Items

fields
    theItems: HArray1OfStartRequestItem from StepAP203;

end StartRequest;
