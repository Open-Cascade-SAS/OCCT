-- Created on: 1996-01-12
-- Created by: Denis PASCAL
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PlanarAngle from DrawDim inherits PlanarDimension from DrawDim

	---Purpose: 

uses Shape    from TopoDS,
     Face    from TopoDS,
     Color   from Draw,
     Display from Draw

is

    Create (plane : Face  from TopoDS;
            line1 : Shape from TopoDS; 
            line2 : Shape from TopoDS)
    returns PlanarAngle from DrawDim;    

    Create (line1 : Shape from TopoDS; 
            line2 : Shape from TopoDS)
    returns PlanarAngle from DrawDim;
    
    Sector (me : mutable; inverted, reversed : Boolean from Standard);
    
    Position (me : mutable; value : Real from Standard);
    
    DrawOn (me; dis : in out Display);
    
fields

    myLine1 : Shape from TopoDS;
    myLine2 : Shape from TopoDS;
    myIsReversed : Boolean from Standard;
    myIsInverted : Boolean from Standard;
    myPosition   : Real from Standard; -- par rapport au point d'intersection    	    
		
end PlanarAngle;

