-- Created on: 2004-03-05
-- Created by: Mikhail KUZMITCHEV
-- Copyright (c) 2004-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package QANCollection

uses
    Draw,
    TCollection, 
    TColStd,
    gp

is
    imported ListOfPnt;
    imported ListIteratorOfListOfPnt;
    imported DataMapOfRealPnt;
    imported DataMapIteratorOfDataMapOfRealPnt;
    imported IndexedDataMapOfRealPnt;
    imported DoubleMapOfRealInteger;
    imported DoubleMapIteratorOfDoubleMapOfRealInteger;

    Commands(DI : in out Interpretor from Draw);
    CommandsSimple(DI : in out Interpretor from Draw);
    CommandsTest(DI : in out Interpretor from Draw);
    CommandsPerf(DI : in out Interpretor from Draw);
    CommandsAlloc(DI : in out Interpretor from Draw);
    CommandsStl(DI : in out Interpretor from Draw);

end;
