-- Created on: 1997-01-09
-- Created by: Yves FRICAUD
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



private class ShapesSet from TNaming 

	---Purpose: 

uses
    Shape                   from TopoDS,
    ShapeEnum               from TopAbs,
    MapOfShape              from TopTools

is
    Create returns ShapesSet from TNaming;
    	---C++: inline

    Create (S    : Shape        from TopoDS;
    	    Type : ShapeEnum    from TopAbs = TopAbs_SHAPE)
    returns ShapesSet from TNaming;

---Category: Modification
   
    Clear(me : in out)
	---Level: Public
	---Purpose: Removes all Shapes
	---C++: inline
    is static;
    
    Add(me : in out; S : Shape from TopoDS) returns Boolean
	---Level: Public
	---Purpose: Adds the Shape <S>
	---C++: inline
    is static;

    Contains(me; S : Shape ) returns Boolean
	---Level: Public
	---Purpose: Returns True  if <S> is in <me>
	---C++: inline
    is static;
    
    Remove(me : in out; S : Shape ) returns Boolean
	---Level: Public
	---Purpose: Removes <S> in <me>.
        ---C++: inline
    is static;


    -- Modification with an other ShapesSet--

    Add    (me : in out; Shapes : ShapesSet from TNaming);
    	---Purpose: Adds the shapes contained in <Shapes>.
    
    Filter (me : in out; Shapes : ShapesSet from TNaming);
      	---Purpose: Erases in <me> the shapes not 
     	--          contained in <Shapes>

               
    Remove (me : in out; Shapes : ShapesSet from TNaming);
    	---Purpose: Removes in <me> the shapes contained in <Shapes>


---Category: Querying
    
    IsEmpty(me) returns Boolean from Standard;
    	---C++: inline

    NbShapes (me) returns Integer from Standard;   
    	---C++: inline

    ChangeMap(me: in out) returns MapOfShape from TopTools;
    	---C++: return &
    	---C++: inline

    Map(me) returns MapOfShape from TopTools;
    	---C++: return const&
    	---C++: inline

fields
    myMap   : MapOfShape              from TopTools;

end ShapesSet;


