-- Created on: 1997-12-08
-- Created by: Serguei ZARITCHNY
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class FilletRadiusPresentation from DsgPrs

        ---Purpose: A framework for displaying radii of fillets.
uses
    Presentation from Prs3d,
    Pnt from gp,
    Dir from gp,
    Drawer from Prs3d,
    ExtendedString from TCollection,
    ArrowSide from DsgPrs,
    TrimmedCurve from Geom,
    Circle  from Geom,
    Ax1 from gp
is
    Add( myclass; aPresentation : Presentation from Prs3d;
    	    	  aDrawer       : Drawer from Prs3d;
		  thevalue      : Real from Standard;
		  aText         : ExtendedString from TCollection;
		  aPosition     : Pnt from gp;
		  aNormalDir    : Dir from gp;
		  aBasePnt      : Pnt from gp;
		  aFirstPoint   : Pnt from gp;
		  aSecondPoint  : Pnt from gp;
		  aCenter       : Pnt from gp;
		  ArrowPrs      : ArrowSide from DsgPrs; 
		  drawRevers    : Boolean from Standard; 
    	    	  DrawPosition  : out Pnt from gp;
    	    	  EndOfArrow    : out Pnt from gp;
    	    	  TrimCurve     : out TrimmedCurve from Geom;
    	    	  HasCircle     : out Boolean from Standard);
    	---Purpose: Adds a display of the radius of a fillet to the
    	-- presentation aPresentation. The display ttributes
    	-- defined by the attribute manager aDrawer. the value
    	-- specifies the length of the radius.
		  
end FilletRadiusPresentation;
