-- Created on: 1995-07-24
-- Created by: Modelistation
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Plane from StdPrs
	 
inherits Root from Prs3d

    	---Purpose: A framework to display infinite planes.
          
uses 
    Surface           from Adaptor3d,
    Presentation      from Prs3d,
    Drawer            from Prs3d,
    TypeOfLinePicking from Prs3d,
    Length            from Quantity
    
is
    Add(myclass; aPresentation: Presentation from Prs3d; 
         	 aPlane       : Surface      from Adaptor3d;
    	    	 aDrawer      : Drawer       from Prs3d);
		 
    	---Purpose: Defines display of infinite planes.
    	-- The infinite plane aPlane is added to the display
    	-- aPresentation, and the attributes of the display are
    	-- defined by the attribute manager aDrawer.

    Match(myclass; X,Y,Z   : Length  from Quantity;
    	          aDistance: Length  from Quantity;
                  aPlane   : Surface from Adaptor3d;
    	          aDrawer  : Drawer  from Prs3d)
    returns Boolean from Standard;

    	---Purpose: returns true if the distance between the point (X,Y,Z) and the
    	--          plane is less than aDistance.


end Plane;
