-- Created on: 1991-02-27
-- Created by: Jean Claude Vauthier
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class UniformDeflection from CPnts 
 
        ---Purpose : This classe defines an algorithm to create a set of points at the
        --  positions of constant deflection of a given curve or a trimmed 
        --  circle.
        --  The continuity of the curve must be at least C2.
        --
        --  the usage of the is the following.
        --          
        --  class myUniformDFeflection instantiates
        --                     UniformDeflection(Curve, Tool);
        --
        --      
        -- Curve C; // Curve inherits from Curve or Curve2d from Adaptor2d
        -- myUniformDeflection Iter1;
        -- DefPntOfmyUniformDeflection P;
        --        
        -- for(Iter1.Initialize(C, Deflection, EPSILON, True); 
        --     Iter1.More();
        --     Iter1.Next()) {
        --   P = Iter1.Value();
        --   ... make something with P
        -- }
        -- if(!Iter1.IsAllDone()) {
        --    ... something wrong happened 
        -- }
uses
    Curve   from Adaptor3d,
    Curve2d from Adaptor2d,
    Pnt     from gp

raises DomainError from Standard, 
       NotDone     from StdFail, 
       OutOfRange  from Standard

is


        --        
  
  Create 
  ---Purpose: creation of a indefinite UniformDeflection
  returns UniformDeflection;

  Create(C : Curve from Adaptor3d; Deflection,  Resolution  : Real; 
                                 WithControl : Boolean )
        --- Purpose :  Computes a uniform deflection distribution of points
        --  on the curve <C>.
        --  <Deflection> defines the constant deflection value.
        --  The algorithm computes the number of points and the points.
        --  The curve <C> must be at least C2 else the computation can fail.
        --  If just some parts of the curve is C2 it is better to give the 
        --  parameters bounds and to use the below constructor .
        --  if <WithControl> is True, the algorithm controls the estimate 
        --  deflection
        --  when the curve is singular at the point P(u),the algorithm 
        --  computes the next point as  
        --  P(u + Max(CurrentStep,Abs(LastParameter-FirstParameter)))
        --  if the singularity is at the first point ,the next point
        --  calculated is the P(LastParameter)   
     returns UniformDeflection;

  Create(C : Curve2d from Adaptor2d; Deflection,  Resolution  : Real; 
                                   WithControl : Boolean )
	---Purpose: As above with 2d curve
     returns UniformDeflection;

  Create(C : Curve from Adaptor3d; Deflection, U1, U2, Resolution : Real; 
                    WithControl : Boolean)
        --- Purpose :
        --  Computes an uniform deflection distribution of points on a part of
        --  the curve <C>. Deflection defines the step between the points.
        --  <U1> and <U2> define the distribution span. 
        --  <U1> and <U2> must be in the parametric range of the curve.
     returns UniformDeflection
     raises DomainError;
        --  raised if U1 and U2 are not in the parametric bounds of the curve.

  Create(C : Curve2d from Adaptor2d; Deflection, U1, U2, Resolution : Real; 
                    WithControl : Boolean)
        --- Purpose : As above with 2d curve
     returns UniformDeflection
     raises DomainError;
        --  raised if U1 and U2 are not in the parametric bounds of the curve.

    Initialize(me : in out; C : Curve from Adaptor3d; 
                            Deflection, Resolution : Real; 
                            WithControl : Boolean)
    	---Purpose: Initialize the algoritms with <C>, <Deflection>, <UStep>,
    	--          <Resolution> and <WithControl>
        is static;
     
    Initialize(me : in out; C : Curve2d from Adaptor2d; 
                            Deflection, Resolution : Real; 
                            WithControl : Boolean)
    	---Purpose: Initialize the algoritms with <C>, <Deflection>, <UStep>,
    	--          <Resolution> and <WithControl>
        is static;
     
    Initialize(me : in out; C : Curve from Adaptor3d; 
                            Deflection, U1, U2, Resolution : Real; 
                            WithControl : Boolean)
    	---Purpose: Initialize the algoritms with <C>, <Deflection>, <UStep>,
    	--          <U1>, <U2> and <WithControl>
     	raises DomainError
	is static;
  
    Initialize(me : in out; C : Curve2d from Adaptor2d; 
                            Deflection, U1, U2, Resolution : Real; 
                            WithControl : Boolean)
    	---Purpose: Initialize the algoritms with <C>, <Deflection>, <UStep>,
    	--          <U1>, <U2> and <WithControl>
     	raises DomainError
	is static;
  
    IsAllDone (me)
        --- Purpose : To know if all the calculus were done successfully
        --  (ie all the points have been computed). The calculus can fail if
        --  the Curve is not C1 in the considered domain.
        --  Returns True if the calculus was successful.
        ---C++: inline
        returns Boolean
     	is static;

    Next(me : in out)
        ---Purpose: go to the next Point.
        ---C++: inline
    	raises OutOfRange
    	is static;  

    More(me : in out)
        ---Purpose: returns True if it exists a next Point.
    	returns Boolean
      	is static;
  
    Value(me) returns Real
        ---Purpose : return the computed parameter
        ---C++: inline
    	is static;


    Point(me) returns Pnt from gp
        ---Purpose : return the computed parameter
        ---C++: inline
    	is static;
	
    Perform (me : in out)  
        ---Purpose: algorithm 
    	is static private;
	
fields

    myDone       : Boolean;
    my3d         : Boolean;
    myCurve      : Address from Standard;
    myFinish     : Boolean;
    myTolCur     : Real;
    myControl    : Boolean;
    myIPoint     : Integer;
    myNbPoints   : Integer;
    myParams     : Real[3];
    myPoints     : Pnt from gp [3] ;
    myDwmax      : Real;
    myDeflection : Real;
    myFirstParam : Real;
    myLastParam  : Real;
    myDu         : Real;
    
end UniformDeflection;





