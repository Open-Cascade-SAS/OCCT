-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class TrimmedCurve from StepGeom 

inherits BoundedCurve from StepGeom 

uses

	Curve from StepGeom, 
	HArray1OfTrimmingSelect from StepGeom, 
	Boolean from Standard, 
	TrimmingPreference from StepGeom, 
	TrimmingSelect from StepGeom, 
	HAsciiString from TCollection
is

	Create returns mutable TrimmedCurve;
	---Purpose: Returns a TrimmedCurve


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aBasisCurve : mutable Curve from StepGeom;
	      aTrim1 : mutable HArray1OfTrimmingSelect from StepGeom;
	      aTrim2 : mutable HArray1OfTrimmingSelect from StepGeom;
	      aSenseAgreement : Boolean from Standard;
	      aMasterRepresentation : TrimmingPreference from StepGeom) is virtual;

	-- Specific Methods for Field Data Access --

	SetBasisCurve(me : mutable; aBasisCurve : mutable Curve);
	BasisCurve (me) returns mutable Curve;
	SetTrim1(me : mutable; aTrim1 : mutable HArray1OfTrimmingSelect);
	Trim1 (me) returns mutable HArray1OfTrimmingSelect;
	Trim1Value (me; num : Integer) returns TrimmingSelect;
	NbTrim1 (me) returns Integer;
	SetTrim2(me : mutable; aTrim2 : mutable HArray1OfTrimmingSelect);
	Trim2 (me) returns mutable HArray1OfTrimmingSelect;
	Trim2Value (me; num : Integer) returns TrimmingSelect;
	NbTrim2 (me) returns Integer;
	SetSenseAgreement(me : mutable; aSenseAgreement : Boolean);
	SenseAgreement (me) returns Boolean;
	SetMasterRepresentation(me : mutable; aMasterRepresentation : TrimmingPreference);
	MasterRepresentation (me) returns TrimmingPreference;

fields

	basisCurve : Curve from StepGeom;
	trim1 : HArray1OfTrimmingSelect from StepGeom; -- a SelectType
	trim2 : HArray1OfTrimmingSelect from StepGeom; -- a SelectType
	senseAgreement : Boolean from Standard;
	masterRepresentation : TrimmingPreference from StepGeom; -- an Enumeration

end TrimmedCurve;
