-- Created on: 1992-11-17
-- Created by: Christian CAILLET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class SelectionIterator  from IFSelect

    ---Purpose : Defines an Iterator on a list of Selections

uses Selection, HSeqOfSelection, TSeqOfSelection

raises NoSuchObject

is

    Create  returns SelectionIterator;
    ---Purpose : Creates an empty iterator, ready to be filled

    Create (sel : Selection) returns SelectionIterator;
    ---Purpose : Creates an iterator from a Selection : it lists the Selections
    --           from which <sel> depends (given by its method FillIterator)

    AddFromIter (me : in out;  iter : in out SelectionIterator)  is static;
    ---Purpose : Adds to an iterator the content of another one
    --           (each selection is present only once in the result)

    AddItem     (me : in out; sel : any Selection)               is static;
    ---Purpose : Adds a Selection to an iterator (if not yet noted)

    AddList     (me : in out; list : TSeqOfSelection)            is static;
    ---Purpose : Adds a list of Selections to an iterator (this list comes
    --           from the description of a Selection or a Dispatch, etc...)


    More (me) returns Boolean  is static;
    ---Purpose : Returns True if there are more Selections to get

    Next (me : in out)  is static;
    ---Purpose : Sets iterator to the next item

    Value (me) returns any Selection  raises NoSuchObject  is static;
    ---Purpose : Returns the current Selction beeing iterated
    --           Error if count of Selection has been passed
    ---C++ : return const &

fields

    thecurr : Integer;
    thelist : HSeqOfSelection;

end SelectionIterator;
