-- Created on: 1995-12-04
-- Created by: Laurent BOURESCHE
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class TgtField from GeomFill inherits TShared from MMgt

	---Purpose: Root class defining the methods we need to make an
	--          algorithmic tangents field.

uses
    Vec from gp,
    BSpline from Law

is

    IsScalable(me) returns Boolean from Standard is virtual;
    Scale(me : mutable; Func : BSpline from Law) is virtual;

    Value(me; W : Real from Standard)
    returns Vec from gp
    ---Purpose: Computes  the value  of the    field of tangency    at
    --          parameter W.
    is deferred;

    D1(me; W : Real from Standard)
    returns Vec from gp
    ---Purpose: Computes the  derivative of  the field of  tangency at
    --          parameter W.
    is deferred;

    D1(me; W : Real from Standard; V, DV : out Vec from gp)
    ---Purpose: Computes the value and the  derivative of the field of
    --          tangency at parameter W.
    is deferred;

end TgtField;
