-- File:	QANewModTopOpe_ReShaper.cdl
-- Created:	Thu Feb  7 12:05:56 2002
-- Author:	Igor FEOKTISTOV <ifv@nnov.matra-dtv.fr>
-- Copyright:	SAMTECH S.A. 2002

-- Lastly modified by :
-- +---------------------------------------------------------------------------+
-- !       ifv ! Creation                                ! 7-02-2002! 3.0-00-1!
-- +---------------------------------------------------------------------------+

class ReShaper from QANewModTopOpe inherits TShared from  MMgt 
    	---Purpose: to remove  "floating" objects from compound.
	-- "floating" objects are wires, edges, vertices that do not belong
	-- solids, shells or faces.

uses 
    Shape from TopoDS, 
    HSequenceOfShape  from  TopTools, 
    MapOfShape  from  TopTools 
is 
 
    Create(TheInitialShape  :  Shape from TopoDS) 
     
    returns  mutable  ReShaper; 
     
    Create(TheInitialShape  :  Shape from TopoDS;   
    	   TheMap  :  MapOfShape  from  TopTools) 
     
    returns  mutable  ReShaper; 
     
    Create(TheInitialShape  :  Shape from TopoDS;   
           TheShapeToBeRemoved  : HSequenceOfShape  from  TopTools) 
     
    returns  mutable  ReShaper; 
     
    Remove(me  :  mutable;  TheS  :  Shape from TopoDS); 
     
    Perform(me  :  mutable); 
     
    Clear(me  :  mutable);  
    ---Purpose:  to  clear  all  added  for  removing  shapes  from  inner  map.
     
    GetResult(me)  returns  Shape  from  TopoDS; 
	---C++: return const &
	---C++: alias "Standard_EXPORT operator TopoDS_Shape() const;"
     
fields 
 
    myInitShape  :  Shape  from  TopoDS; 
    myResult     :  Shape  from  TopoDS;  
    myMap        :  MapOfShape  from  TopTools;  
    
end;    

-- @@SDM: begin

-- Copyright SAMTECH ..........................................Version    3.0-00
-- Lastly modified by : ifv                                    Date :  7-02-2002

-- File history synopsis (creation,modification,correction)
-- +---------------------------------------------------------------------------+
-- ! Developer !              Comments                   !   Date   ! Version  !
-- +-----------!-----------------------------------------!----------!----------+
-- !       ifv ! Creation                                ! 7-02-2002! 3.0-00-1!
-- +---------------------------------------------------------------------------+

-- @@SDM: end
