-- Created by: DAUTRY Philippe
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

--      	----------------

---Version:	0.0
--Version	Date		Purpose
--		0.0	Mar 11 1997	Creation


class CopyTool from TDF

	---Purpose: This class provides services to build, copy or
	--          paste a set of information.
	--          
	--          Copy methods:
	--          -------------
	--          
	--          * Copy(aSourceDataSet, aTargetLabel,
	--          aRelocationTable) copies a source DataSet under
	--          its target place (see below: IMPORTANT NOTICE 1).
	--          
	--          * Copy(aSourceDataSet, anTargetLabel,
	--          aRelocationTable, aFilter) does the same job as
	--          the previous method. But <aFilter> gives a list of
	--          IDs for which a target attribute prevails over a
	--          source one. In this special case, the source
	--          attribute will be copied only if there will be no
	--          target attribute.
	--          
	--          
	--          IMPORTANT NOTICE : Label pre-binding
	--          ------------------
	--          
	--          For it is possible to copy root labels in another
	--          place in the same Data or in a different one with
	--          other tags, it is necessary to inform the Copy
	--          algorithm about the target place. To do so:
	--          
	--          * first get or create new target root labels;
	--          
	--          * then bind them with the source root labels using
	--          the relocation table method:
	--          SetRelocation(aSourceLabel, aTargetLabel);
	--          
	--          * finally call Copy(...) with the relocation table
	--          previously set. In this way, this method will take
	--          these relocations in account.


uses

    Boolean             from Standard,
    Label               from TDF,
    Attribute           from TDF,
    DataSet             from TDF,
    RelocationTable     from TDF,
    AttributeMap        from TDF,
    AttributeDataMap    from TDF,
    LabelDataMap        from TDF,
    LabelMap            from TDF,
    IDFilter            from TDF,
    ClosureMode         from TDF


is

    Copy(myclass;
    	 aSourceDataSet   : DataSet from TDF;
	 aRelocationTable : mutable RelocationTable from TDF);
	---Purpose:  Copy   <aSourceDataSet> with using  and  updating
	--           <aRelocationTable>. This  method ignores   target
	--          attributes privilege over source ones.

    Copy(myclass;
    	 aSourceDataSet   : DataSet from TDF;
	 aRelocationTable : mutable RelocationTable from TDF;
    	 aPrivilegeFilter : IDFilter from TDF);
	---Purpose:    Copy  <aSourceDataSet>  using      and updating
	--          <aRelocationTable>. Use <aPrivilegeFilter> to give
	--           a list  of   IDs for which  the target  attribute
	--          prevails over the source one.


    -- Copy method piloting self contained attitude.
    -- ----------------------------------------------

    Copy(myclass;
    	 aSourceDataSet   : DataSet from TDF;
	 aRelocationTable : mutable RelocationTable from TDF;
    	 aPrivilegeFilter : IDFilter from TDF;
    	 aRefFilter       : IDFilter from TDF;
    	 setSelfContained : Boolean from Standard);
	---Purpose:   Copy    <aSourceDataSet>   using and    updating
	--          <aRelocationTable>. Use <aPrivilegeFilter> to give
	--           a  list of IDs   for which  the target  attribute
	--             prevails    over    the    source     one.   If
	--            <setSelfContained>   is   set  to   true,  every
	--          TDF_Reference will  be replaced  by the referenced
	--          structure according to <aRefFilter>.
	--          
	--          NB: <aRefFilter> is used only if
	--          <setSelfContained> is true.



    -- ----------------------------------------------------------------------
    -- 
    -- Private methods
    -- 
    -- ----------------------------------------------------------------------

    
    ---Purpose: Internal root label copy recursive method.    
    CopyLabels(myclass;
    	       aSLabel          : Label from TDF;
	       aTargetLabel     : in out Label from TDF;
	       aLabMap          : in out LabelDataMap from TDF;
	       aAttMap          : in out AttributeDataMap from TDF;
    	       aSrcLabelMap     : LabelMap from TDF;
    	       aSrcAttributeMap : AttributeMap from TDF)
    is private;

    ---Purpose: Internal root label copy recursive method.
    CopyAttributes(myclass;
    	    	   aSLabel          : Label from TDF;
    	    	   aTargetLabel     : in out Label from TDF;
    	    	   aAttMap          : in out AttributeDataMap from TDF;
    	    	   aSrcAttributeMap : AttributeMap from TDF)
    is private;
    ---Purpose: Internal attribute copy method.


end CopyTool;
