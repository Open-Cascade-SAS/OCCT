-- Created by: Peter KURNEV
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Point from BOPDS 

	---Purpose: 
    	-- The class BOPDS_Point is to store  
    	-- the information about intersection point 
uses
    Pnt from gp, 
    Pnt2d from gp 
    
--raises

is 
    Create 
    	returns Point from BOPDS; 
    ---C++: alias "virtual ~BOPDS_Point();" 
    ---C++: inline 
    	---Purpose:  
    	--- Empty contructor  
    	---  
	
    SetPnt(me:out; 
    	    thePnt:Pnt from gp); 
    ---C++: inline 
    	---Purpose: 
    	--- Modifier   
	--- Sets 3D point <thePnt>  
	
    Pnt(me)  
    	returns Pnt from gp; 
    ---C++: return const & 
    ---C++: inline  
    	---Purpose: 
    	--- Selector   
	--- Returns 3D point 
    
    SetPnt2D1(me:out; 
    	    thePnt:Pnt2d from gp); 
    ---C++: inline	 
     	---Purpose: 
    	--- Modifier   
	--- Sets 2D point on the first face <thePnt> 
	 
    Pnt2D1(me)  
    	returns Pnt2d from gp; 
    ---C++: return const & 
    ---C++: inline  
    	---Purpose: 
    	--- Selector 
	--- Returns 2D point on the first face <thePnt> 
    SetPnt2D2(me:out; 
    	    thePnt:Pnt2d from gp); 
    ---C++: inline 
    	---Purpose: 
    	--- Modifier   
	--- Sets 2D point on the second face <thePnt> 	 
     
    Pnt2D2(me)  
    	returns Pnt2d from gp; 
    ---C++: return const & 
    ---C++: inline  
    	---Purpose: 
    	--- Selector 
	--- Returns 2D point on the second face <thePnt>  
	
    SetIndex(me:out;  
    	    theIndex: Integer from Standard); 
    ---C++: inline      
     	---Purpose: 
    	--- Modifier
	--- Sets the index of the vertex <theIndex>
    Index(me)  
    	returns Integer from Standard; 
    ---C++: inline  
    	---Purpose: 
    	--- Selector 
	--- Returns index of the vertex   
	
fields
    myPnt :Pnt from gp is protected; 
    myPnt2D1:Pnt2d from gp is protected; 
    myPnt2D2:Pnt2d from gp is protected; 
    myIndex : Integer from Standard is protected;    

end Point;
