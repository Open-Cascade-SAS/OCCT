-- Created on: 2000-11-23
-- Created by: Michael KLOKOV
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class FaceFace from IntTools

    	---Purpose: This class provides the intersection of 
    	---	    face's underlying surfaces.

uses 

    TopolTool from Adaptor3d, 
    HSurface  from GeomAdaptor, 
    ListOfPntOn2S from IntSurf ,
    Intersection from IntPatch,
    Face from TopoDS,
    SequenceOfCurves from IntTools,
    LineConstructor from IntTools,
    SequenceOfPntOn2Faces from IntTools, 
    Context from BOPInt
    
    

raises NotDone from StdFail
is

    Create 
    	returns FaceFace from IntTools; 
    	---Purpose: 
    	--- Empty constructor.
	---


    SetParameters(me: in out;  
    	    	    ApproxCurves    : Boolean from Standard;
    	    	    ComputeCurveOnS1: Boolean from Standard;
    	    	    ComputeCurveOnS2: Boolean from Standard;
    	    	    ApproximationTolerance: Real from Standard);
    	---Purpose:
	--- Modifier
	---

    Perform(me: in out;  
    	    	    F1: Face from TopoDS;
    	    	    F2: Face from TopoDS);
    	---Purpose: 
    	--- Intersects underliing surfaces of F1 and F2
	--- Use sum of tolerance of F1 and F2 as intersection
	--- criteria
	---
	
    IsDone(me)
    	returns Boolean from Standard;
    	---Purpose: 
    	--- Returns True if the intersection was successful
	---

    Lines(me)
    	returns SequenceOfCurves from IntTools;
    	---C++: return const&	
    	---Purpose: 
    	--- Returns sequence of 3d curves as result of intersection
	---
	 
    Points(me)
    	returns  SequenceOfPntOn2Faces from IntTools;
    	---C++: return const&	 
    	---Purpose: 
    	--- Returns sequence of 3d curves as result of intersection
	---

    TolReached3d(me)  
    	returns Real from Standard;
	---Purpose:
	--- Returns tolerance reached during approximation.
	--- If approximation was not done, returns zero.
	---

    TolReached2d(me)  
    	returns Real from Standard;
	---Purpose:
    	--- Returns tolerance reached during approximation.
	--- If approximation was not done, returns zero.
	---
	     
    Face1  (me) 
    	returns  Face  from  TopoDS; 
	---C++: return const& 
	---Purpose:
	--- Returns first of processed faces
	---
	 
    Face2  (me) 
    	returns  Face  from  TopoDS; 
	---C++: return const& 
	---Purpose:
	--- Returns second of processed faces
	---
     
    TangentFaces  (me)
    	returns Boolean from Standard; 
	---Purpose:
	--- Returns True if faces are tangent
	--- 
    PrepareLines3D (me:out; 
    	    bToSplit: Boolean from Standard=Standard_True);
    	---Purpose: 
    	--- Provides post-processing the result lines. 
        --- <bToSplit> - the flag.    		     
    	--  In case of <bToSplit> is true the closed 3D-curves will be splitted  
        --  on parts. 
        --  In case of <bToSplit> is false the closed 3D-curves remain untouched.  
    
    SetList (me: in out;  
    	    ListOfPnts: in out ListOfPntOn2S from IntSurf);
    
    ----------------------------------------------------------
    --                  private  block
    ----------------------------------------------------------
    MakeCurve(me: in out; Index   : Integer from Standard;
    	                  D1      : TopolTool from Adaptor3d;
    	                  D2      : TopolTool from Adaptor3d)
	is protected; 
	
    ComputeTolReached3d(me:out) 
    	is  protected; 
 
    SetContext(me:out; 
    	  aContext : Context from BOPInt); 
     	---Purpose:
	--- Sets the intersecton context 
	
    Context(me) 
    	returns Context from BOPInt; 
    ---C++:  return const & 	
    	---Purpose:
	--- Gets the intersecton context	
	---	  
fields 
 
    myIsDone       : Boolean         from Standard;
    myIntersector  : Intersection    from IntPatch;
    myLConstruct   : LineConstructor from IntTools;
    myHS1          : HSurface        from GeomAdaptor;
    myHS2          : HSurface        from GeomAdaptor;
    myNbrestr      : Integer         from Standard;

    myTolReached2d : Real            from Standard;
    myTolReached3d : Real            from Standard;
    
    myApprox       : Boolean         from Standard;
    myApprox1      : Boolean         from Standard;
    myApprox2      : Boolean         from Standard;
    myTolApprox    : Real            from Standard;
    
    mySeqOfCurve : SequenceOfCurves from IntTools;

    myTangentFaces: Boolean         from Standard; 
    myFace1       : Face from TopoDS;  
    myFace2       : Face from TopoDS;  
    myPnts        : SequenceOfPntOn2Faces from IntTools;
    
    myListOfPnts  : ListOfPntOn2S from IntSurf;   
    
    myContext     : Context from  BOPInt;	 

end FaceFace from IntTools;

