-- Created on: 1999-08-04
-- Created by: Denis PASCAL
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class DriverTable from TPrsStd inherits TShared from MMgt

    ---Purpose:   This class is   a  container to record  (AddDriver)
    --          binding between  GUID and  TPrsStd_Driver. 
        -- You create a new instance of TPrsStd_Driver
-- and use the method AddDriver to load it into the driver table. the method
 

uses Boolean    from Standard,
     Attribute  from TDF,
     Label      from TDF,
     GUID       from Standard,
     IDList     from TDF,
     Driver     from TPrsStd,
     DataMapOfGUIDDriver from TPrsStd

is

    Get (myclass) returns mutable DriverTable from TPrsStd;
    ---Purpose: Returns the static table.
    --          If it does not exist, creates it and fills it with standard drivers.

    Create returns mutable DriverTable from TPrsStd;
    ---Purpose: Default constructor

    InitStandardDrivers (me : mutable);
    ---Purpose: Fills the table with standard drivers


    AddDriver (me : mutable; guid   : GUID   from Standard;
    	    	    	     driver : Driver from TPrsStd)
    ---Purpose: Returns true if the driver has been added successfully to the driver table.
    returns Boolean from Standard;

    FindDriver (me; guid   :     GUID   from Standard;
	 	    driver : out Driver from TPrsStd)
    ---Purpose: Returns true if the driver was found.
    returns Boolean from Standard;

    RemoveDriver (me : mutable; guid : GUID from Standard)
    ---Purpose:
-- Removes a driver with the given GUID.
  --      Returns true if the driver has been removed successfully.
    returns Boolean from Standard;

    Clear (me : mutable);
    ---Purpose: Removes all drivers. Returns
 -- true if the driver has been removed successfully.
 -- If this method is used, the InitStandardDrivers method should be
 -- called to fill the table with standard drivers.

fields

    myDrivers : DataMapOfGUIDDriver from TPrsStd;

end DriverTable;
