-- Created on: 1994-02-07
-- Created by: Modelistation
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package BRepIntCurveSurface 

	---Purpose: Inttantiates IntCurveSurface with Surfaces from BRep 
	--          and Curves from Adaptor

        ---Level: Public
        --
        -- All the methods of the classes of this package are public.
        -- 

uses  
--modified by NIZNHY-PKV Sun Dec 15 16:54:16 2002  f
    BRepTopAdaptor, 
--modified by NIZNHY-PKV Sun Dec 15 16:54:28 2002  t     
    IntCurveSurface, 
     BRepAdaptor,
     Geom2dInt,
     GeomAdaptor, 
     TopoDS,
     BRepClass, 
     TopAbs, 
     TopExp,
     StdFail,
     gp

is

    --------------------------------------------------
    -- Instantiation of IntCurveSurfaces algorithms --
    -- The intersection is computed on the surfaces --
    -- with their natural boundaries.               --
    --------------------------------------------------

--    class ICSSurfaceTool instantiates 
--          SurfaceTool from IntCurveSurface(
----	    HSurface     from BRepAdaptor) ;
--
----	    
--    class ICSCurveTool instantiates 
----    	  CurveTool from IntCurveSurface(
--	    HCurve       from GeomAdaptor) ;
----
--   
----    class ICSInter instantiates 
--          Inter from IntCurveSurface(
----	     HCurve           from GeomAdaptor,
-- 	     ICSCurveTool    from BRepIntCurveSurface,
----	     HSurface         from BRepAdaptor,
--             ICSSurfaceTool  from BRepIntCurveSurface);
--

    ------------------------------------------------------
    -- The Inter class provides intersection between    --
    --  - a BRepAdaptor surface and a GeomAdaptor curve --
    --  - a Shape               and a GeomAdaptor curve --
    -- Only the points which are inside the surface     --
    -- are returned.                                    --
    ------------------------------------------------------

    class Inter; 
    
    
    
    
end BRepIntCurveSurface;
