-- Created on: 2003-10-10
-- Created by: Alexander SOLOVYOV
-- Copyright (c) 2003-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


deferred class DataSource from MeshVS inherits TShared from MMgt

	---Purpose: The deferred class using for the following tasks:
	-- 1) Receiving geometry data about single element of node by its number;
	-- 2) Receiving type of element or node by its number;
 	-- 3) Receiving topological information about links between element and nodes it consist of;
        -- 4) Receiving information about what element cover this node;
        -- 5) Receiving information about all nodes and elements the object consist of 
	-- 6) Activation of advanced mesh selection. In the advanced mesh selection mode there is created: 
	--    - one owner for the whole mesh and for all selection modes
        --    - one sensitive entity for the whole mesh and for each selection mode	 
	--    Receiving of IDs of detected entities (nodes and elements) in a viewer is achieved by  
        --    implementation of a group of methods GetDetectedEntities. 
	 
uses
  Integer from Standard,
  Boolean from Standard,
  Address from Standard,

  Array1OfReal       from TColStd, 
  Array1OfInteger    from TColStd,
  PackedMapOfInteger from TColStd, 
  HPackedMapOfInteger from TColStd,
  HArray1OfReal      from TColStd, 
  Array1OfPnt2d      from TColgp,

  EntityType                 from MeshVS,
  HArray1OfSequenceOfInteger from MeshVS, 
   
  Box2d  from Bnd, 
  Box    from Bnd, 
   
  Mesh   from MeshVS  

is

  GetGeom ( me; ID     : Integer;
            IsElement  : Boolean;
            Coords     : out Array1OfReal from TColStd;
            NbNodes    : out Integer;
            Type       : out EntityType from MeshVS ) returns Boolean is deferred;
	---Purpose: Returns geometry information about node or element
        -- ID is the numerical identificator of node or element
        -- IsElement indicates this ID describe node ( if Standard_False ) or element ( if Standard_True )
        -- Coords is an array of co-ordinates of node(s).
        --     For node it is only 3 numbers: X, Y, Z in the strict order
        --     For element it is 3*n numbers, where n is number of this element vertices
        --     The order is strict also: X1, Y1, Z1, X2,...., where Xi, Yi, Zi are co-ordinates of vertices
        -- NbNodes is number of nodes. It is recommended this parameter to be set to 1 for node.
        -- Type is type of node or element (from enumeration). It is recommended this parameter to be set to
        --     MeshVS_ET_Node for node.

  GetGeomType ( me; ID     : Integer;
                IsElement  : Boolean;
                Type       : out EntityType from MeshVS ) returns Boolean is deferred;
	---Purpose: This method is similar to GetGeom, but returns only element or node type.
        --This method is provided for finer performance.

  Get3DGeom( me; ID      : Integer;
                 NbNodes : out Integer;
                 Data    : out HArray1OfSequenceOfInteger from MeshVS ) returns Boolean is virtual;
	---Purpose: This method returns topology information about 3D-element
        -- Returns false if element with ID isn't 3D or because other troubles


  GetAddr ( me; ID     : Integer;
            IsElement  : Boolean   ) returns Address is deferred;
	---Purpose: This method returns pointer which represents element or node data structure.
        -- This address will be saved in MeshVS_MeshEntityOwner, so that you can access to data structure fast
        -- by the method Owner(). In the redefined method you can return NULL.
        -- ID is the numerical identificator of node or element
        -- IsElement indicates this ID describe node ( if Standard_False ) or element ( if Standard_True )
 
  GetNodesByElement ( me; ID  : Integer;
		      NodeIDs : out Array1OfInteger from TColStd;
		      NbNodes : out Integer ) returns Boolean is deferred;
	---Purpose: This method returns information about nodes this element consist of.
        -- ID is the numerical identificator of element.
        -- NodeIDs is the output array of nodes IDs in correct order,
	-- the same as coordinates returned by GetGeom().
        -- NbNodes is number of nodes (number of items set in NodeIDs).
	-- Returns False if element does not exist

  GetAllNodes    ( me ) returns PackedMapOfInteger from TColStd is deferred;
	---C++: return const &
	---Purpose: This method returns map of all nodes the object consist of.

  GetAllElements ( me ) returns PackedMapOfInteger from TColStd is deferred;
	---C++: return const &
	---Purpose: This method returns map of all elements the object consist of.

  GetNormal ( me; Id : Integer; Max : Integer;
                  nx, ny, nz : out Real ) returns Boolean is virtual;
	---Purpose: This method calculates normal of face, which is using for correct reflection presentation.
        --   There is default method, for advance reflection this method can be redefined.
        -- Id is the numerical identificator of only element!
        -- Max is maximal number of nodes an element can consist of
        -- nx, ny, nz  are values whose represent co-ordinates of normal (will be returned)
        --   In the redefined method you can return normal with length more then 1, but in this case
        --   the appearance of element will be more bright than usual. For ordinary brightness you must return
        --   normal with length 1

  GetNodeNormal ( me; ranknode : Integer; ElementId : Integer;
                  nx, ny, nz : out Real ) returns Boolean is virtual;
	---Purpose: This method return normal of node ranknode of face Id, 
        --          which is using for smooth shading presentation.
        --          Returns false if normal isn't defined.

  GetNormalsByElement( me; Id       : Integer; 
                           IsNodal  : Boolean;
                           MaxNodes : Integer;
                           Normals  : out HArray1OfReal from TColStd ) returns Boolean is virtual;
	---Purpose: This method puts components of normal vectors at each node of a mesh face (at each face of a mesh volume)
    	-- into the output array.
    	-- Returns false if some problem was detected during calculation of normals.
    	-- Id is an identifier of the mesh element.
    	-- IsNodal, when true, means that normals at mesh element nodes are needed. If nodal normals
    	-- are not available, or IsNodal is false, or the mesh element is a volume, then the output array contents 
    	-- depend on the element type: 
    	--   face: a normal calculated by GetNormal() is duplicated for each node of the face;
    	--   volume: normals to all faces of the volume are computed (not for each node!).
    	-- MaxNodes is maximal number of nodes an element can consist of.
    	-- Normals contains the result.

  GetAllGroups ( me; Ids : out PackedMapOfInteger from TColStd ) is virtual;
	---Purpose: This method returns map of all groups the object contains.

  GetGroup ( me; Id : Integer; Type : out EntityType from MeshVS; 
                 Ids : out PackedMapOfInteger from TColStd ) returns Boolean is virtual;
	---Purpose: This method returns map of all group elements.

  GetGroupAddr ( me; ID : Integer ) returns Address is virtual;
	---Purpose: This method returns pointer which represents group data structure.
        -- This address will be saved in MeshVS_MeshOwner, so that you can access to data structure fast
        -- by the method Owner(). In the redefined method you can return NULL.
        -- ID is the numerical identificator of group

  IsAdvancedSelectionEnabled( me )
  returns Boolean from Standard is virtual;
    	---Purpose: Returns True if advanced mesh selection is enabled. 
        --          Default implementation returns False.  
	--          It should be redefined to return True for advanced
        --          mesh selection activation.

  GetBoundingBox( me ) returns Box from Bnd is virtual;
        ---Purpose: Returns the bounding box of the whole mesh.
        --          It is used in advanced selection mode to define roughly
        --          the sensitive area of the mesh.
        --          It can be redefined to get access to a box computed in advance.

  GetDetectedEntities( me : mutable;  Prs        : Mesh from MeshVS;    
    	    	    	              X,Y        : Real from Standard;
            	    	              aTol       : Real from Standard; 
			              Nodes      : out HPackedMapOfInteger from TColStd; 
    	    	    	              Elements   : out HPackedMapOfInteger from TColStd;
    	    	    	              DMin       : out Real from Standard )
  returns Boolean is virtual;
	---Purpose: Returns maps of entities (nodes and elements) detected
        --          by mouse click at the point (X,Y) on the current view plane, 
	--          with the tolerance aTol. 
	--          DMin - is out argument should return actual detection tolerance.
	--          Returns True if something is detected.
        --          It should be redefined if the advanced mesh selection is 
        --          activated. Default implementation returns False.
	 
  GetDetectedEntities( me : mutable;  Prs                     : Mesh from MeshVS; 
    	    	    	              XMin, YMin, XMax, YMax  : Real;
             	    	              aTol                    : Real; 
    	    	    	              Nodes                   : out HPackedMapOfInteger from TColStd;  
    	    	    	              Elements                : out HPackedMapOfInteger from TColStd )
  returns Boolean is virtual;
	---Purpose: Returns maps of entities (nodes and elements) detected 
	--          by mouse selection with rectangular box (XMin, YMin, XMax, YMax)
	--          on the current veiw plane, with the tolerance aTol. 
	--          Returns True if something is detected.
        --          It should be redefined if the advanced mesh selection is 
        --          activated. Default implementation returns False.
	 
  GetDetectedEntities( me : mutable;  Prs       : Mesh from MeshVS; 
    	    	    	              Polyline  : Array1OfPnt2d from TColgp;
                                      aBox      : Box2d; 
             	    	              aTol      : Real; 
			              Nodes     : out HPackedMapOfInteger from TColStd; 
    	    	    	              Elements  : out HPackedMapOfInteger from TColStd )
  returns Boolean is virtual;
	---Purpose: Returns maps of entities (nodes and elements) detected 
	--          by mouse selection with the polyline <Polyline> 
	--          on the current veiw plane, with the tolerance aTol. 
	--          Returns True if something is detected.
        --          It should be redefined if the advanced mesh selection is 
        --          activated. Default implementation returns False.

  GetDetectedEntities( me : mutable; Prs      : Mesh from MeshVS; 
                                     Nodes    : in out HPackedMapOfInteger from TColStd;
                                     Elements : in out HPackedMapOfInteger from TColStd )
  returns Boolean is virtual;
	---Purpose: Filter out the maps of mesh entities so as to keep
	--          only the entities that are allowed to be selected
	--          according to the current context.
	--          Returns True if any of the maps has been changed.
        --          It should be redefined if the advanced mesh selection is 
        --          activated. Default implementation returns False.
				   
end DataSource;
