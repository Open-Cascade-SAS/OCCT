-- Created on: 1994-08-03
-- Created by: Modeling
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package MeshTest 

	---Purpose: Provides methods for testing the mesh algorithms.

uses 
     TColStd,
     Draw,
     TopoDS,
     BRepMesh

is

    imported DrawableMesh from MeshTest;

    Commands(DI : in out Interpretor from Draw);
	---Purpose: Defines meshing commands 

    PluginCommands(DI : in out Interpretor from Draw);
    	---Purpose: Defines plugin commands 

end MeshTest;
