-- File:	IGESType.cdl
-- Created:	Mon Apr  6 14:24:36 1992
-- Author:	Christian CAILLET
--		<cky@phobox>
---Copyright:	 Matra Datavision 1992


class IGESType  from IGESData

    ---Purpose : taken from directory part of an entity (from file or model),
    --           gives "type" and "form" data, used to recognize entity's type

uses Integer

is

    Create returns IGESType;  -- default constructor (gives type = form = 0)

    Create (atype, aform : Integer) returns IGESType;

    Type (me) returns Integer  is static;
    ---Purpose : returns "type" data

    Form (me) returns Integer  is static;
    ---Purpose : returns "form" data

    IsEqual (me; another : IGESType) returns Boolean  is static;
    ---Purpose : compares two IGESTypes, avoiding comparing their fields
    ---C++ : alias operator ==

    Nullify (me : in out)  is static;
    ---Purpose : resets fields (usefull when an IGESType is stored as mask)

fields

    thetype : Integer;
    theform : Integer;

end IGESType;
