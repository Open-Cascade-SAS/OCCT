-- Created on: 2002-12-12
-- Created by: data exchange team
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class UniformSurfaceSection from StepElement
inherits SurfaceSection from StepElement

    ---Purpose: Representation of STEP entity UniformSurfaceSection

uses
    MeasureOrUnspecifiedValue from StepElement

is
    Create returns UniformSurfaceSection from StepElement;
	---Purpose: Empty constructor

    Init (me: mutable; aSurfaceSection_Offset: MeasureOrUnspecifiedValue from StepElement;
                       aSurfaceSection_NonStructuralMass: MeasureOrUnspecifiedValue from StepElement;
                       aSurfaceSection_NonStructuralMassOffset: MeasureOrUnspecifiedValue from StepElement;
                       aThickness: Real;
                       aBendingThickness: MeasureOrUnspecifiedValue from StepElement;
                       aShearThickness: MeasureOrUnspecifiedValue from StepElement);
	---Purpose: Initialize all fields (own and inherited)

    Thickness (me) returns Real;
	---Purpose: Returns field Thickness
    SetThickness (me: mutable; Thickness: Real);
	---Purpose: Set field Thickness

    BendingThickness (me) returns MeasureOrUnspecifiedValue from StepElement;
	---Purpose: Returns field BendingThickness
    SetBendingThickness (me: mutable; BendingThickness: MeasureOrUnspecifiedValue from StepElement);
	---Purpose: Set field BendingThickness

    ShearThickness (me) returns MeasureOrUnspecifiedValue from StepElement;
	---Purpose: Returns field ShearThickness
    SetShearThickness (me: mutable; ShearThickness: MeasureOrUnspecifiedValue from StepElement);
	---Purpose: Set field ShearThickness

fields
    theThickness: Real;
    theBendingThickness: MeasureOrUnspecifiedValue from StepElement;
    theShearThickness: MeasureOrUnspecifiedValue from StepElement;

end UniformSurfaceSection;
