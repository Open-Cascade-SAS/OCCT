-- Created on: 1992-09-22
-- Created by: Christian CAILLET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



package IFGraph

    	---Purpose : Provides tools to operate on an InterfaceModel and its
    	--           Entities as on a Graph. These Tools are based on classes
    	--           Graph and GraphContent  from Interface

uses Interface, GraphTools, TColStd, Standard

is

--  (sub-classes of GraphContent from Interface)
    	class AllShared;
	class AllConnected;
    	class Cumulate;
    	class Compare;
	class ExternalSources;

    	class Articulations;

    class SubPartsIterator;  -- result as several subsets
    	class ConnectedComponants;
    	class StrongComponants;
	class Cycles;
	class SCRoots;

--    class SortedStrongsFrom  instantiates  SortedStrgCmptsFromIterator from GraphTools
--    	(Graph from Interface,Transient,
--    	 MapTransientHasher from TColStd,GraphContent from Interface);

--    class SortedStrongs instantiates SortedStrgCmptsIterator from GraphTools
--    	(Graph from Interface,Transient,
--    	 GraphContent from Interface,SortedStrongsFrom from IFGraph);

--    class SortedStrongs instantiates SortedStrgCmptsIterator
--    	(Graph,Transient,GraphContent,GraphContent);

end IFGraph;
