-- Created on: 1999-02-24
-- Created by: Christian CAILLET
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class RemoveCurves  from IGESSelect    inherits ModelModifier from IGESSelect

    ---Purpose : Removes Curves UV or 3D (not both !) from Faces, those
    --           designated by the Selection. No Selection means all the file

uses AsciiString from TCollection,
     IGESModel, CopyTool, ContextModif
 
is

    Create (UV : Boolean) returns mutable RemoveCurves;
    ---Purpose : Creates a RemoveCurves from Faces (141/142/143/144)
    --           UV True  : Removes UV Curves (pcurves)
    --           UV False : Removes 3D Curves

    Performing (me; ctx : in out ContextModif;
                target  : mutable IGESModel;
                TC      : in out CopyTool);
    ---Purpose : Specific action : Removes the Curves
 
    Label (me) returns AsciiString from TCollection;
    ---Purpose : Returns a text which is
    --           "Remove Curves UV on Face"  or  "Remove Curves 3D on Face"

fields

    theUV : Boolean;

end RemoveCurves;
