-- Created on: 2000-05-24
-- Created by: Edward AGAPOV
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DocumentStorageDriver from XCAFDrivers 
inherits DocumentStorageDriver from MDocStd
		    
	---Purpose: storage driver of a  XS document
		    
uses
    ASDriverTable from MDF,
    MessageDriver from CDM

is
    Create returns mutable DocumentStorageDriver from XCAFDrivers;

    AttributeDrivers(me : mutable; theMessageDriver : MessageDriver from CDM)
    returns ASDriverTable from MDF
    is redefined;

end DocumentStorageDriver;
    
