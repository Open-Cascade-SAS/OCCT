-- Created on: 1999-11-09
-- Created by: data exchange team
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package RWStepAP203 

    ---Purpose: Reading & Writing tools for classes from StepAP203

uses
    Interface,
    StepData,
    StepAP203

is

    class RWCcDesignApproval;
    class RWCcDesignCertification;
    class RWCcDesignContract;
    class RWCcDesignDateAndTimeAssignment;
    class RWCcDesignPersonAndOrganizationAssignment;
    class RWCcDesignSecurityClassification;
    class RWCcDesignSpecificationReference;
    class RWChange;
    class RWChangeRequest;
    class RWStartRequest;
    class RWStartWork;

end RWStepAP203;
