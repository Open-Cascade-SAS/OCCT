-- Created on: 1991-10-04
-- Created by: Remi GILET
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class BPoint from GccInt  

inherits Bisec from GccInt 
     ---Purpose: Describes a point as a bisecting object between two 2D geometric objects.
        
uses Pnt2d from gp,
     IType  from GccInt


is

Create(Point : Pnt2d) returns BPoint;
    ---Purpose: Constructs a bisecting object whose geometry is the 2D point Point.
    
Point(me) returns Pnt2d from gp
    is redefined;
    ---Purpose: Returns a 2D point which is the geometry of this bisecting object.
    
ArcType(me) returns IType from GccInt
    is static;
    --- Purpose: Returns GccInt_Pnt, which is the type of any GccInt_BPoint bisecting object.
    
fields

    pnt : Pnt2d from gp;
    ---Purpose: The bisecting line.

end BPoint;    

