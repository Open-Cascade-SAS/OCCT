-- File:	IntImp_ZerCOnSSParFunc.cdl
-- Created:	Mon Feb 14 12:15:50 1994
-- Author:	Jacques GOUSSARD
--		<jag@topsn2>
---Copyright:	 Matra Datavision 1994


generic class ZerCOnSSParFunc from IntImp 
    (ThePSurface     as any;
     ThePSurfaceTool as any;   --as PSurfaceTool from IntImp(ThePSurface)
     TheCurveOnSurf  as any;
     TheCurveTool    as any     --as COnSCurveTool from IntImp(TheCurve)
    )
    
inherits FunctionSetWithDerivatives from math

      	---Purpose: this function is associated to the intersection between 
      	--          a curve on surface and a surface  .


uses Vector from math,
     Matrix from math,
     Pnt from gp

is
    Create( S1 : ThePSurface;
    	    C  : TheCurveOnSurf;
            S2 : ThePSurface )

	---Purpose: S1 is the surface on which the intersection is searched.
	--          C is a curve on the surface S2.

    	returns ZerCOnSSParFunc from IntImp;
	    

    NbVariables(me) returns Integer from Standard
    is static;
    
    NbEquations(me) returns Integer from Standard
    is static;
    
    Value(me : in out; X : in Vector from math;
    	    	       F : out Vector from math)
    returns Boolean from Standard
    is static;
    
    Derivatives(me : in out;X : in  Vector from math;
    	    	    	    D : out Matrix from math)
    returns Boolean from Standard
    is static;
    
    Values(me : in out;
    	   X  : in Vector from math;
	   F  : out Vector from math; D: out Matrix from math)
    returns Boolean from Standard
    is static;

    Point(me)
    	---C++: return const&
    	returns Pnt from gp
    	is static;
    
    Root(me) returns Real from Standard
    is static;
    
    AuxillarSurface(me)
    	---C++: return const&
    	returns ThePSurface
    	is static;

    AuxillarCurve(me)
    	---C++: return const&
    	returns TheCurveOnSurf
    	is static;
    
fields
     curve    : Address from Standard; --- TheCurveOnSurf;
     surface1 : Address from Standard; --- ThePSurface;
     surface2 : Address from Standard; --- ThePSurface;
     p	      : Pnt from gp;
     f        : Real from Standard;
     
end ZerCOnSSParFunc;
