-- File:	DefSwitch.cdl
-- Created:	Mon Apr  6 14:40:25 1992
-- Author:	Christian CAILLET
--		<cky@phobox>
---Copyright:	 Matra Datavision 1992


class DefSwitch  from IGESData  inherits Storable

    ---Purpose : description of a directory componant which can be either
    --           undefined (let Void), defined as a Reference to an entity,
    --           or as a Rank, integer value adressing a builtin table
    --           The entity reference is not included here, only reference
    --           status is kept (because entity type must be adapted)

uses Integer, DefType

is

    Create returns DefSwitch;
    ---Purpose : creates a DefSwitch as Void

    SetVoid (me : in out)  is static;
    ---Purpose : sets DefSwitch to "Void" status (in file : Integer = 0)

    SetReference (me : in out)  is static;
    ---Purpose : sets DefSwitch to "Reference" Status (in file : Integer < 0)

    SetRank (me : in out; val : Integer)  is static;
    ---Purpose : sets DefSwitch to "Rank" with a Value (in file : Integer > 0)

    DefType (me) returns DefType  is static;
    ---Purpose : returns DefType status (Void,Reference,Rank)

    Value (me) returns Integer  is static;
    ---Purpose : returns Value as Integer (sensefull for a Rank)

fields

    theval : Integer;

end DefSwitch;
