-- File:        StyledItem.cdl
-- Created:     Mon Dec  4 12:02:31 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWStyledItem from RWStepVisual

	---Purpose : Read & Write Module for StyledItem

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     StyledItem from StepVisual,
     EntityIterator from Interface

is

	Create returns RWStyledItem;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable StyledItem from StepVisual);

	WriteStep (me; SW : in out StepWriter; ent : StyledItem from StepVisual);

	Share(me; ent : StyledItem from StepVisual; iter : in out EntityIterator);

end RWStyledItem;
