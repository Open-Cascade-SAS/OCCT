-- Created by: Tanya COOL
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Radius from Prs2d inherits Dimension from Prs2d

 ---Purpose: Constructs the primitive Radius

uses

	Drawer	           from Graphic2d,
	GraphicObject      from Graphic2d,
	Pnt2d              from gp,
	Circ2d             from gp,
	ExtendedString     from TCollection,
	ArrowSide          from Prs2d,
	TypeOfDist         from Prs2d,
	TypeOfArrow        from Prs2d,
    	FStream            from Aspect 

raises 

  ConstructionError from Standard

is
	Create( aGraphicObject: GraphicObject  from Graphic2d;
	        anAttachPnt   : Pnt2d          from gp;
		aCircle       : Circ2d         from gp;
            	aText         : ExtendedString from TCollection;
		aTxtScale     : Real           from Standard = 10.0; 
		anArrAngle    : Real           from Standard = 20.0;
		anArrLength   : Real           from Standard = 25.0;
            	anArrType     : TypeOfArrow    from Prs2d    = Prs2d_TOA_OPENED;
		anArrow       : ArrowSide      from Prs2d    = Prs2d_AS_BOTHAR;
		IsReverseArrow: Boolean        from Standard = Standard_False )
	returns mutable Radius from Prs2d;

    ---Purpose: Creates the radius of the circle passing through 
    --          the point <anAttachPnt>

    	--------------------------------------
	-- Category: Inquire methods
	--------------------------------------
    
    Values( me; anAttPnt: out Pnt2d from gp; 
            aCirc: out Circ2d from gp ); 
    ---Level: Internal
    ---Purpose: allows to get the properties of the diameter

	--------------------------
	-- Category: Draw and Pick
	--------------------------

    Draw( me : mutable; aDrawer: Drawer from Graphic2d )
	is static protected;
    ---Level: Internal
    ---Purpose: Draws the angle <me>.

    DrawElement( me : mutable; aDrawer: Drawer from Graphic2d;
                 anIndex: Integer from Standard)
        is redefined protected;
    ---Level: Internal
    ---Purpose: Draws element <anIndex> of the radius <me>.

    DrawVertex( me : mutable; aDrawer: Drawer from Graphic2d;
                anIndex: Integer from Standard)
        is redefined protected;
    ---Level: Internal
    ---Purpose: Draws vertex <anIndex> of the radius <me>.

    Pick( me : mutable; X, Y: ShortReal from Standard;
      	  aPrecision: ShortReal from Standard;
       	  aDrawer: Drawer from Graphic2d)
	returns Boolean from Standard
	is static protected;
    ---Level: Internal
    ---Purpose: Returns Standard_True if the radius <me> is picked,
    --	    Standard_False if not.

	Save( me; aFStream: in out FStream from Aspect ) is virtual;
	
	CalcTxtPos(me:mutable; theFromAbs: 
    	    	    Boolean from Standard=Standard_False) 
    	---C++: inline 
    	is redefined protected;
				 										
fields
 
	myX1   : ShortReal  from Standard;
	myY1   : ShortReal  from Standard;
	myX2   : ShortReal  from Standard;
	myY2   : ShortReal  from Standard;
    	myPnt  : Pnt2d      from gp;
    	myCirc : Circ2d     from gp;
    	
end Radius from Prs2d;
