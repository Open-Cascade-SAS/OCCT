-- Created on: 1992-06-22
-- Created by: Gilles DEBARBOUILLE
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



private class Sentence from Units 

	---Purpose: This class describes all the methods to create and
	--          compute an expression contained in a string.

uses

    Token          from Units,
    TokensSequence from Units,
    Lexicon        from Units

--raises

is

    Create(alexicon : Lexicon from Units ; astring : CString)
    
    ---Level: Internal 
    
    ---Purpose: Creates and  returns  a   Sentence, by  analyzing  the
    --          string <astring> with the lexicon <alexicon>.
    
    returns Sentence from Units;
    
    SetConstants(me : in out)
    
    ---Level: Internal 
    
    ---Purpose: For each constant encountered, sets the value.
    
    is static;
    
    Sequence(me) returns any TokensSequence from Units
    
    ---Level: Internal 
    
    ---C++: inline
    
    ---Purpose: Returns <thesequenceoftokens>.
    
    is static;
    
    Sequence(me : in out ; asequenceoftokens : any TokensSequence from Units)
    
    ---Level: Internal 
    
    ---C++: inline
    
    ---Purpose: Sets the field <thesequenceoftokens> to <asequenceoftokens>.
    
    is static;
    
    Evaluate(me : in out)returns mutable Token from Units
    
    ---Level: Internal 
    
    ---Purpose: Computes and  returns in a   token the result  of  the
    --          expression.
    
    is static;
    
    IsDone(me) returns Boolean from Standard
    ---Level: Internal 
    ---C++: inline
    ---Purpose: Return True if number of created tokens > 0
    --          (i.e creation of sentence is succesfull)
    is static;

    Dump(me)
    
    ---Level: Internal 
    
    ---C++: inline
    
    ---Purpose: Useful for debugging.
    
    is static;

fields

    thesequenceoftokens : TokensSequence from Units;

end Sentence;
