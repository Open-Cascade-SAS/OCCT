-- File:	RWStepFEA_RWArbitraryVolume3dElementCoordinateSystem.cdl
-- Created:	Thu Dec 12 17:51:03 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWArbitraryVolume3dElementCoordinateSystem from RWStepFEA

    ---Purpose: Read & Write tool for ArbitraryVolume3dElementCoordinateSystem

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    ArbitraryVolume3dElementCoordinateSystem from StepFEA

is
    Create returns RWArbitraryVolume3dElementCoordinateSystem from RWStepFEA;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : ArbitraryVolume3dElementCoordinateSystem from StepFEA);
	---Purpose: Reads ArbitraryVolume3dElementCoordinateSystem

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: ArbitraryVolume3dElementCoordinateSystem from StepFEA);
	---Purpose: Writes ArbitraryVolume3dElementCoordinateSystem

    Share (me; ent : ArbitraryVolume3dElementCoordinateSystem from StepFEA;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWArbitraryVolume3dElementCoordinateSystem;
