-- Created on: 1991-01-14
-- Created by: Arnaud BOUZY
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class RelationIterator from Expr

	---Purpose: Iterates on every basic relation contained in
	--          a GeneralRelation.
        ---Level : Internal

uses GeneralRelation from Expr,
    SingleRelation from Expr,
    Array1OfSingleRelation from Expr

raises NoMoreObject from Standard,
    NoSuchObject from Standard

is

    Create(rel : GeneralRelation)
    returns RelationIterator;
    
    More(me)
    ---Purpose: Returns False if no other relation remains.
    returns Boolean
    is static;
    
    Next(me : in out)
    raises NoMoreObject
    is static;
    
    Value(me)
    ---Purpose: Returns current basic relation.
    --          Exception is raised if no more relation remains.
    returns  SingleRelation
    raises NoSuchObject
    is static;

fields

    myRelation : Array1OfSingleRelation;
    current : Integer;

end RelationIterator;
