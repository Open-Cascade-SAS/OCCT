-- File:        BackgroundColour.cdl
-- Created:     Fri Dec  1 11:11:15 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class BackgroundColour from StepVisual 

inherits Colour from StepVisual 

uses

	AreaOrView from StepVisual
is

	Create returns mutable BackgroundColour;
	---Purpose: Returns a BackgroundColour

	Init (me : mutable;
	      aPresentation : AreaOrView from StepVisual) is virtual;

	-- Specific Methods for Field Data Access --

	SetPresentation(me : mutable; aPresentation : AreaOrView);
	Presentation (me) returns AreaOrView;

fields

	presentation : AreaOrView from StepVisual; -- a SelectType

end BackgroundColour;
