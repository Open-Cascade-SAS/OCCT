-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class ReversibleTopologyItem from StepShape inherits SelectType from StepData

	-- <ReversibleTopologyItem> is an EXPRESS Select Type construct translation.
	-- it gathers : Edge, Path, Face, FaceBound, ClosedShell, OpenShell

uses

	Edge,
	Path,
	Face,
	FaceBound,
	ClosedShell,
	OpenShell
is

	Create returns ReversibleTopologyItem;
	---Purpose : Returns a ReversibleTopologyItem SelectType

	CaseNum (me; ent : Transient) returns Integer;
	---Purpose: Recognizes a ReversibleTopologyItem Kind Entity that is :
	--        1 -> Edge
	--        2 -> Path
	--        3 -> Face
	--        4 -> FaceBound
	--        5 -> ClosedShell
	--        6 -> OpenShell
	--        0 else

	Edge (me) returns any Edge;
	---Purpose : returns Value as a Edge (Null if another type)

	Path (me) returns any Path;
	---Purpose : returns Value as a Path (Null if another type)

	Face (me) returns any Face;
	---Purpose : returns Value as a Face (Null if another type)

	FaceBound (me) returns any FaceBound;
	---Purpose : returns Value as a FaceBound (Null if another type)

	ClosedShell (me) returns any ClosedShell;
	---Purpose : returns Value as a ClosedShell (Null if another type)

	OpenShell (me) returns any OpenShell;
	---Purpose : returns Value as a OpenShell (Null if another type)


end ReversibleTopologyItem;

