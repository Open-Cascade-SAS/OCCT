-- File:	StepToTopoDS_Builder.cdl
-- Created:	Fri Dec 16 14:49:51 1994
-- Author:	Frederic MAUPAS
--		<fma@stylox>
---Copyright:	 Matra Datavision 1994

class Builder from StepToTopoDS
    inherits Root from StepToTopoDS
    
    ---Purpose:
    --         


uses

    ManifoldSolidBrep           from StepShape,
    BrepWithVoids               from StepShape,
    FacetedBrep                 from StepShape,
    FacetedBrepAndBrepWithVoids from StepShape,
    ShellBasedSurfaceModel      from StepShape,
    EdgeBasedWireframeModel     from StepShape,
    FaceBasedSurfaceModel       from StepShape,
    GeometricSet                from StepShape,
    Shape                       from TopoDS,
    BuilderError                from StepToTopoDS,
    TransientProcess            from Transfer,
    NMTool                      from StepToTopoDS
    
    raises NotDone from StdFail
     
is 

    Create returns Builder from StepToTopoDS;
    
    Create (S  : ManifoldSolidBrep from StepShape;
       	    TP : TransientProcess  from Transfer )
	returns Builder from StepToTopoDS;
     
    Create (S  : BrepWithVoids from StepShape;
            TP : TransientProcess  from Transfer )
    	returns Builder from StepToTopoDS;

    Create ( S : FacetedBrep from StepShape;
            TP : TransientProcess  from Transfer )
    	returns Builder from StepToTopoDS;

    Create (S  : FacetedBrepAndBrepWithVoids from StepShape;
            TP : TransientProcess  from Transfer )
    	returns Builder from StepToTopoDS;

    Create (S      : ShellBasedSurfaceModel from StepShape;
            TP     : TransientProcess  from Transfer;
            NMTool : in out NMTool from StepToTopoDS )
    	returns Builder from StepToTopoDS;

    Create ( S : GeometricSet from StepShape;
            TP : TransientProcess  from Transfer )
    	returns Builder from StepToTopoDS;

    Init (me : in out;
    	  S  : ManifoldSolidBrep from StepShape;
          TP : TransientProcess  from Transfer );

    Init (me : in out;
    	  S  : BrepWithVoids from StepShape;
          TP : TransientProcess  from Transfer );

    Init (me : in out;
    	  S  : FacetedBrep from StepShape;
          TP : TransientProcess  from Transfer );

    Init (me : in out;
    	  S  : FacetedBrepAndBrepWithVoids from StepShape;
          TP : TransientProcess  from Transfer );
	  
    Init (me     : in out;
    	   S     : ShellBasedSurfaceModel from StepShape;
          TP     : TransientProcess  from Transfer;
	  NMTool : in out NMTool from StepToTopoDS );
	  
    Init (me : in out;
    	  S  : EdgeBasedWireframeModel from StepShape;
          TP : TransientProcess  from Transfer );
	  
    Init (me : in out;
    	  S  : FaceBasedSurfaceModel from StepShape;
          TP : TransientProcess  from Transfer );
	  
    Init (me : in out;
    	  S  : GeometricSet from StepShape;
          TP : TransientProcess  from Transfer );
	  
    Value (me) returns Shape from TopoDS
    	raises NotDone
    	is static;
    	---C++: return const&
    
    Error (me) returns BuilderError from StepToTopoDS
    	is static;

fields

    myError  : BuilderError from StepToTopoDS;    
    
    myResult : Shape from TopoDS;
    
end Builder;
