-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class FillStyleSelect from StepVisual inherits SelectType from StepData

	-- <FillStyleSelect> is an EXPRESS Select Type construct translation.
	-- it gathers : FillAreaStyleColour, ExternallyDefinedTileStyle, FillAreaStyleTiles, ExternallyDefinedHatchStyle, FillAreaStyleHatching
	-- Rev4 : only FillAreaStyleColour remains

uses

	FillAreaStyleColour
--	ExternallyDefinedTileStyle,
--	FillAreaStyleTiles,
--	ExternallyDefinedHatchStyle,
--	FillAreaStyleHatching
is

	Create returns FillStyleSelect;
	---Purpose : Returns a FillStyleSelect SelectType

	CaseNum (me; ent : Transient) returns Integer;
	---Purpose: Recognizes a FillStyleSelect Kind Entity that is :
	--        1 -> FillAreaStyleColour
	--        2 -> ExternallyDefinedTileStyle
	--        3 -> FillAreaStyleTiles
	--        4 -> ExternallyDefinedHatchStyle
	--        5 -> FillAreaStyleHatching
	--        0 else

	FillAreaStyleColour (me) returns any FillAreaStyleColour;
	---Purpose : returns Value as a FillAreaStyleColour (Null if another type)


end FillStyleSelect;

