-- Created on: 1993-01-09
-- Created by: CKY / Contract Toubro-Larsen ( TCD )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class LabelDisplay from IGESDraw  inherits LabelDisplayEntity

        ---Purpose: defines IGESLabelDisplay, Type <402> Form <5>
        --          in package IGESDraw
        --
        --          Permits one or more displays for the
        --          entity labels of an entity

uses

        IGESEntity              from IGESData,
        HArray1OfIGESEntity     from IGESData,
        LeaderArrow             from IGESDimen,
        HArray1OfLeaderArrow    from IGESDimen,
        HArray1OfInteger        from TColStd,
        ViewKindEntity          from IGESData,
        HArray1OfViewKindEntity from IGESDraw,
        Pnt                     from gp,
        HArray1OfXYZ            from TColgp

raises DimensionMismatch, OutOfRange

is

        Create returns LabelDisplay;

        -- Specific Methods pertaining to the class

        Init (me                   : mutable;
              allViews             : HArray1OfViewKindEntity;
              allTextLocations     : HArray1OfXYZ;
              allLeaderEntities    : HArray1OfLeaderArrow;
              allLabelLevels       : HArray1OfInteger;
              allDisplayedEntities : HArray1OfIGESEntity)
        raises DimensionMismatch;
        ---Purpose : This method is used to set the fields of the class
        --           LabelDisplay
        --   - allViews             : Pointers to View Entities
        --   - allTextLocations     : Coordinates of text locations in the views
        --   - allLeaderEntities    : Pointers to Leader Entities in the views
        --   - allLabelLevels       : Entity label level numbers in the views
        --   - allDisplayedEntities : Pointers to the entities being displayed
        -- raises exception if Lengths of allViews, allTextLocations,
        -- allLeaderEntities, allLabelLevels and allDisplayedEntities are
        -- not same.

        NbLabels (me) returns Integer;
        ---Purpose : returns the number of label placements in <me>

        ViewItem (me; ViewIndex : Integer) returns ViewKindEntity
        raises OutOfRange;
        ---Purpose : returns the View entity indicated by ViewIndex
        -- raises an exception if ViewIndex <= 0 or ViewIndex > NbLabels().

        TextLocation (me; ViewIndex : Integer) returns Pnt
        raises OutOfRange;
        ---Purpose : returns the 3d-Point coordinates of the text location, in the
        -- view indicated by ViewIndex
        -- raises an exception if ViewIndex <= 0 or ViewIndex > NbLabels().

        LeaderEntity (me; ViewIndex : Integer) returns LeaderArrow
        raises OutOfRange;
        ---Purpose : returns the Leader entity in the view indicated by ViewIndex
        -- raises an exception if ViewIndex <= 0 or ViewIndex > NbLabels().

        LabelLevel (me; ViewIndex : Integer) returns Integer
        raises OutOfRange;
        ---Purpose : returns the Entity label level number in the view indicated
        -- by ViewIndex
        -- raises an exception if ViewIndex <= 0 or ViewIndex > NbLabels().

        DisplayedEntity (me; EntityIndex : Integer) returns IGESEntity
        raises OutOfRange;
        ---Purpose : returns the entity indicated by EntityIndex
        -- raises an exception if EntityIndex <= 0 or EntityIndex > NbLabels().

        TransformedTextLocation (me; ViewIndex : Integer) returns Pnt
        raises OutOfRange;
        ---Purpose : returns the transformed 3d-Point coordinates of the text
        -- location, in the view indicated by ViewIndex
        -- raises an exception if ViewIndex <= 0 or ViewIndex > NbLabels().

fields

--
-- Class    : IGESDraw_LabelDisplay
--
-- Purpose  : Declaration of the variables specific to a Label Display.
--
-- Reminder : A Label Display is defined by :
--                    - Pointers to View Entities
--                    - Coordinates of text locations in the views
--                    - Pointers to Leader Entities in the views
--                    - Entity label level numbers in the views
--                    - Pointers to the entities being displayed
--

        theViews             : HArray1OfViewKindEntity;

        theTextLocations     : HArray1OfXYZ;

        theLeaderEntities    : HArray1OfLeaderArrow;

        theLabelLevels       : HArray1OfInteger;

        theDisplayedEntities : HArray1OfIGESEntity;

end LabelDisplay;
