-- Created on: 2000-07-03
-- Created by: Andrey BETENEV
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1

class RWSpecifiedHigherUsageOccurrence from RWStepRepr

    ---Purpose: Read & Write tool for SpecifiedHigherUsageOccurrence

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    SpecifiedHigherUsageOccurrence from StepRepr

is
    Create returns RWSpecifiedHigherUsageOccurrence from RWStepRepr;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : SpecifiedHigherUsageOccurrence from StepRepr);
	---Purpose: Reads SpecifiedHigherUsageOccurrence

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: SpecifiedHigherUsageOccurrence from StepRepr);
	---Purpose: Writes SpecifiedHigherUsageOccurrence

    Share (me; ent : SpecifiedHigherUsageOccurrence from StepRepr;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWSpecifiedHigherUsageOccurrence;
