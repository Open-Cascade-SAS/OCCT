-- Created on: 1994-03-30
-- Created by: Laurent BUCHARD
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.





class SolidClassifier from BRepClass3d  inherits SClassifier from BRepClass3d
     
     ---Purpose: Provides an algorithm to classify a point in a solid.



uses 
    Pnt           from gp,
    Face          from TopoDS,
    Shape         from TopoDS,
    SolidExplorer from BRepClass3d

raises

    DomainError from Standard
	
is 


    Create
    	---Purpose : empty constructor
    returns SolidClassifier from BRepClass3d;
        
    Load(me:in out; S   :        Shape from TopoDS)
    is static;
    

    Create(S   :        Shape from TopoDS)
    	---Purpose: Constructor from a Shape.
    returns SolidClassifier from BRepClass3d;
    
    
    Create(S   :        Shape from TopoDS; 
           P   :        Pnt from gp;
	   Tol :        Real from Standard)
    	---Purpose: Constructor to classify the point P with the 
    	--          tolerance Tol on the solid S.
    returns SolidClassifier from BRepClass3d;
    

    Perform(me: in out;
            P   :        Pnt from gp;
	    Tol :        Real from Standard)
    	---Purpose: Classify the point P with the 
    	--          tolerance Tol on the solid S.
    is static;

    PerformInfinitePoint(me: in out;
			 Tol :        Real from Standard)
    	---Purpose: Classify an infinite point with the 
    	--          tolerance Tol on the solid S.
    	--          Useful for compute the orientation of a solid. 
    is static;
    
    Destroy(me:in out)
    	---C++: alias ~
    is static;
    

fields
    aSolidLoaded   : Boolean       from Standard;
    explorer       : SolidExplorer from BRepClass3d;
    isaholeinspace : Boolean       from Standard;
end SolidClassifier;
