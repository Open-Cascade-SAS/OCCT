-- Created on: 1997-01-20
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package TestTopOpeDraw

uses 

    TopoDS,
    Draw,
    DrawTrSurf,
    DBRep,
    TCollection,
    Geom2d,
    Geom,
    gp,
    TestTopOpeTools,
    Standard,
    TColgp
        
is
    
    class ListOfPnt2d instantiates List from TCollection(Pnt2d from gp);
    class DrawableSHA;
    class DrawableSUR;
    class DrawableC3D;
    class DrawableC2D;
    class DrawableP3D;
    class Array1OfDrawableP3D instantiates Array1 from TCollection
    (DrawableP3D from TestTopOpeDraw);
    class HArray1OfDrawableP3D instantiates HArray1 from TCollection
    (DrawableP3D from TestTopOpeDraw,Array1OfDrawableP3D from TestTopOpeDraw);
    class DrawableP2D;

    class DrawableMesure;
    class Array1OfDrawableMesure instantiates Array1 from TCollection
    (DrawableMesure from TestTopOpeDraw);
    class HArray1OfDrawableMesure instantiates HArray1 from TCollection
    (DrawableMesure from TestTopOpeDraw,
     Array1OfDrawableMesure from TestTopOpeDraw);

    AllCommands(I : in out Interpretor from Draw);
    OtherCommands(I : in out Interpretor from Draw);

end TestTopOpeDraw;
