-- File:      Intf_InterferencePolygon2d.cdl
-- Created:   Mon Sep 28 17:09:45 1992
-- Author:    Didier PIFFAULT
---Copyright: Matra Datavision 1992


class InterferencePolygon2d from Intf

inherits Interference from Intf

	---Purpose: Computes the  interference between two  polygons or
	--          the    self intersection of    a  polygon  in  two
	--          dimensions.

uses    Pnt2d             from gp,
    	SectionPoint      from Intf,
    	SeqOfSectionPoint from Intf,
    	TangentZone       from Intf,
    	SeqOfTangentZone  from Intf,
        Polygon2d         from Intf

raises  OutOfRange from Standard

is

-- Interface :

    Create          returns InterferencePolygon2d from Intf;
    ---Purpose: Constructs an empty interference of Polygon.


    Create         (Obje1, Obje2 : in Polygon2d) 
    	            returns InterferencePolygon2d from Intf;
    ---Purpose: Constructs and computes an interference between two Polygons.


    Create         (Obje       : in Polygon2d) 
    	            returns InterferencePolygon2d from Intf;
    ---Purpose: Constructs and computes the auto interference of a Polygon.


    Perform        (me         : in out;
    	    	    Obje1, Obje2 : in Polygon2d);
    ---Purpose: Computes an interference between two Polygons.


    Perform        (me         : in out;
    	    	    Obje       : in Polygon2d);
    ---Purpose: Computes the self interference of a Polygon.


    Pnt2dValue     (me;
    	    	    Index      : in Integer)
		    returns Pnt2d from gp
    	    	    raises OutOfRange from Standard
    	    	    is static;
    ---Purpose: Gives the  geometrical 2d point   of the  intersection
    --          point at address <Index> in the interference.


-- Implementation :

    Interference   (me : in out; Obje1, Obje2 : in Polygon2d)
    	    	    is private;

    Interference   (me : in out; Obje : in Polygon2d)
    	    	    is private;

    Clean          (me   : in out) is private;

    Intersect      (me         : in out;
                    iO, iT     : Integer from Standard;
                    BegO, EndO : in Pnt2d from gp;
                    BegT, EndT : in Pnt2d from gp)
    	    	    is private;
    ---Purpose: Computes the intersection between two segments 
    --          <BegO><EndO> et <BegT><EndT>.

fields

    oClos, tClos         : Boolean from Standard;
    nbso                 : Integer from Standard;

end InterferencePolygon2d;
