-- Created on: 1999-06-10
-- Created by: Vladislav ROMASHKO
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


package TFunction 
    --- Purpose: Function attributes separate data from
    -- algorithms. Each function contains the ID of a function driver.
uses  

    Standard, 
    TCollection,  
    TColStd,
    TDF, 
    TDataStd
 
is 
  
    enumeration ExecutionStatus is
    	ES_WrongDefinition,
	ES_NotExecuted,
	ES_Executing,
	ES_Succeeded,
	ES_Failed;

    deferred class Driver;         

    class DriverTable;   

    class Logbook;

    class DataMapOfGUIDDriver
    instantiates DataMap from TCollection(GUID   from Standard, 
	    	 		       	  Driver from TFunction, 
				          GUID   from Standard);
    class Array1OfDataMapOfGUIDDriver
    instantiates Array1 from TCollection(DataMapOfGUIDDriver from TFunction);
    class HArray1OfDataMapOfGUIDDriver
    instantiates HArray1 from TCollection(DataMapOfGUIDDriver from TFunction,
    	    	    	    	    	  Array1OfDataMapOfGUIDDriver from TFunction);

    class Function; 
    class GraphNode;
    class Scope;

    class IFunction;
    class Iterator;

    class DataMapOfLabelListOfLabel
    instantiates DataMap from TCollection(Label          from TDF, 
	    	 		       	  LabelList      from TDF, 
				          LabelMapHasher from TDF);     
    class DoubleMapOfIntegerLabel
    instantiates DoubleMap from TCollection(Integer from Standard,
    	    	    	    	    	    Label from TDF,
					    MapIntegerHasher from TColStd,
					    LabelMapHasher from TDF);

end TFunction;    
