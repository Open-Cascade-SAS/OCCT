-- Created on: 2000-04-09
-- Created by: Sergey MOZOKHIN
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



package STEPCAFControl

    ---Purpose : This package provides external access and control for STEP,
    --           on the level of CAF (shapes with attributes, external 
    --           references etc.)

uses 
    Dico,
    TCollection,
    TColStd,
    TopTools,
    TopoDS,
    IFSelect,
    Transfer,
    XSControl,
    STEPControl,
    STEPConstruct,
    StepShape,
    StepRepr,
    StepBasic,
    ShapeBuild,
    TDF,
    TDocStd,
    XCAFDoc,
    MoniTool

is

    class Reader;
    	---Purpose: Reader for DECAF documents
    
    class Writer;
    	---Purpose: Writer for DECAF documents

    class ExternFile;
        ---Purpose: Auxiliary class to store results of translation of external file

    class ActorWrite;
    class Controller;
    	---Purpose: Extensions of standard STEP tools for DECAF specifics
    
    class DictionaryOfExternFile instantiates 
    	  Dictionary from Dico (ExternFile from STEPCAFControl);

    class DataMapOfShapeSDR instantiates 
    	  DataMap from TCollection (Shape from TopoDS,
	    	    	    	    ShapeDefinitionRepresentation from StepShape,
				    ShapeMapHasher from TopTools);

    --- skl
    class DataMapOfShapePD instantiates 
    	  DataMap from TCollection (Shape from TopoDS,
	    	    	    	    ProductDefinition from StepBasic,
				    ShapeMapHasher from TopTools);

    class DataMapOfSDRExternFile instantiates 
    	  DataMap from TCollection (ShapeDefinitionRepresentation from StepShape,
				    ExternFile from STEPCAFControl,
				    MapTransientHasher from TColStd);

    --- skl
    class DataMapOfPDExternFile instantiates 
    	  DataMap from TCollection (ProductDefinition from StepBasic,
				    ExternFile from STEPCAFControl,
				    MapTransientHasher from TColStd);

    class DataMapOfLabelShape instantiates
    	  DataMap from TCollection (Label from TDF,
				    Shape from TopoDS,
	    	    	    	    LabelMapHasher from TDF);

    class DataMapOfLabelExternFile instantiates
    	  DataMap from TCollection (Label from TDF,
				    ExternFile from STEPCAFControl,
	    	    	    	    LabelMapHasher from TDF);

end STEPCAFControl;
