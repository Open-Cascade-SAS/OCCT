-- Created on: 1994-04-05
-- Created by: Didier PIFFAULT
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ComparatorOfIndexedVertexOfDelaun from BRepMesh

  ---Purpose: Sort two point in a given direction.


  uses  Boolean from Standard,
        XY from gp,
        DataStructureOfDelaun from BRepMesh

  is      Create (theDir : XY from gp; 
                  TheTol : Real from Standard;
                  HDS    : DataStructureOfDelaun from BRepMesh) 
           returns ComparatorOfIndexedVertexOfDelaun;


         IsLower (me; Left, Right: Integer)
           ---Purpose: returns True if <Left> is lower than <Right>
           returns Boolean from Standard;

         IsGreater (me; Left, Right: Integer)
           ---Purpose: returns True if <Left> is greater than <Right>
           returns Boolean from Standard;

         IsEqual(me; Left, Right: Integer)
           ---Purpose: returns True when <Right> and <Left> are equal.
           returns Boolean from Standard;


         fields  IndexedStructure : DataStructureOfDelaun from BRepMesh;
                 DirectionOfSort  : XY from gp;
                 Tolerance        : Real from Standard;

end ComparatorOfIndexedVertexOfDelaun;
