-- File:	IntImp_COnSCurveTool.cdl
-- Created:	Mon Feb 14 12:19:01 1994
-- Author:	Jacques GOUSSARD
--		<jag@topsn2>
---Copyright:	 Matra Datavision 1994


deferred generic class COnSCurveTool from IntImp (Curve as any)

	---Purpose: Template class for the methods on a curve on surface.
	--          It is possible to implement this class with
	--          an instantiation of the Curve2dTool from Adaptor3d.

uses Pnt2d from gp,
     Vec2d from gp


is

    FirstParameter(myclass;C : Curve ) returns Real;
    
    LastParameter(myclass;C : Curve ) returns Real;

    Value (myclass; C : Curve; U : Real) returns Pnt2d from gp;
    
    D1(myclass; C : Curve ; U : Real; 
    	    	P : out Pnt2d from gp; V : out Vec2d from gp);
		
    Resolution(myclass; C : Curve; Tol3d: Real from Standard)
    
        ---Purpose :  Returns the parametric  resolution corresponding
        --         to the space resolution Tol3d.

    	returns Real from Standard;

end COnSCurveTool;
