-- Created on: 1994-11-17
-- Created by: Marie Jose MARTZ
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class GeomCurve from GeomToIGES inherits GeomEntity from GeomToIGES

    ---Purpose: This class implements the transfer of the Curve Entity from Geom
    --          To IGES. These can be :
    --          Curve
    --            . BoundedCurve
    --               * BSplineCurve
    --               * BezierCurve
    --               * TrimmedCurve
    --            . Conic     
    --               * Circle
    --               * Ellipse
    --               * Hyperbloa
    --               * Line
    --               * Parabola
    --            . OffsetCurve     
  

uses

    Curve                from Geom,
    BoundedCurve         from Geom,
    BSplineCurve         from Geom,
    BezierCurve          from Geom,
    TrimmedCurve         from Geom,
    Conic                from Geom,
    Circle               from Geom,
    Ellipse              from Geom,
    Hyperbola            from Geom,
    Line                 from Geom,
    Parabola             from Geom,
    OffsetCurve          from Geom,
    IGESEntity           from IGESData,
    GeomEntity           from GeomToIGES
    
    
is 
    
    Create returns GeomCurve from GeomToIGES;


    Create(GE : GeomEntity from GeomToIGES)  
    	 returns GeomCurve from GeomToIGES;
    ---Purpose : Creates a tool GeomCurve ready to run and sets its
    --         fields as GE's.

    TransferCurve (me    : in out;
                   start : Curve from Geom;
		   Udeb  : Real  from Standard;
		   Ufin  : Real  from Standard)
    	 returns mutable IGESEntity from IGESData;
    ---Purpose :  Transfert  a  GeometryEntity which  answer True  to  the
    --            member : BRepToIGES::IsGeomCurve(Geometry).  If this
    --            Entity could not be converted, this member returns a NullEntity.


    TransferCurve (me    : in out;
                   start : BoundedCurve from Geom;
		   Udeb  : Real         from Standard;
		   Ufin  : Real         from Standard)
    	 returns mutable IGESEntity from IGESData;


    TransferCurve (me    : in out;
                   start : BSplineCurve from Geom;
		   Udeb  : Real         from Standard;
		   Ufin  : Real         from Standard)
    	 returns mutable IGESEntity from IGESData;


    TransferCurve (me    : in out;
                   start : BezierCurve from Geom;
          	   Udeb  : Real        from Standard;
		   Ufin  : Real        from Standard)
    	 returns mutable IGESEntity from IGESData;

	 
    TransferCurve (me    : in out;
                   start : TrimmedCurve from Geom;
          	   Udeb  : Real        from Standard;
		   Ufin  : Real        from Standard)
    	 returns mutable IGESEntity from IGESData;


    TransferCurve (me    : in out;
                   start : Conic from Geom;
		   Udeb  : Real  from Standard;
		   Ufin  : Real  from Standard)
    	 returns mutable IGESEntity from IGESData;


    TransferCurve (me    : in out;
                    start : Circle from Geom;
 		    Udeb  : Real   from Standard;
		    Ufin  : Real   from Standard)
    	 returns mutable IGESEntity from IGESData;


    TransferCurve (me    : in out;
                   start : Ellipse from Geom;
		   Udeb  : Real    from Standard;
		   Ufin  : Real    from Standard)
    	 returns mutable IGESEntity from IGESData;


    TransferCurve (me    : in out;
                   start : Hyperbola from Geom;
		   Udeb  : Real      from Standard;
		   Ufin  : Real      from Standard)
    	 returns mutable IGESEntity from IGESData;


    TransferCurve (me    : in out;
                   start : Line from Geom;
		   Udeb  : Real from Standard;
		   Ufin  : Real from Standard)
    	 returns mutable IGESEntity from IGESData;


    TransferCurve (me    : in out;
                   start : Parabola from Geom;
	           Udeb  : Real     from Standard;
		   Ufin  : Real     from Standard)
    	 returns mutable IGESEntity from IGESData;


    TransferCurve (me    : in out;
                   start : OffsetCurve from Geom;
 		   Udeb  : Real        from Standard;
		   Ufin  : Real        from Standard)
    	 returns mutable IGESEntity from IGESData;


end GeomCurve;


