-- Created on: 2008-12-10
-- Created by: Pavel TELKOV
-- Copyright (c) 2008-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class MaterialToolDriver from BinMXCAFDoc inherits ADriver from BinMDF

uses
    MessageDriver    from CDM,
    SRelocationTable from BinObjMgt,
    RRelocationTable from BinObjMgt,
    Persistent       from BinObjMgt,
    Attribute        from TDF

is
    Create (theMsgDriver:MessageDriver from CDM)
    returns mutable MaterialToolDriver from BinMXCAFDoc;

    NewEmpty (me)  returns mutable Attribute from TDF
    is redefined;

    Paste(me; theSource     : Persistent from BinObjMgt;
              theTarget     : mutable Attribute from TDF;
              theRelocTable : out RRelocationTable from BinObjMgt)
    returns Boolean from Standard is redefined;

    Paste(me; theSource     : Attribute from TDF;
              theTarget     : in out Persistent from BinObjMgt;
              theRelocTable : out SRelocationTable from BinObjMgt)
    is redefined;

end;
