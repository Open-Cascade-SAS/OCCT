-- Created on: 2000-08-21
-- Created by: Andrey BETENEV
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package ShapeProcess 

    	---Purpose: Shape Processing module
	-- allows to define and apply general Shape Processing as a
	-- customizable sequence of Shape Healing operators. The
	-- customization is implemented via user-editable resource
	-- file which defines sequence of operators to be executed
	-- and their parameters.

uses

    Dico,
    Resource,
    TCollection,
    TColStd,
    GeomAbs,
    TopAbs,
    TopoDS,
    TopTools,
    BRepTools,
    Message,
    ShapeExtend,
    ShapeBuild

is

    class Context; 

    	class ShapeContext;

    deferred class Operator;

	primitive OperFunc;
	class UOperator;

    class OperLibrary;

    class DictionaryOfOperator instantiates 
    	  Dictionary from Dico (Operator from ShapeProcess);

    RegisterOperator (name: CString; op: Operator from ShapeProcess)
    returns Boolean;
    	---Purpose: Registers operator to make it visible for Performer

    FindOperator (name: CString; op: out Operator from ShapeProcess)
    returns Boolean;
    	---Purpose: Finds operator by its name

    Perform (context: Context from ShapeProcess; seq: CString) 
    returns Boolean;
    	---Purpose: Performs a specified sequence of operators on Context
	--          Resource file and other data should be already loaded
	--          to Context (including description of sequence seq)

end ShapeProcess;
