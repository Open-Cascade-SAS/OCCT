-- Created on: 1993-03-10
-- Created by: JCV
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class ConicalSurface from Geom inherits ElementarySurface from Geom

        ---Purpose :  Describes a cone.
    	--    A cone is defined by the half-angle at its apex, and
    	--    is positioned in space by a coordinate system (a
    	--    gp_Ax3 object) and a reference radius as follows:
    	-- - The "main Axis" of the coordinate system is the
    	--   axis of revolution of the cone.
    	-- - The plane defined by the origin, the "X Direction"
    	--   and the "Y Direction" of the coordinate system is
    	--   the reference plane of the cone. The intersection
    	--   of the cone with this reference plane is a circle of
    	--   radius equal to the reference radius.
    	-- - The apex of the cone is on the negative side of
    	--   the "main Axis" of the coordinate system if the
    	--   half-angle is positive, and on the positive side if
    	--   the half-angle is negative.
    	--   This coordinate system is the "local coordinate
    	--   system" of the cone. The following apply:
    	-- - Rotation around its "main Axis", in the
    	--   trigonometric sense given by the "X Direction"
    	--   and the "Y Direction", defines the u parametric direction.
    	-- - Its "X Axis" gives the origin for the u parameter.
    	-- - Its "main Direction" is the v parametric direction of the cone.
    	-- - Its origin is the origin of the v parameter.
    	--   The parametric range of the two parameters is:
    	-- - [ 0, 2.*Pi ] for u, and - ] -infinity, +infinity [ for v
    	--   The parametric equation of the cone is:  P(u, v) =
    	--   O + (R + v*sin(Ang)) * (cos(u)*XDir + sin(u)*YDir) + v*cos(Ang)*ZDir where:
    	-- - O, XDir, YDir and ZDir are respectively
    	--   the origin, the "X Direction", the "Y Direction" and
    	--   the "Z Direction" of the cone's local coordinate system,
    	-- - Ang is the half-angle at the apex of the cone,   and
    	-- - R is the reference radius.
        

uses Ax3      from gp,
     Cone     from gp,
     Pnt      from gp,
     Trsf     from gp,
     GTrsf2d  from gp,
     Vec      from gp,
     Curve    from Geom, 
     Geometry from Geom

raises ConstructionError from Standard,
       RangeError        from Standard

is

  Create (A3 : Ax3; Ang : Real; Radius : Real) 
     returns mutable ConicalSurface
        ---Purpose :
        --  A3 defines the local coordinate system of the conical surface.
        --  Ang is the conical surface semi-angle ]0, PI/2[.
        --  Radius is the radius of the circle Viso in the placement plane 
        --  of the conical surface defined with "XAxis" and "YAxis".
        --  The "ZDirection" of A3 defines the direction of the surface's
        --  axis of symmetry.
        --  If the location point of A3 is the apex of the surface 
        --  Radius = 0 .
        --  At the creation the parametrization of the surface is defined
        --  such that the normal Vector (N = D1U ^ D1V) is oriented towards
        --  the "outside region" of the surface. 
     raises ConstructionError;
        ---Purpose :
        --  Raised if Radius < 0.0 or Ang < Resolution from gp or 
        --  Ang >= PI/2 - Resolution


  Create (C : Cone)   returns mutable ConicalSurface;
        ---Purpose :
        --  Creates a ConicalSurface from a non transient Cone from 
        --  package gp.


  SetCone (me : mutable; C : Cone);
        ---Purpose :
        --  Set <me> so that <me> has the same geometric properties as C.


  SetRadius (me : mutable; R : Real)
        ---Purpose :
        --  Changes the radius of the conical surface in the placement
        --  plane (Z = 0, V = 0).  The local coordinate system is not
        --  modified.
     raises ConstructionError;
        ---Purpose : Raised if R < 0.0


  SetSemiAngle (me : mutable; Ang : Real)
        ---Purpose :
        --  Changes the semi angle of the conical surface.
     raises ConstructionError;
        ---Purpose :
        --  Raised if Ang < Resolution or Ang >= PI/2 - Resolution 


  Cone (me) returns Cone;
        ---Purpose :
        --  returns a non transient cone with the same geometric properties
        --  as <me>.


  UReversedParameter (me; U : Real ) returns Real;
	---Purpose: return 2.PI - U.


  VReversedParameter (me; V : Real ) returns Real;
	---Purpose: Computes the u (or v) parameter on the modified
    	-- surface, when reversing its u (or v) parametric
    	-- direction, for any point of u parameter U (or of v
    	-- parameter V) on this cone.
    	-- In the case of a cone, these functions return respectively:
    	-- - 2.*Pi - U, -V.
  
  
  VReverse (me : mutable)
    	---Purpose : Changes the orientation of this cone in the v
    	-- parametric direction. The bounds of the surface are
    	-- not changed but the v parametric direction is reversed.
    	-- As a consequence, for a cone:
    	-- - the "main Direction" of the local coordinate system
    	--   is reversed, and
    	-- - the half-angle at the apex is inverted.
  is redefined;

  TransformParameters(me; U,V : in out Real; T : Trsf from gp)
	---Purpose: Computes the  parameters on the  transformed  surface for
	--          the transform of the point of parameters U,V on <me>.
	--          
	--          me->Transformed(T)->Value(U',V')
	--          
	--          is the same point as
	--          
	--          me->Value(U,V).Transformed(T)
	--          
	--          Where U',V' are the new values of U,V after calling
	--          
	--          me->TranformParameters(U,V,T)
	--          
	--          This methods multiplies V by T.ScaleFactor()
     is redefined;  

  ParametricTransformation(me; T : Trsf from gp) returns GTrsf2d from gp
	---Purpose: Returns a 2d transformation  used to find the  new
	--          parameters of a point on the transformed surface.
	--          
	--          me->Transformed(T)->Value(U',V')
	--          
	--          is the same point as
	--          
	--          me->Value(U,V).Transformed(T)
	--          
	--          Where U',V' are  obtained by transforming U,V with
	--          th 2d transformation returned by
	--          
	--          me->ParametricTransformation(T)
	--          
	--          This  methods  returns  a scale  centered  on  the
	--          U axis with T.ScaleFactor
     is redefined;  

  Apex (me)  returns Pnt;
    	---Purpose : Computes the apex of this cone. It is on the negative
    	-- side of the axis of revolution of this cone if the
    	-- half-angle at the apex is positive, and on the positive
    	-- side of the "main Axis" if the half-angle is negative.
     


  Bounds (me; U1, U2, V1, V2 : out Real);
        ---Purpose :
        --  The conical surface is infinite in the V direction so 
        --  V1 = Realfirst from Standard and V2 = RealLast.  
        --  U1 = 0 and U2 = 2*PI.


  Coefficients (me; A1, A2, A3, B1, B2, B3, C1, C2, C3, D : out Real);
        ---Purpose :
        --  Returns the coefficients of the implicit equation of the
        --  quadric in the absolute cartesian coordinate system :
        --  These coefficients are normalized.
        --  A1.X**2 + A2.Y**2 + A3.Z**2 + 2.(B1.X.Y + B2.X.Z + B3.Y.Z) +
        --  2.(C1.X + C2.Y + C3.Z) + D = 0.0


  RefRadius (me)   returns Real;
        ---Purpose : Returns the reference radius of this cone.
        -- The reference radius is the radius of the circle formed
        -- by the intersection of this cone and its reference
        -- plane (i.e. the plane defined by the origin, "X
        -- Direction" and "Y Direction" of the local coordinate
        -- system of this cone).
        -- If the apex of this cone is on the origin of the local
        -- coordinate system of this cone, the returned value is 0.
       
     
  SemiAngle (me)  returns Real;
        ---Purpose :
        --  returns the semi-angle of the conical surface ]0.0, PI/2[.


  IsUClosed (me)  returns Boolean;
        ---Purpose : returns True.


  IsVClosed (me)  returns Boolean;
        ---Purpose : returns False.


  IsUPeriodic (me)  returns Boolean;
        ---Purpose : Returns True.


  IsVPeriodic (me)  returns Boolean;
        ---Purpose : Returns False.


  UIso (me; U : Real)  returns mutable Curve;
        ---Purpose : Builds the U isoparametric line of this cone. The
    	--  origin of this line is on the reference plane of this
    	--  cone (i.e. the plane defined by the origin, "X Direction"
    	--  and "Y Direction" of the local coordinate system of this cone).
        

  VIso (me; V : Real)   returns mutable Curve;
        ---Purpose : Builds the V isoparametric circle of this cone. It is the
    	-- circle on this cone, located in the plane of Z
    	-- coordinate V*cos(Semi-Angle) in the local coordinate system of this
    	-- cone. The "Axis" of this circle is the axis of revolution
    	-- of this cone. Its starting point is defined by the "X
    	-- Direction" of this cone.
    	-- Warning
    	-- If the V isoparametric circle is close to the apex of
    	-- this cone, the radius of the circle becomes very small.
    	-- It is possible to have a circle with radius equal to 0.0.
       


  D0 (me; U, V : Real; P : out Pnt);
        ---Purpose :
        --  Computes the  point P (U, V) on the surface.
        --  P (U, V) = Loc +
        --  (RefRadius + V * sin (Semi-Angle)) * (cos (U) * XDir + sin (U) * YDir) +
        --  V * cos (Semi-Angle) * ZDir
        --  where Loc is the origin of the placement plane (XAxis, YAxis)
        --  XDir is the direction of the XAxis and YDir the direction of
        --  the YAxis.


  D1 (me; U, V : Real; P : out Pnt; D1U, D1V : out Vec);
        ---Purpose :
        --  Computes the current point and the first derivatives in the
        --  directions U and V.


  D2 (me; U, V : Real; P : out Pnt; D1U, D1V, D2U, D2V, D2UV : out Vec);
        ---Purpose :
        --  Computes the current point, the first and the second derivatives
        --  in the directions U and V.


  D3 (me; U, V : Real; P : out Pnt;
      D1U, D1V, D2U, D2V, D2UV, D3U, D3V, D3UUV, D3UVV :out Vec);
        ---Purpose :
        --  Computes the current point, the first,the second and the third 
        --  derivatives in the directions U and V.


  DN (me; U, V : Real; Nu, Nv : Integer)   returns Vec
        ---Purpose: Computes the derivative of order Nu in the u
    	-- parametric direction, and Nv in the v parametric
    	-- direction at the point of parameters (U, V) of this cone. 
    	-- Exceptions
    	-- Standard_RangeError if:
    	-- - Nu + Nv is less than 1,
    	-- - Nu or Nv is negative.
    raises RangeError;


  Transform (me : mutable; T : Trsf);
    	---Purpose: Applies the transformation T to this cone.
  Copy (me)  returns mutable like me;

    	---Purpose: Creates a new object which is a copy of this cone.
fields

  radius    : Real;
  semiAngle : Real;

end;
