-- Created on: 1991-09-18
-- Created by: Arnaud BOUZY
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class UnknownIterator from Expr 

	---Purpose: Describes an iterator on NamedUnknowns contained 
	--          in any GeneralExpression.
        ---Level : Internal

uses GeneralExpression from Expr,
    NamedUnknown from Expr,
    MapOfNamedUnknown from Expr

raises NoMoreObject from Standard,
    NoSuchObject from Standard

is

    Create(exp : GeneralExpression)
    returns UnknownIterator;
    
    Perform(me: in out; exp : GeneralExpression)
    is static private;
    
    More(me)
    returns Boolean
    is static;
    
    Next(me : in out)
    raises NoMoreObject
    is static;
    
    Value(me)
    returns NamedUnknown
    raises NoSuchObject
    is static;

fields

    myMap : MapOfNamedUnknown;
    myCurrent : Integer;

end UnknownIterator;
