-- File:	IntTools_FClass2d.cdl
-- Created:	Wed Mar 22 09:29:42 1995
-- Author:	Laurent BUCHARD
--		<lbr@mastox>
---Copyright:	 Matra Datavision 1995


class FClass2d from IntTools

    	---Purpose: Class provides an algorithm to classify a 2d Point
    	---         in 2d space of face using boundaries of the face.

uses  
    Pnt2d             from gp, 
    Face              from TopoDS,
    State             from TopAbs,
    SequenceOfInteger from TColStd,
    SeqOfPtr          from BRepTopAdaptor    

is 
    Create   
    	returns FClass2d from IntTools; 
	---Purpose:
	--- Empty constructor
	---
	    	
    Create( F: Face from TopoDS;  
    	    Tol: Real from Standard)
    	returns FClass2d from IntTools;
	---Purpose:
	--- Initializes algorithm by the face F
	--- and tolerance Tol
	---

    Init  (me:out; 
    	   F: Face from TopoDS;  
    	   Tol: Real from Standard);
    	---Purpose:
	--- Initializes algorithm by the face F
	--- and tolerance Tol
	---
    
    PerformInfinitePoint(me) 
    	returns State from TopAbs;
	---Purpose:
	--- Returns state of infinite 2d point relatively to (0, 0)
	---
    
    Perform(me;  
    	    Puv: Pnt2d from gp;  
    	    RecadreOnPeriodic: Boolean from Standard=Standard_True) 
    	returns State from TopAbs;
	---Purpose:
	--- Returns state of the 2d point Puv.
	--- If RecadreOnPeriodic is true (defalut value),
	--- for the periodic surface 2d point, adjusted to period, is
	--- classified.
	---
    
    Destroy(me: in out);
    	---C++: alias ~
    	---Purpose:
	--- Destructor
	---


    TestOnRestriction(me;  
    	    	    	Puv: Pnt2d from gp; 
                        Tol: Real from Standard;
                        RecadreOnPeriodic: Boolean from Standard  =  Standard_True) 
    	returns State from TopAbs;
    	---Purpose: 
    	--- Test a point with +- an offset (Tol) and returns
    	--- On if some points are OUT an some are IN
    	--  (Caution: Internal use . see the code for more details)
	---

--modified by NIZNHY-PKV Mon May 29 10:47:52 2006f 
    IsHole(me) 
	returns Boolean from Standard; 
--modified by NIZNHY-PKV Mon May 29 10:47:54 2006t

fields 

    TabClass    : SeqOfPtr          from BRepTopAdaptor;
    TabOrien    : SequenceOfInteger from TColStd;
    Toluv       : Real              from Standard;
    Face        : Face              from TopoDS;
    U1          : Real              from Standard;
    V1          : Real              from Standard;    
    U2          : Real              from Standard;
    V2          : Real              from Standard;
    
    Umin        : Real              from Standard;  
    Umax        : Real              from Standard;
    Vmin        : Real              from Standard;  
    Vmax        : Real              from Standard; 
    --modified by NIZNHY-PKV Mon May 29 10:44:12 2006f 
    myIsHole    : Boolean           from Standard; 
    --modified by NIZNHY-PKV Mon May 29 10:44:14 2006t


end FClass2d ;
