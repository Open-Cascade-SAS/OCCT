-- Created on: 1995-01-27
-- Created by: Marie Jose MARTZ
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class BRShell from BRepToIGES inherits BREntity from BRepToIGES

    ---Purpose: This class implements the transfer of Shape Entities from Geom
    --          To IGES. These can be :
    --            . Vertex
    --            . Edge
    --            . Wire
  

uses

    Shape                from TopoDS,
    Face                 from TopoDS,
    Shell                from TopoDS,
    IGESEntity           from IGESData,
    BREntity             from BRepToIGES    
    
is 
    
    Create 
    	returns BRShell from BRepToIGES;
    
    Create (BR : BREntity from BRepToIGES)
    	returns BRShell from BRepToIGES;    


    TransferShell (me    : in out;
                   start : Shape from TopoDS)
    	returns mutable IGESEntity from IGESData;
    ---Purpose :  Transfert an Shape entity from TopoDS to IGES
    --            This entity must be a Face or a Shell.
    --            If this Entity could not be converted, this member returns a NullEntity.


    TransferShell (me    : in out;
                   start : Shell from TopoDS)
    	returns mutable IGESEntity from IGESData;
    ---Purpose :  Transfert an Shell entity from TopoDS to IGES
    --            If this Entity could not be converted, this member returns a NullEntity.


    TransferFace (me    : in out;
                  start : Face from TopoDS)
    	returns mutable IGESEntity from IGESData;
    ---Purpose :  Transfert a Face entity from TopoDS to IGES
    --            If this Entity could not be converted, this member returns a NullEntity.


end BRShell;
