-- File:	RWStepShape_RWSubedge.cdl
-- Created:	Fri Jan  4 17:42:45 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class RWSubedge from RWStepShape

    ---Purpose: Read & Write tool for Subedge

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    Subedge from StepShape

is
    Create returns RWSubedge from RWStepShape;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : Subedge from StepShape);
	---Purpose: Reads Subedge

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: Subedge from StepShape);
	---Purpose: Writes Subedge

    Share (me; ent : Subedge from StepShape;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWSubedge;
