-- Created on: 1996-01-12
-- Created by: Denis PASCAL
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PlanarRadius from DrawDim inherits PlanarDimension from DrawDim

	---Purpose: 

uses Shape   from TopoDS,
     Face    from TopoDS,
     Color   from Draw,
     Display from Draw

is

    Create (plane  : Face  from TopoDS;
            circle : Shape from TopoDS)
    returns mutable PlanarRadius from DrawDim;    

    Create (circle : Shape from TopoDS)
    returns mutable PlanarRadius from DrawDim;
    
    DrawOn(me; dis : in out Display);
    

fields

    myCircle : Shape from TopoDS;

end PlanarRadius;
