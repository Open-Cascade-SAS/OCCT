-- Created on: 1999-03-10
-- Created by: data exchange team
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class AppliedOrganizationAssignment from StepAP214 
inherits OrganizationAssignment from StepBasic
       
uses
    	HArray1OfOrganizationItem from StepAP214, 
	OrganizationItem from StepAP214, 
	Organization from StepBasic,
	OrganizationRole from StepBasic


is
    
    Create returns mutable AppliedOrganizationAssignment;
	---Purpose: Returns a AppliedOrganizationAssignment


	Init (me : mutable;
	      aAssignedOrganization : mutable Organization from StepBasic;
	      aRole : mutable OrganizationRole from StepBasic) is redefined;

	Init (me : mutable;
	      aAssignedOrganization : mutable Organization from StepBasic;
	      aRole : mutable OrganizationRole from StepBasic;
	      aItems : mutable HArray1OfOrganizationItem from StepAP214) is virtual;

	-- Specific Methods for Field Data Access --

	SetItems(me : mutable; aItems : mutable HArray1OfOrganizationItem);
	Items (me) returns mutable HArray1OfOrganizationItem;
	ItemsValue (me; num : Integer) returns OrganizationItem;
	NbItems (me) returns Integer;
    
fields

    	items : HArray1OfOrganizationItem from StepAP214; -- a SelectType

end AppliedOrganizationAssignment;
