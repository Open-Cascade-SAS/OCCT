-- Created on: 1997-01-22
-- Created by: Mister rmi
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class FWOSDriver from CDF  inherits MetaDataDriver from CDF
uses
    MetaData from CDM,
    Document from CDM,
    ExtendedString from TCollection
is
    Create
    returns FWOSDriver from CDF;
    ---Purpose: initializes the MetaDatadriver with its specific name.


    	
    Find(me: mutable; aFolder, aName, aVersion: ExtendedString from TCollection)
    returns Boolean from Standard;
    ---Purpose: indicate whether a file exists corresponding to the folder and the name
    
    HasReadPermission(me: mutable; aFolder, aName, aVersion: ExtendedString from TCollection)
    returns Boolean from Standard;

    
    MetaData(me: mutable; aFolder, aName, aVersion: ExtendedString from TCollection)
    returns MetaData from CDM
    is  private;
    
    CreateMetaData(me: mutable; aDocument: Document from CDM;
    	         aFileName: ExtendedString from TCollection)
    returns  MetaData from CDM
    is  private;
    
    FindFolder(me: mutable; aFolder: ExtendedString from TCollection)
    returns Boolean from Standard;


   DefaultFolder(me: mutable) returns ExtendedString from TCollection;
   
   BuildFileName(me: mutable; aDocument: Document from CDM)
   returns ExtendedString from TCollection;
    
   Concatenate(myclass; aFolder,aName:  ExtendedString from TCollection)
   returns ExtendedString from TCollection
   is private;


   BuildMetaData(me: mutable; aFileName: ExtendedString from TCollection)
   returns MetaData from CDM
   is  private;

   SetName(me: mutable; aDocument: Document from CDM; aName: ExtendedString from TCollection)
   returns ExtendedString from TCollection
   is redefined;
   
end FWOSDriver from CDF;
