-- Created on: 2001-12-28
-- Created by: Andrey BETENEV
-- Copyright (c) 2001-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1

class ConnectedEdgeSet from StepShape
inherits TopologicalRepresentationItem from StepShape

    ---Purpose: Representation of STEP entity ConnectedEdgeSet

uses
    HAsciiString from TCollection,
    HArray1OfEdge from StepShape

is
    Create returns ConnectedEdgeSet from StepShape;
	---Purpose: Empty constructor

    Init (me: mutable; aRepresentationItem_Name: HAsciiString from TCollection;
                       aCesEdges: HArray1OfEdge from StepShape);
	---Purpose: Initialize all fields (own and inherited)

    CesEdges (me) returns HArray1OfEdge from StepShape;
	---Purpose: Returns field CesEdges
    SetCesEdges (me: mutable; CesEdges: HArray1OfEdge from StepShape);
	---Purpose: Set field CesEdges

fields
    theCesEdges: HArray1OfEdge from StepShape;

end ConnectedEdgeSet;
