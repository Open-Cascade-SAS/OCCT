-- Created on: 1998-02-04
-- Created by: Christian CAILLET
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



deferred class SignType  from Interface    inherits SignText from MoniTool

    	---Purpose : Provides the basic service to get a type name, according
    	--           to a norm
    	--           It can be used for other classes (general signatures ...)

uses CString, Transient, AsciiString, InterfaceModel

is

--    Name (me) returns CString  is deferred;  already in SignText
    ---Purpose : Returns an identification of the Signature (a word), given at
    --           initialization time

    Text  (me; ent : any Transient; context : any Transient)
    	returns AsciiString from TCollection;
    ---Purpose : Specialised to consider context as an InterfaceModel


    Value (me; ent : any Transient; model : InterfaceModel)
    	returns CString  is deferred;
    ---Purpose : Returns the Signature for a Transient object. It is specific
    --           of each sub-class of Signature. For a Null Handle, it should
    --           provide ""
    --           It can work with the model which contains the entity

    ClassName (myclass; typnam : CString) returns CString;
    ---Purpose : From a CDL Type Name, returns the Class part (package dropped)
    --           WARNING : buffered, to be immediately copied or printed

end SignType;
