-- Created on: 1993-05-07
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class VPointInterIterator from TopOpeBRep

    -- ==========================
    -- Restriction Point iterator
    -- ==========================

uses

    LineInter from TopOpeBRep,
    PLineInter from TopOpeBRep,
    VPointInter from TopOpeBRep

is

    Create returns VPointInterIterator from TopOpeBRep;
    Create(LI : LineInter from TopOpeBRep)  
    returns VPointInterIterator from TopOpeBRep;

    Init(me:in out; LI : LineInter from TopOpeBRep;
    	    	    checkkeep : Boolean from Standard = Standard_False) is static;
    Init(me:in out) is static;
    More(me) returns Boolean is static;
    Next(me:in out) is static;
 
    CurrentVP(me:in out) returns VPointInter from TopOpeBRep is static;
    ---C++: return const &

    CurrentVPIndex(me) returns Integer is static;

    ChangeCurrentVP(me:in out) returns VPointInter from TopOpeBRep is static;
    ---C++: return &

    PLineInterDummy(me) returns PLineInter from TopOpeBRep;
    
fields

    myLineInter : PLineInter from TopOpeBRep;
    myVPointIndex : Integer;    
    myVPointNb : Integer;
    mycheckkeep : Boolean from Standard;

end VPointInterIterator from TopOpeBRep;
