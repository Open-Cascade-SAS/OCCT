-- Created on: 1993-01-14
-- Created by: Philippe DAUTRY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Builder from BRepSweep 

	---Purpose: implements the abstract Builder with the BRep Builder

uses
    Builder from BRep,
        
    Shape	from TopoDS,
    Shell	from TopoDS,
    Face	from TopoDS,
    Wire	from TopoDS,
    Edge	from TopoDS,
    Vertex	from TopoDS,
    
    Orientation from TopAbs
    
is

    Create(aBuilder : Builder from BRep) returns Builder from BRepSweep;
	---Purpose: Creates a Builder.
	
    Builder(me) returns Builder from BRep
	---C++: inline
	---C++: return const &
    is static;
	
        -- implements the Builder methods

    MakeCompound (me; aCompound : out Shape from TopoDS)
    	---Purpose: Returns an empty Compound.
    is static;

    MakeCompSolid (me; aCompSolid : out Shape from TopoDS)
    	---Purpose: Returns an empty CompSolid.
    is static;

    MakeSolid (me; aSolid : out Shape from TopoDS)
    	---Purpose: Returns an empty Solid.
    is static;

    MakeShell (me; aShell : out Shape from TopoDS)
    	---Purpose: Returns an empty Shell.
    is static;

    MakeWire (me; aWire : out Shape from TopoDS)
    	---Purpose: Returns an empty Wire.
    is static;

    
    Add(me; aShape1 : in out Shape from TopoDS; 
	    aShape2 : in     Shape from TopoDS;
    	    Orient  : in     Orientation from TopAbs)
    	---Purpose: Adds the Shape 1 in the Shape 2, set to
    	--          <Orient> orientation.
    is static;
    
    Add(me; aShape1 : in out Shape from TopoDS; 
	    aShape2 : in     Shape from TopoDS)
    	---Purpose: Adds the Shape 1 in the Shape 2.
    is static;

fields

    myBuilder : Builder from BRep;

end Builder;

