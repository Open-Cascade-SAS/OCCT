-- Created on: 1999-06-18
-- Created by: Sergei ZERTCHANINOV
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class FaceConnect  from ShapeFix

    ---Purpose : 

uses 
    DataMapOfShapeListOfShape from TopTools,
    Face from TopoDS, Shell from TopoDS

is

    Create returns FaceConnect from ShapeFix;

    Add (me : in out; aFirst : Face from TopoDS; aSecond : Face from TopoDS)
    returns Boolean from Standard;
    ---Purpose : 

    Build (me : in out; shell : Shell from TopoDS;
    	   sewtoler : Real from Standard; fixtoler : Real from Standard)
    returns Shell from TopoDS;
    ---Purpose : 

    Clear (me : in out);
    ---Purpose : Clears internal data structure

fields

    myConnected    : DataMapOfShapeListOfShape from TopTools;
    	-- Map of pairs (face, list of connected faces) - to store connectivity info
    myOriFreeEdges : DataMapOfShapeListOfShape from TopTools;
    	-- Map of pairs (face, list of original free edges)
    myResFreeEdges : DataMapOfShapeListOfShape from TopTools;
    	-- Map of pairs (free edge, list of result free edges)
    myResSharEdges : DataMapOfShapeListOfShape from TopTools;
    	-- Map of pairs (free edge, list of result shared edges)

end FaceConnect;
