-- Created on: 1996-04-01
-- Created by: Philippe MANGIN
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



private class DistributionOfJerk from FairCurve inherits  DistributionOfEnergy  from FairCurve

	---Purpose: Compute the "Jerk" distribution.

uses  Vector        from math, 
      FunctionSet   from math,
      HArray1OfReal  from TColStd,
      HArray1OfPnt2d from TColgp,
      BattenLaw  from FairCurve


is
    Create( BSplOrder :  Integer;
            FlatKnots :  HArray1OfReal;
	    Poles     :  HArray1OfPnt2d;
	    DerivativeOrder : Integer; 
	    Law       :  BattenLaw;
            NbValAux  : Integer = 0) returns DistributionOfJerk;
	    

    Value(me: in out; X: Vector; F: out Vector)
    	---Purpose: computes the values <F> of the functions for the 
    	--          variable <X>.
    	--          returns True if the computation was done successfully, 
    	--          False otherwise.

    returns Boolean is redefined;
    

fields
    MyLaw           : BattenLaw;
end DistributionOfJerk;
