-- Created on: 1992-11-05
-- Created by: Remi LEQUETTE
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class Torus from BRepPrim inherits Revolution from BRepPrim

	---Purpose: Implements the torus primitive

uses
    Face from TopoDS,
    
    Pnt from gp,
    Ax2 from gp    

raises
    DomainError

is
    Create(Position : Ax2 from gp; Major : Real; Minor : Real)
    returns Torus from BRepPrim
	   ---Purpose: the STEP definition
	   --          Position : center and axes
	   --          Major, Minor : Radii
	   --          
	   --          Errors : Major < Resolution
	   --                   Minor < Resolution
    raises DomainError;

    Create(Major,Minor : Real)
    returns Torus from BRepPrim
	---Purpose: Torus centered at origin
    raises DomainError;
    
    Create(Center : Pnt from gp; Major, Minor : Real)
    returns Torus from BRepPrim
	---Purpose: Torus at Center
    raises DomainError;
    
    MakeEmptyLateralFace(me) returns Face from TopoDS
	---Purpose: The surface normal should be directed  towards the
	--          outside.
    is redefined;
    
    SetMeridian(me : in out)
    is static private;
    
fields
    myMajor     : Real;
    myMinor     : Real;

end Torus;
