-- Created on: 2005-04-18
-- Created by: Eugeny NAPALKOV <eugeny.napalkov@opencascade.com>
-- Copyright (c) 2005-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package BinXCAFDrivers

uses
    Standard,
    CDM,
    BinMDF,
    BinDrivers
is
    class DocumentStorageDriver;
    class DocumentRetrievalDriver;

    Factory (theGUID : GUID from Standard) returns Transient from Standard;
    ---C++: return const &

    AttributeDrivers (MsgDrv : MessageDriver from CDM)
    	returns ADriverTable from BinMDF;
    	---Purpose: Creates the table of drivers of types supported
end;    
