-- Created on: 2000-10-31
-- Created by: Vladislav ROMASHKO
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Limitation from QANewBRepNaming inherits BooleanOperationFeat from QANewBRepNaming

uses

    Label from TDF, 
    MakeShape from BRepBuilderAPI,
    Limitation from QANewModTopOpe

is
 
    Create returns Limitation from QANewBRepNaming;

    Create(ResultLabel : Label from TDF) 
    returns Limitation from QANewBRepNaming;

    Load (me; MakeShape : in out Limitation from QANewModTopOpe); 
     
    LoadContent(me; MakeShape : in out Limitation from QANewModTopOpe)
    ---Purpose: Loads the content of the result.
    is protected;

    LoadResult(me; MakeShape : in out Limitation from QANewModTopOpe)
    ---Purpose: Loads the result.
    is protected;

    LoadDegenerated(me; MakeShape : in out Limitation from QANewModTopOpe)
    ---Purpose: Loads the deletion of the degenerated edges.
    is protected;    


    LoadWire(me; MakeShape : in out Limitation from QANewModTopOpe)
    ---Purpose: A default implementation for naming of a wire as an object of
    --          a boolean operation.
    is protected;

    LoadShell(me; MakeShape : in out Limitation from QANewModTopOpe)
    ---Purpose: A default implementation for naming of a shell as an object of
    --          a boolean operation.
    is protected;

end Limitation;
