-- File:        ContextDependentInvisibility.cdl
-- Created:     Mon Dec  4 12:02:24 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWContextDependentInvisibility from RWStepVisual

	---Purpose : Read & Write Module for ContextDependentInvisibility

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     ContextDependentInvisibility from StepVisual,
     EntityIterator from Interface

is

	Create returns RWContextDependentInvisibility;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable ContextDependentInvisibility from StepVisual);

	WriteStep (me; SW : in out StepWriter; ent : ContextDependentInvisibility from StepVisual);

	Share(me; ent : ContextDependentInvisibility from StepVisual; iter : in out EntityIterator);

end RWContextDependentInvisibility;
