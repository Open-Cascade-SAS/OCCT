-- Created on: 2000-07-03
-- Created by: Andrey BETENEV
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1

class ProductDefinitionRelationship from StepBasic
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity ProductDefinitionRelationship

uses
    HAsciiString from TCollection,
    ProductDefinition from StepBasic

is
    Create returns ProductDefinitionRelationship from StepBasic;
	---Purpose: Empty constructor

    Init (me: mutable; aId: HAsciiString from TCollection;
                       aName: HAsciiString from TCollection;
                       hasDescription: Boolean;
                       aDescription: HAsciiString from TCollection;
                       aRelatingProductDefinition: ProductDefinition from StepBasic;
                       aRelatedProductDefinition: ProductDefinition from StepBasic);
	---Purpose: Initialize all fields (own and inherited)

    Id (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Id
    SetId (me: mutable; Id: HAsciiString from TCollection);
	---Purpose: Set field Id

    Name (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Name
    SetName (me: mutable; Name: HAsciiString from TCollection);
	---Purpose: Set field Name

    Description (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Description
    SetDescription (me: mutable; Description: HAsciiString from TCollection);
	---Purpose: Set field Description
    HasDescription (me) returns Boolean;
	---Purpose: Returns True if optional field Description is defined

    RelatingProductDefinition (me) returns ProductDefinition from StepBasic;
	---Purpose: Returns field RelatingProductDefinition
    SetRelatingProductDefinition (me: mutable; RelatingProductDefinition: ProductDefinition from StepBasic);
	---Purpose: Set field RelatingProductDefinition

    RelatedProductDefinition (me) returns ProductDefinition from StepBasic;
	---Purpose: Returns field RelatedProductDefinition
    SetRelatedProductDefinition (me: mutable; RelatedProductDefinition: ProductDefinition from StepBasic);
	---Purpose: Set field RelatedProductDefinition

fields
    theId: HAsciiString from TCollection;
    theName: HAsciiString from TCollection;
    theDescription: HAsciiString from TCollection; -- optional
    theRelatingProductDefinition: ProductDefinition from StepBasic;
    theRelatedProductDefinition: ProductDefinition from StepBasic;
    defDescription: Boolean; -- flag "is Description defined"

end ProductDefinitionRelationship;
