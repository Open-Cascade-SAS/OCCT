-- Created on: 1996-12-05
-- Created by: Flore Lantheaume/Odile Olivier
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ConcentricRelation from AIS inherits Relation from AIS

	---Purpose: A framework to define a constraint by a relation of
    	-- concentricity between two or more interactive datums.
    	-- The display of this constraint is also defined.
    	-- A plane is used to create an axis along which the
    	-- relation of concentricity can be extended.

uses

    PresentationManager3d from PrsMgr,
    Presentation          from Prs3d,
    Selection             from SelectMgr,
    Shape                 from TopoDS,
    Pnt                   from gp,
    Dir                   from gp,
    Projector             from Prs3d,
    Transformation        from Geom,
    Plane                 from Geom
    
is
    Create (aFShape     : Shape          from TopoDS;
    	    aSShape     : Shape          from TopoDS;
	    aPlane      : Plane          from Geom)
	 ---Purpose: Constructs the display object for concentric relations
    	 -- between shapes.
    	 -- This object is defined by the two shapes, aFShape
    	 -- and aSShape and the plane aPlane.
    	 -- aPlane is provided to create an axis along which the
    	 -- relation of concentricity can be extended. 
    returns mutable ConcentricRelation from AIS;

    -- Methods from PresentableObject
    
    Compute(me            : mutable;
  	    aPresentationManager: PresentationManager3d from PrsMgr;
    	    aPresentation : mutable Presentation from Prs3d;
    	    aMode         : Integer from Standard= 0) 
    is redefined static private;
    
    Compute(me:mutable;
    	        aProjector: Projector from Prs3d;
                aPresentation: mutable Presentation from Prs3d)
    is redefined static private;     
    
    Compute(me            : mutable;
    	    aProjector    : Projector from Prs3d;
    	    aTrsf         : Transformation from Geom;
	    aPresentation : mutable Presentation from Prs3d)
    is redefined;
	 ---Purpose: computes the presentation according to a point of view
	 --          given by <aProjector>. 
         --          To be Used when the associated degenerated Presentations 
	 --          have been transformed by <aTrsf> which is not a Pure
	 --          Translation. The HLR Prs can't be deducted automatically
	 --          WARNING :<aTrsf> must be applied
	 --           to the object to display before computation  !!!

    ComputeTwoEdgesConcentric(me:mutable;
    	    	    	      aPresentationManager: Presentation from Prs3d)
    is private;	
			      
    ComputeEdgeVertexConcentric(me:mutable;
    	    	    	        aPresentationManager: Presentation from Prs3d)
    is private;	
    
    ComputeTwoVerticesConcentric(me:mutable;
    	    	    	         aPresentationManager: Presentation from Prs3d)
    is private;	
    
    -- Methods from SelectableObject
   
    ComputeSelection(me         : mutable;
    	    	     aSelection : mutable Selection from SelectMgr;
    	    	     aMode      : Integer from Standard)
    is redefined private;
    
fields
    
    myCenter    : Pnt   from gp;
    myRad       : Real  from Standard;
    myDir       : Dir   from gp;
    myPnt       : Pnt   from gp;

end ConcentricRelation;
