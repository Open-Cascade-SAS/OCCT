-- Created on: 1999-07-22
-- Created by: data exchange team
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ShapeDivideClosed from ShapeUpgrade inherits ShapeDivide from ShapeUpgrade

	---Purpose: Divides all closed faces in the shape. Class 
    	--          ShapeUpgrade_ClosedFaceDivide is used as divide tool.

uses

    Shape from TopoDS

is
    Create (S: Shape from TopoDS) returns ShapeDivideClosed from ShapeUpgrade;
    	---Purpose: Initialises tool with shape and default parameter.
    
    SetNbSplitPoints (me: in out; num: Integer);
    	---Purpose: Sets the number of cuts applied to divide closed faces.
	--          The number of resulting faces will be num+1.
    

end ShapeDivideClosed;
