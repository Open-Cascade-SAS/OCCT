-- Created on: 1993-06-23
-- Created by: Didier PIFFAULT
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Tool from Intf

	---Purpose: Provides services to create box for infinites 
	--          lines in a given contexte. 

uses    Integer from Standard,
    	Real from Standard,
	Box2d from Bnd,
	Lin2d from gp,
	Hypr2d from gp,
	Parab2d from gp,
	Conic from IntAna2d,
	Box from Bnd,
	Lin from gp,
	Hypr from gp,
	Parab from gp


raises  OutOfRange  from Standard


is      Create returns Tool from Intf;

    	Lin2dBox   (me         : in out;
    	    	    theLin2d   : in  Lin2d   from gp;
    	    	    bounding   : in  Box2d   from Bnd;
    	    	    boxLin     : out Box2d   from Bnd)
    	    is static;

    	Hypr2dBox  (me         : in out;
    	    	    theHypr2d  : in  Hypr2d  from gp;
    	    	    bounding   : in  Box2d   from Bnd;
    	    	    boxHypr    : out Box2d   from Bnd)
    	    is static;

    	Inters2d   (me         : in out;
    	    	    theCurve   : in  Hypr2d  from gp;
    	    	    Domain     : in  Box2d   from Bnd)
    	    	returns Integer from Standard is static private;

    	Parab2dBox (me         : in out;
    	    	    theParab2d : in  Parab2d from gp;
    	    	    bounding   : in  Box2d   from Bnd;
    	    	    boxHypr    : out Box2d   from Bnd)
    	    is static;

    	Inters2d   (me         : in out;
    	    	    theCurve   : in  Parab2d from gp;
    	    	    Domain     : in  Box2d   from Bnd)
    	    	returns Integer from Standard is static private;


    	LinBox     (me       : in out;
    	    	    theLin   : in  Lin from gp;
    	    	    bounding : in  Box from Bnd;
    	    	    boxLin   : out Box from Bnd)
    	    is static;

    	HyprBox    (me       : in out;
    	    	    theHypr  : in  Hypr from gp;
    	    	    bounding : in  Box  from Bnd;
    	    	    boxHypr  : out Box  from Bnd)
    	    is static;

    	Inters3d   (me         : in out;
    	    	    theCurve   : in  Hypr  from gp;
    	    	    Domain     : in  Box   from Bnd)
    	    	returns Integer from Standard is static private;

    	ParabBox   (me       : in out;
    	    	    theParab : in  Parab from gp;
    	    	    bounding : in  Box   from Bnd;
    	    	    boxHypr  : out Box   from Bnd)
    	    is static;

    	Inters3d   (me         : in out;
    	    	    theCurve   : in Parab from gp;
    	    	    Domain     : in Box   from Bnd)
    	    	returns Integer from Standard is static private;


    	NbSegments (me)
	    	returns Integer from Standard
    	    is static;

    	BeginParam (me;
	    	    SegmentNum : Integer from Standard)
		returns Real from Standard
    	    	raises OutOfRange  from Standard
    	    is static;

    	EndParam   (me;
	    	    SegmentNum : Integer from Standard)
		returns Real from Standard
    	    	raises OutOfRange  from Standard
    	    is static;


fields  nbSeg         : Integer from Standard;
    	beginOnCurve  : Real    from Standard [6];
    	endOnCurve    : Real    from Standard [6];
      
      -- Code of every side of BndBox. 
        bord          : Integer from Standard [12];
        
        xint          : Real    from Standard [12];
        yint          : Real    from Standard [12];
        zint          : Real    from Standard [12];
        parint        : Real    from Standard [12];

end Tool;
