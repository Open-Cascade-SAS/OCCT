-- Created on: 1991-02-22
-- Created by: Jean Claude Vauthier
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




package GCPnts
        --- Purpose :
        --  This package  contains the geometric  algorithmes  used to
        --  compute characteristic points on parametrized curves.
        --  
        --  They are  high  level  algorithms based  on  the low level
        --  algorithms in CPnts.
    	---Level : Public. 
    	--  All methods of all  classes will be public.

uses Standard, TCollection, CPnts, Adaptor3d, Adaptor2d  , gp, GeomAbs,
     TColgp, StdFail, TColStd

is

   enumeration AbscissaType 
         is LengthParametrized, Parametrized, AbsComposite end;
	 
   enumeration DeflectionType 
         is Linear, Circular, Curved, DefComposite end;

   class AbscissaPoint;
   
   class UniformAbscissa;
   
   class UniformDeflection;

   class QuasiUniformDeflection;

   class QuasiUniformAbscissa;

   class TangentialDeflection;
   
end GCPnts;





