-- Created on: 1997-11-19
-- Created by: Denis PASCAL
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- modified     Sergey Zaritchny



class Geometry from PDataXtd inherits Attribute from PDF

	---Purpose: 

uses Integer          from Standard,
     Real             from PDataStd,
     HAttributeArray1 from PDF
    
is

    Create returns mutable Geometry from  PDataXtd;
    
    Create (Type : Integer from Standard)
    returns mutable Geometry from PDataXtd;
    
    GetType (me) returns Integer from Standard;
    
    SetType (me : mutable; Type : Integer from Standard);
    
fields

    myType : Integer from Standard;

end Geometry;
