-- Created on: 1994-11-04
-- Created by: Christian CAILLET
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

generic class Mapper from Transfer
    (TheKey    as  any;
     TheHasher as  any;
     TheInfo   as  any)
        inherits Finder

    ---Purpose : a Mapper defines a Finder for a specific input class
    --           its definition includes the value of the Key to be mapped,
    --           and the HashCoder associated to the class of the Key
    --           
    --           TheKey defines the class to be keyed
    --           TheHasher is the associated Hasher
    --           TheInfo   is an additionnal class which helps to provide
    --             informations on the value (template : see DataInfo)

uses CString

is

    Create (akey : any TheKey) returns Mapper;
    ---Purpose : Creates a Mapper with a Value. This Value can then not be
    --           changed. It is used by the Hasher to compute the HashCode,
    --           which will then be stored for an immediate reading.

    Value (me) returns any TheKey  is static;
    ---Purpose : Returns the contained value
    ---C++ : return const &

    Equates (me; other : Finder) returns Boolean;
    ---Purpose : Specific testof equallity : defined as False if <other> has
    --           not the same true Type, else contents are compared (by
    --           C++ operator ==)

    ValueType    (me) returns Type  is redefined;
    ---Purpose : Returns the Type of the Value. By default, returns the
    --           DynamicType of <me>, but can be redefined

    ValueTypeName (me) returns CString  is redefined;
    ---Purpose : Returns the name of the Type of the Value. Default is name
    --           of ValueType, unless it is for a non-handled object

fields

    theval  : TheKey;

end Mapper;
