-- File:	RWStepBasic_RWCharacterizedObject.cdl
-- Created:	Thu May 11 16:38:00 2000 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class RWCharacterizedObject from RWStepBasic

    ---Purpose: Read & Write tool for CharacterizedObject

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    CharacterizedObject from StepBasic

is
    Create returns RWCharacterizedObject from RWStepBasic;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : CharacterizedObject from StepBasic);
	---Purpose: Reads CharacterizedObject

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: CharacterizedObject from StepBasic);
	---Purpose: Writes CharacterizedObject

    Share (me; ent : CharacterizedObject from StepBasic;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWCharacterizedObject;
