-- Created on: 1992-10-22
-- Created by: Laurent BUCHARD
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Geom2dCurveTool from Geom2dInt


	---Purpose: This class provides a Geom2dCurveTool as < Geom2dCurveTool from IntCurve >
	--          from a Tool as < Geom2dCurveTool from Adaptor3d > .

uses 

     Pnt2d        from gp,
     Vec2d        from gp,
     Lin2d        from gp,
     Circ2d       from gp,
     Elips2d      from gp,
     Parab2d      from gp,
     Hypr2d       from gp,
     Array1OfReal from TColStd,
     CurveType    from GeomAbs,
     Curve2d      from Adaptor2d


is


    GetType(myclass; C: Curve2d from Adaptor2d)
    	---C++: inline
    	returns CurveType from GeomAbs;

    IsComposite(myclass; C:  Curve2d from Adaptor2d)
        ---C++: inline
    	returns Boolean from Standard;

    Line(myclass; C: Curve2d from Adaptor2d)
    
	---Purpose: Returns the Lin2d from gp corresponding to the curve C.
	--          This method is called only when TheType returns
	--          GeomAbs_Line.
        ---C++: inline
    	returns Lin2d from gp;

 
    Circle(myclass; C: Curve2d from Adaptor2d)
    
	---Purpose: Returns the Circ2d from gp corresponding to the curve C.
	--          This method is called only when TheType returns
	--          GeomAbs_Circle.
        ---C++: inline
    	returns Circ2d from gp;


    Ellipse(myclass; C: Curve2d from Adaptor2d)
    
	---Purpose: Returns the Elips2d from gp corresponding to the curve C.
	--          This method is called only when TheType returns
	--          GeomAbs_Ellipse.
        ---C++: inline
    	returns Elips2d from gp;


    Parabola(myclass; C: Curve2d from Adaptor2d)
    
	---Purpose: Returns the Parab2d from gp corresponding to the curve C.
	--          This method is called only when TheType returns
	--          GeomAbs_Parabola.
        ---C++: inline
    	returns Parab2d from gp;


    Hyperbola(myclass; C: Curve2d from Adaptor2d)
    
	---Purpose: Returns the Hypr2d from gp corresponding to the curve C.
	--          This method is called only when TheType returns
	--          GeomAbs_Hyperbola.
        ---C++: inline
    	returns Hypr2d from gp;


-- The following method are used only when TheType returns  IntCurve_Other.


    EpsX (myclass; C: Curve2d from Adaptor2d)
        ---C++: inline
    	returns Real;

    EpsX (myclass; C: Curve2d from Adaptor2d;
                   Eps_XYZ : Real from Standard)
        ---C++: inline
    	returns Real;


    NbSamples(myclass; C: Curve2d from Adaptor2d)

    	returns Integer;

    NbSamples(myclass; C: Curve2d from Adaptor2d; U0,U1: Real from Standard)

    	returns Integer;


    FirstParameter(myclass; C:Curve2d from Adaptor2d)
        ---C++: inline
    	returns Real;


    LastParameter(myclass; C:Curve2d from Adaptor2d)
        ---C++: inline
    	returns Real;
	

    Value (myclass; C: Curve2d from Adaptor2d; X: Real)
        ---C++: inline
    	returns Pnt2d from gp;


    D0 (myclass; C: Curve2d from Adaptor2d; U: Real ; 
                 P: out Pnt2d);
        ---C++: inline

    D1 (myclass; C: Curve2d from Adaptor2d; U: Real ; 
                 P: out Pnt2d; T: out Vec2d);
         ---C++: inline

    D2 (myclass; C: Curve2d from Adaptor2d; U: Real ; 
                 P: out Pnt2d; T,N: out Vec2d);
         ---C++: inline
    
    D3 (myclass; C: Curve2d from Adaptor2d; U: Real ; 
                 P: out Pnt2d; T,N,V: out Vec2d);
         ---C++: inline
    
    DN(myclass; C: Curve2d from Adaptor2d; U: Real ; 
                 N: Integer from Standard)
         returns Vec2d;
         ---C++: inline

   NbIntervals(myclass ; C:  Curve2d from Adaptor2d) 
        ---Purpose : output the number of interval of continuity C2 of 
        --           the curve
        ---C++: inline
        returns Integer from Standard;
        
   Intervals         (myclass; C:  Curve2d from Adaptor2d
		       ; Tab    : out    Array1OfReal from TColStd);
	---Purpose: compute Tab. 
        ---C++: inline

   GetInterval (myclass; C:  Curve2d from Adaptor2d
                       ; Index  : Integer from Standard
		       ; Tab    : Array1OfReal from TColStd
    	    	       ; U1, U2 : out Real from Standard);
        ---Purpose : output the bounds of interval of index <Index>
        --           used if Type == Composite.
        ---C++: inline

   Degree(myclass; C : Curve2d from Adaptor2d) returns Integer from Standard;
     	---C++: inline


end Geom2dCurveTool;




