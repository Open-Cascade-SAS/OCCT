-- Created on: 1994-10-03
-- Created by: Christian CAILLET
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ShapeListBinder  from TransferBRep  inherits Binder from Transfer

    ---Purpose : This binder binds several (a list of) shapes with a starting
    --           entity, when this entity itself corresponds to a simple list
    --           of shapes. Each part is not seen as a sub-result of an
    --           independant componant, but as an item of a built-in list

uses CString, Type,
     ShapeEnum from TopAbs,  Shape from TopoDS ,
      Vertex from TopoDS,  Edge  from TopoDS,  Wire  from TopoDS,
      Face   from TopoDS,  Shell from TopoDS,  Solid from TopoDS,
      CompSolid from TopoDS,    Compound from TopoDS ,
      HSequenceOfShape from TopTools

raises TypeMismatch, OutOfRange

is

    Create returns mutable ShapeListBinder;

    Create (list : mutable HSequenceOfShape from TopTools)
    	 returns mutable ShapeListBinder;

    IsMultiple (me) returns Boolean  is redefined;
    -- returns True if more than one result

    ResultType (me) returns Type;
    -- returns TopoDS_Shape

    ResultTypeName (me) returns CString;
    -- returns list(TopoDS_Shape)

    AddResult (me : mutable; res : Shape);
    ---Purpose : Adds an item to the result list

    Result (me) returns HSequenceOfShape from TopTools;

    SetResult (me : mutable; num : Integer; res : Shape);
    ---Purpose : Changes an already defined sub-result

    NbShapes (me) returns Integer;

    Shape (me; num : Integer) returns Shape
    	raises OutOfRange;
    ---C++ : return const &

    ShapeType (me; num : Integer) returns ShapeEnum;

    -- different sub-types for the Result. Shape(num) returns a Shape

    Vertex    (me; num : Integer) returns Vertex    raises TypeMismatch, OutOfRange;
    Edge      (me; num : Integer) returns Edge      raises TypeMismatch, OutOfRange;
    Wire      (me; num : Integer) returns Wire      raises TypeMismatch, OutOfRange;
    Face      (me; num : Integer) returns Face      raises TypeMismatch, OutOfRange;
    Shell     (me; num : Integer) returns Shell     raises TypeMismatch, OutOfRange;
    Solid     (me; num : Integer) returns Solid     raises TypeMismatch, OutOfRange;
    CompSolid (me; num : Integer) returns CompSolid raises TypeMismatch, OutOfRange;
    Compound  (me; num : Integer) returns Compound  raises TypeMismatch, OutOfRange;

fields

    theres :  HSequenceOfShape from TopTools;

end ShapeListBinder;
