-- Created on: 2002-12-12
-- Created by: data exchange team
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class RWCurveElementSectionDerivedDefinitions from RWStepElement

    ---Purpose: Read & Write tool for CurveElementSectionDerivedDefinitions

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    CurveElementSectionDerivedDefinitions from StepElement

is
    Create returns RWCurveElementSectionDerivedDefinitions from RWStepElement;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : CurveElementSectionDerivedDefinitions from StepElement);
	---Purpose: Reads CurveElementSectionDerivedDefinitions

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: CurveElementSectionDerivedDefinitions from StepElement);
	---Purpose: Writes CurveElementSectionDerivedDefinitions

    Share (me; ent : CurveElementSectionDerivedDefinitions from StepElement;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWCurveElementSectionDerivedDefinitions;
