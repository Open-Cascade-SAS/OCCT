-- File:        PrecisionQualifier.cdl
-- Created:     Mon Dec  4 12:02:23 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWPrecisionQualifier from RWStepShape

	---Purpose : Read & Write Module for PrecisionQualifier

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     PrecisionQualifier from StepShape

is

	Create returns RWPrecisionQualifier;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable PrecisionQualifier from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : PrecisionQualifier from StepShape);

end RWPrecisionQualifier;
