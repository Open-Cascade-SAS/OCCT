-- Created on: 2002-12-12
-- Created by: data exchange team
-- Copyright (c) 2002-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class SymmetricTensor22d from StepFEA
inherits SelectType from StepData

    ---Purpose: Representation of STEP SELECT type SymmetricTensor22d

uses
    HArray1OfReal from TColStd

is
    Create returns SymmetricTensor22d from StepFEA;
	---Purpose: Empty constructor

    CaseNum (me; ent: Transient) returns Integer;
	---Purpose: Recognizes a kind of SymmetricTensor22d select type
	--          1 -> HArray1OfReal from TColStd
	--          0 else

    AnisotropicSymmetricTensor22d (me) returns HArray1OfReal from TColStd;
	---Purpose: Returns Value as AnisotropicSymmetricTensor22d (or Null if another type)

end SymmetricTensor22d;
