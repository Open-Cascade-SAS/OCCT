-- Created on: 1997-02-10
-- Created by: Alexander BRIVIN and Dmitry TARASOV
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Material from Vrml inherits  TShared  from  MMgt

	---Purpose: defines a Material node of VRML specifying properties of geometry
	---          and its appearance.
    	--  This node defines the current surface material properties for all subsequent shapes.
        --  Material sets several components of the current material during traversal. Different shapes
        --  interpret materials with multiple values differently. To bind materials to shapes, use a
        --  MaterialBinding node. 

    	--  The lighting parameters defined by the Material node are the same parameters defined by
        --  the OpenGL lighting model. 
uses 
 
    HArray1OfColor  from   Quantity, 
    HArray1OfReal   from   TColStd

is
 
    Create  (  aAmbientColor   :  HArray1OfColor  from   Quantity; 
    	       aDiffuseColor   :  HArray1OfColor  from   Quantity;
    	       aSpecularColor  :  HArray1OfColor  from   Quantity; 
	       aEmissiveColor  :  HArray1OfColor  from   Quantity; 
	       aShininess      :  HArray1OfReal   from   TColStd; 
	       aTransparency   :  HArray1OfReal   from   TColStd ) 
	  returns mutable Material from Vrml; 

    Create  returns mutable Material from Vrml;

    SetAmbientColor  ( me : mutable; aAmbientColor   :  HArray1OfColor  from  Quantity );
    AmbientColor  ( me )  returns  HArray1OfColor  from  Quantity;

    SetDiffuseColor  ( me : mutable; aDiffuseColor   :  HArray1OfColor  from  Quantity );
    DiffuseColor  ( me )  returns  HArray1OfColor  from  Quantity;

    SetSpecularColor ( me : mutable; aSpecularColor  :  HArray1OfColor  from  Quantity );
    SpecularColor ( me )  returns  HArray1OfColor  from  Quantity;

    SetEmissiveColor ( me : mutable; aEmissiveColor  :  HArray1OfColor  from  Quantity );
    EmissiveColor ( me )  returns  HArray1OfColor  from  Quantity;

    SetShininess  ( me : mutable;  aShininess : HArray1OfReal from TColStd  ); 
    Shininess  ( me )  returns  HArray1OfReal from TColStd; 

    SetTransparency  ( me : mutable;
    	    	aTransparency  :  HArray1OfReal from TColStd  ); 
    Transparency  ( me )  returns  HArray1OfReal from TColStd; 

    Print  ( me; anOStream: in out OStream from Standard) returns OStream from Standard;
    ---C++:  return  & 

fields
 
    myAmbientColor   :  HArray1OfColor  from   Quantity;	-- Ambient color
    myDiffuseColor   :  HArray1OfColor  from   Quantity;	-- Diffuse color
    mySpecularColor  :  HArray1OfColor  from   Quantity;	-- Specular color
    myEmissiveColor  :  HArray1OfColor  from   Quantity;	-- Emissive color
    myShininess      :  HArray1OfReal   from   TColStd;	        -- Shininess
    myTransparency   :  HArray1OfReal   from   TColStd;    	-- Transparency

end Material;
