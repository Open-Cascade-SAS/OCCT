-- Created on: 2001-08-24
-- Created by: Alexander GRIGORIEV
-- Copyright (c) 2001-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- modified     13.04.2009 Sergey Zaritchny

class GeometryDriver from BinMDataXtd  inherits ADriver from BinMDF

        ---Purpose: Attribute Driver.

uses
    SRelocationTable from BinObjMgt,
    RRelocationTable from BinObjMgt,
    Persistent       from BinObjMgt,
    MessageDriver    from CDM,
    Attribute        from TDF

is
    Create (theMessageDriver:MessageDriver from CDM)
        returns mutable GeometryDriver from BinMDataXtd;

    NewEmpty (me)  returns mutable Attribute from TDF;

    Paste(me; Source     : Persistent from BinObjMgt;
              Target     : mutable Attribute from TDF;
              RelocTable : out RRelocationTable from BinObjMgt)
        returns Boolean from Standard;

    Paste(me; Source     : Attribute from TDF;
              Target     : in out Persistent from BinObjMgt;
              RelocTable : out SRelocationTable from BinObjMgt);

end GeometryDriver;
