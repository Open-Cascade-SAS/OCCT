-- Created on: 1992-04-06
-- Created by: Christian CAILLET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class DefSwitch  from IGESData  inherits Storable

    ---Purpose : description of a directory componant which can be either
    --           undefined (let Void), defined as a Reference to an entity,
    --           or as a Rank, integer value adressing a builtin table
    --           The entity reference is not included here, only reference
    --           status is kept (because entity type must be adapted)

uses Integer, DefType

is

    Create returns DefSwitch;
    ---Purpose : creates a DefSwitch as Void

    SetVoid (me : in out)  is static;
    ---Purpose : sets DefSwitch to "Void" status (in file : Integer = 0)

    SetReference (me : in out)  is static;
    ---Purpose : sets DefSwitch to "Reference" Status (in file : Integer < 0)

    SetRank (me : in out; val : Integer)  is static;
    ---Purpose : sets DefSwitch to "Rank" with a Value (in file : Integer > 0)

    DefType (me) returns DefType  is static;
    ---Purpose : returns DefType status (Void,Reference,Rank)

    Value (me) returns Integer  is static;
    ---Purpose : returns Value as Integer (sensefull for a Rank)

fields

    theval : Integer;

end DefSwitch;
