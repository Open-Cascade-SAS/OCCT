-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class QuasiUniformCurveAndRationalBSplineCurve from StepGeom 

inherits BSplineCurve from StepGeom 


	--- This classe is an implementation of EXPRESS
	--  ANDOR Subtype Declaration.
uses

	QuasiUniformCurve from StepGeom, 
	RationalBSplineCurve from StepGeom, 
	HAsciiString from TCollection, 
	Integer from Standard, 
	HArray1OfCartesianPoint from StepGeom, 
	BSplineCurveForm from StepGeom, 
	Logical from StepData, 
	HArray1OfReal from TColStd, 
	Real from Standard
is

	Create returns QuasiUniformCurveAndRationalBSplineCurve;
	---Purpose: Returns a QuasiUniformCurveAndRationalBSplineCurve


	Init (me : mutable;
	      aName : HAsciiString from TCollection;
	      aDegree : Integer from Standard;
	      aControlPointsList : HArray1OfCartesianPoint from StepGeom;
	      aCurveForm : BSplineCurveForm from StepGeom;
	      aClosedCurve : Logical from StepData;
	      aSelfIntersect : Logical from StepData) is redefined;

	Init (me : mutable;
	      aName : HAsciiString from TCollection;
	      aDegree : Integer from Standard;
	      aControlPointsList : HArray1OfCartesianPoint from StepGeom;
	      aCurveForm : BSplineCurveForm from StepGeom;
	      aClosedCurve : Logical from StepData;
	      aSelfIntersect : Logical from StepData;
	      aQuasiUniformCurve : QuasiUniformCurve from StepGeom;
	      aRationalBSplineCurve : RationalBSplineCurve from StepGeom) is virtual;

	Init (me : mutable;
	      aName : HAsciiString from TCollection;
	      aDegree : Integer from Standard;
	      aControlPointsList : HArray1OfCartesianPoint from StepGeom;
	      aCurveForm : BSplineCurveForm from StepGeom;
	      aClosedCurve : Logical from StepData;
	      aSelfIntersect : Logical from StepData;
	      aWeightsData : HArray1OfReal from TColStd) is virtual;

	-- Specific Methods for Field Data Access --

	SetQuasiUniformCurve(me : mutable; aQuasiUniformCurve : QuasiUniformCurve);
	QuasiUniformCurve (me) returns QuasiUniformCurve;
	SetRationalBSplineCurve(me : mutable; aRationalBSplineCurve : RationalBSplineCurve);
	RationalBSplineCurve (me) returns RationalBSplineCurve;

	-- Specific Methods for ANDOR Field Data Access --


	-- Specific Methods for ANDOR Field Data Access --

	SetWeightsData(me : mutable; aWeightsData : HArray1OfReal);
	WeightsData (me) returns HArray1OfReal;
	WeightsDataValue (me; num : Integer) returns Real;
	NbWeightsData (me) returns Integer;

fields

	quasiUniformCurve : QuasiUniformCurve from StepGeom;
	rationalBSplineCurve : RationalBSplineCurve from StepGeom;

end QuasiUniformCurveAndRationalBSplineCurve;
