-- Created on: 1992-03-26
-- Created by: Herve LEGRAND
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


package Geom2dLProp

    ---Purpose: Handles local properties of curves and surfaces from the 
    --          packages Geom and Geom2d.
    -- SeeAlso: Package LProp.


    ---Level : Public. 
    --  All methods of all  classes will be public.

uses Standard, gp, Geom2d, LProp

is
    
    class Curve2dTool;
    
    class CLProps2d from Geom2dLProp 
            instantiates CLProps from LProp(Curve         from Geom2d,
	                                    Vec2d         from gp,
					    Pnt2d         from gp,
					    Dir2d         from gp,
					    Curve2dTool   from Geom2dLProp); 
    class CurAndInf2d; 
    
    private class NumericCurInf2d instantiates NumericCurInf from LProp( 
    	    	    	    	    	       Curve         from Geom2d,
	                                       Vec2d         from gp,
					       Pnt2d         from gp,
					       Dir2d         from gp,
					       Curve2dTool   from Geom2dLProp); 
					    
end Geom2dLProp;    




