-- File     : Prs2d_Diameter.cdl
-- Created  : April  2000
-- Author   : Tanya COOL
---Copyright: Matra Datavision 2000

class Diameter from Prs2d inherits Dimension from Prs2d

 ---Purpose: Constructs the primitive Radius

uses

	Drawer		   from Graphic2d,
	GraphicObject	   from Graphic2d,
	Pnt2d              from gp,
	Circ2d             from gp,
	ExtendedString     from TCollection,
	ArrowSide          from Prs2d,
	TypeOfDist         from Prs2d,
	TypeOfArrow        from Prs2d,
        FStream            from Aspect 

raises 

    ConstructionError from Standard

is
	Create( aGraphicObject: GraphicObject  from Graphic2d;
	        anAttachPnt   : Pnt2d          from gp;
            	aCircle       : Circ2d         from gp;
          	aText         : ExtendedString from TCollection;
		aTxtScale     : Real           from Standard = 10.0;
            	anArrAngle    : Real           from Standard = 20.0;
		anArrLength   : Real           from Standard = 25.0;
	    	anArrType     : TypeOfArrow    from Prs2d = Prs2d_TOA_OPENED;
		anArrow       : ArrowSide      from Prs2d = Prs2d_AS_BOTHAR;
            	IsReverseArrow: Boolean        from Standard = Standard_False )

	returns mutable Diameter from Prs2d;

    	---Purpose: Creates the radius of the circle passing through 
    	--          the point <anAttachPnt>

    	--------------------------------------
	-- Category: Inquire methods
	--------------------------------------
    
    Values( me; anAttPnt: out Pnt2d from gp; 
            aCirc: out Circ2d from gp ); 
    	---Level: Internal
    	---Purpose: allows to get the properties of the diameter

    --------------------------
    -- Category: Draw and Pick
    --------------------------

    Draw( me : mutable; aDrawer: Drawer from Graphic2d )
	is static protected;
    	---Level: Internal
    	---Purpose: Draws the angle <me>.

    DrawElement( me : mutable; aDrawer: Drawer from Graphic2d;
                 anIndex: Integer from Standard)
        is redefined protected;
    	---Level: Internal
    	---Purpose: Draws element <anIndex> of the diameter <me>.

    DrawVertex( me : mutable; aDrawer: Drawer from Graphic2d;
                anIndex: Integer from Standard)
        is redefined protected;
    	---Level: Internal
    	---Purpose: Draws vertex <anIndex> of the diameter <me>.

    Pick( me : mutable; X, Y: ShortReal from Standard;
	  aPrecision: ShortReal from Standard;
	  aDrawer: Drawer from Graphic2d)
	returns Boolean from Standard
	is static protected;
    	---Level: Internal
    	---Purpose: Returns Standard_True if the diameter <me> is picked,
    	--	    Standard_False if not.

    Save( me; aFStream: in out FStream from Aspect ) is virtual;

    
    CalcTxtPos(me:mutable; theFromAbs: 
    	        Boolean from Standard=Standard_False) 
    	---C++: inline
    	is redefined protected;	
    
fields
 
	myX1   : ShortReal  from Standard;
	myY1   : ShortReal  from Standard;
	myX2   : ShortReal  from Standard;
	myY2   : ShortReal  from Standard;
    	myPnt  : Pnt2d      from gp;
        myCirc : Circ2d     from gp;
--enk fields. Coordinates of appendix. 
	myAppX1   : ShortReal  from Standard;
	myAppY1   : ShortReal  from Standard;
	myAppX2   : ShortReal  from Standard;
	myAppY2   : ShortReal  from Standard;
    	myInside  : Boolean    from Standard;
end Diameter from Prs2d;
