-- Created on: 1993-06-03
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



generic class SurfFunction from Contap 
    (TheSurface as any;
     TheSurfaceTool as any;
     TheSurfProps   as any; -- as SurfProps from Contap(TheSurface,
                            --                          TheSurfaceTool)
     TheContTool    as any)

inherits FunctionSetWithDerivatives from math			       
    
	---Purpose: This class describes the function on a parametric surface.
	--          the form of the function is F(u,v) = 0 where u and v are
	--          the parameteric coordinates of a point on the surface,
	--          to compute the contours of the surface.

uses Vector    from math,
     Matrix    from math,
     Pnt       from gp,
     Vec       from gp,
     Dir       from gp,
     Dir2d     from gp,
     TFunction from Contap


raises UndefinedDerivative from StdFail

is

    Create
    
    	returns SurfFunction from Contap;


    Set(me: in out; S: TheSurface)

    	is static;


    Set(me: in out; Eye: Pnt from gp)
    
    	---C++: inline
    	is static;


    Set(me: in out; Dir: Dir from gp)
    
    	---C++: inline
    	is static;


    Set(me: in out; Dir: Dir from gp; Angle: Real from Standard)
    
    	---C++: inline
    	is static;


    Set(me: in out; Eye: Pnt from gp; Angle: Real from Standard)
    
    	---C++: inline
    	is static;


    Set(me: in out; Tolerance: Real from Standard)
    
    	---C++: inline
    	is static;


    NbVariables(me)

	---Purpose: This method has to return 2.
    	returns Integer from Standard;


    NbEquations(me)

	---Purpose: This method has to return 1.
    	returns Integer from Standard;


    Value(me : in out; X : Vector from math;
                       F : out Vector from math)

	---Purpose: The dimension of F is 1.

    	returns Boolean from Standard;


    Derivatives(me : in out; X : Vector from math;
                             D : out Matrix from math)

	---Purpose: The dimension of D is (1,2).

    	returns Boolean from Standard;


    Values(me : in out; X : Vector from math;
                        F : out Vector from math;
                        D : out Matrix from math)

    	returns Boolean from Standard;


    Root(me)

	---Purpose: Root is the value of the function at the solution.
	--          It is a vector of dimension 1, i-e a real.

    	returns Real from Standard
	---C++: inline
    	is static;


    Tolerance(me)
    
	---Purpose: Returns the value Tol so that if Abs(Func.Root())<Tol
	--          the function is considered null.
	--          
	---C++: inline
    
    	returns Real from Standard
	is static;


    Point(me)

	---Purpose: Returns the value of the solution point on the surface.

    	returns Pnt from gp
	---C++: return const&
	---C++: inline
    	is static;
    

    IsTangent(me : in out)

    	returns Boolean from Standard 
    	is static;
    

    Direction3d(me: in out)

    	returns Vec from gp
	---C++: return const&
	---C++: inline
    	raises UndefinedDerivative from StdFail
    	is static;
    

    Direction2d(me: in out)

    	returns Dir2d from gp
	---C++: return const&
	---C++: inline
    	raises UndefinedDerivative from StdFail
    	is static;


    FunctionType(me)
    
    	returns TFunction from Contap
	---C++: inline
	is static;


    Eye(me)
    
    	returns Pnt from gp
	---C++: return const&
	---C++: inline
	is static;


    Direction(me)
    
    	returns Dir from gp
	---C++: return const&
	---C++: inline
	is static;


    Angle(me)
    
    	returns Real from Standard
	---C++: inline
	is static;


    Surface(me)
    
    	returns any TheSurface
	---C++: return const&
	---C++: inline
	is static;
	


fields

    mySurf   : TheSurface;
    myMean   : Real      from Standard;
    myType   : TFunction from Contap;
    myDir    : Dir       from gp;
    myEye    : Pnt       from gp;
    myAng    : Real      from Standard;
    myCosAng : Real      from Standard;
    tol      : Real      from Standard;

    solpt  : Pnt   from gp;
    valf   : Real  from Standard;
    Usol   : Real  from Standard;
    Vsol   : Real  from Standard;
    Fpu    : Real  from Standard;
    Fpv    : Real  from Standard;
    d2d    : Dir2d from gp;
    d3d    : Vec   from gp;
    
    tangent   : Boolean from Standard;
    computed  : Boolean from Standard;
    derived   : Boolean from Standard;

end SurfFunction;
