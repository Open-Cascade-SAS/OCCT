-- File:	C2d2TanRad.cdl
-- Created:	Tue Oct 20 16:23:30 1992
-- Author:	Remi GILET
--		<reg@sdsun1>
---Copyright:	 Matra Datavision 1992

class Circ2d2TanRad from Geom2dGcc

	---Purpose: This class implements the algorithms used to 
	--          create 2d circles tangent to one curve and a
	--          point/line/circle/curv and with a given radius.
    	--          For each construction methods arguments are:
    	--            - Two Qualified elements for tangency constrains.
    	--            (for example EnclosedCirc if we want the 
    	--            solution inside the argument EnclosedCirc).
    	--            - Two Reals. One (Radius) for the radius and the 
    	--            other (Tolerance) for the tolerance.
    	--          Tolerance is only used for the limit cases.
    	--          For example : 
    	--          We want to create a circle inside a circle C1 and 
    	--          inside a curve Cu2 with a radius Radius and a 
    	--          tolerance Tolerance.
    	--          If we did not used Tolerance it is impossible to 
    	--          find a solution in the the following case : Cu2 is 
    	--          inside C1 and there is no intersection point 
    	--          between the two elements.
    	--          with Tolerance we will give a solution if the 
    	--          lowest distance between C1 and Cu2 is lower than or 
    	--          equal Tolerance.

-- inherits Entity from Standard

uses QualifiedCurve   from Geom2dGcc,
     Integer          from Standard,
     Boolean          from Standard,
     Pnt2d            from gp,
     Point            from Geom2d,
     Circ2d           from gp,
     Array1OfPnt2d    from TColgp,
     Array1OfCirc2d   from TColgp,
     Array1OfInteger  from TColStd,
     Array1OfReal     from TColStd,
     Circ2d2TanRad    from GccAna,
     MyCirc2d2TanRad  from Geom2dGcc,
     Position         from GccEnt,
     Array1OfPosition from GccEnt
     
raises OutOfRange    from Standard,
       BadQualifier  from GccEnt,
       NotDone       from StdFail,
       NegativeValue from Standard

is

Create(Qualified1 : QualifiedCurve from Geom2dGcc ;
       Qualified2 : QualifiedCurve from Geom2dGcc ;
       Radius     : Real           from Standard  ;
       Tolerance  : Real           from Standard  ) 
returns Circ2d2TanRad from Geom2dGcc
raises BadQualifier, NegativeValue;

Create(Qualified1 : QualifiedCurve from Geom2dGcc ;
       Point      : Point          from Geom2d    ;
       Radius     : Real           from Standard  ;
       Tolerance  : Real           from Standard  ) 
returns Circ2d2TanRad from Geom2dGcc
raises BadQualifier, NegativeValue;

Create(Point1     : Point          from Geom2d    ;
       Point2     : Point          from Geom2d    ;
       Radius     : Real           from Standard  ;
       Tolerance  : Real           from Standard  ) 
returns Circ2d2TanRad from Geom2dGcc
raises NegativeValue;

    	---Purpose: These constructors create one or more 2D circles of radius Radius either
    	-- -   tangential to the 2 curves Qualified1 and Qualified2,   or
    	-- -   tangential to the curve Qualified1 and passing through the point Point, or
    	-- -   passing through two points Point1 and Point2.
    	-- Tolerance is a tolerance criterion used by the algorithm
    	-- to find a solution when, mathematically, the problem
    	-- posed does not have a solution, but where there is
    	-- numeric uncertainty attached to the arguments.
    	-- For example, take two circles C1 and C2, such that C2
    	-- is inside C1, and almost tangential to C1. There is, in
    	-- fact, no point of intersection between C1 and C2. You
    	-- now want to find a circle of radius R (smaller than the
    	-- radius of C2), which is tangential to C1 and C2, and
    	-- inside these two circles: a pure mathematical resolution
    	-- will not find a solution. This is where the tolerance
    	-- criterion is used: the algorithm considers that C1 and
    	-- C2 are tangential if the shortest distance between these
    	-- two circles is less than or equal to Tolerance. Thus, a
    	-- solution is found by the algorithm.
    	-- Exceptions
    	-- GccEnt_BadQualifier if a qualifier is inconsistent with
    	-- the argument it qualifies (for example, enclosing for a line).
    	-- Standard_NegativeValue if Radius is negative.


Results(me   : in out                         ;
    	Circ :        Circ2d2TanRad from GccAna)
is static;

Results(me   : in out                              ;
    	Circ :        MyCirc2d2TanRad from Geom2dGcc)
is static;

IsDone(me) returns Boolean from Standard
is static;
    	---Purpose: This method returns True if the algorithm succeeded.
    	-- Note: IsDone protects against a failure arising from a
    	-- more internal intersection algorithm, which has reached its numeric limits.

NbSolutions(me) returns Integer from Standard
raises NotDone
is static;
    	---Purpose: This method returns the number of solutions.
    	--          NotDone is raised if the algorithm failed.
    	-- Exceptions
    	-- StdFail_NotDone if the construction fails.
    
ThisSolution(me ; Index : Integer from Standard) returns Circ2d from gp 
raises OutOfRange, NotDone
is static;
    	---Purpose: Returns the solution number Index and raises OutOfRange 
    	-- exception if Index is greater than the number of solutions.
    	-- Be carefull: the Index is only a way to get all the 
    	-- solutions, but is not associated to theses outside the context of the algorithm-object.
    	-- Warning
    	-- This indexing simply provides a means of consulting the
    	-- solutions. The index values are not associated with
    	-- these solutions outside the context of the algorithm object.
    	-- Exceptions
    	-- Standard_OutOfRange if Index is less than zero or
    	-- greater than the number of solutions computed by this algorithm.
    	-- StdFail_NotDone if the construction fails.    

WhichQualifier(me                                  ;
    	       Index   :     Integer  from Standard;
	       Qualif1 : out Position from GccEnt  ;
	       Qualif2 : out Position from GccEnt  )
raises OutOfRange, NotDone
is static;
    	---Purpose: Returns the qualifiers Qualif1 and Qualif2 of the
    	-- tangency arguments for the solution of index Index
    	-- computed by this algorithm.
    	-- The returned qualifiers are:
    	-- -   those specified at the start of construction when the
    	--   solutions are defined as enclosed, enclosing or
    	--   outside with respect to the arguments, or
    	-- -   those computed during construction (i.e. enclosed,
    	--   enclosing or outside) when the solutions are defined
    	--   as unqualified with respect to the arguments, or
    	-- -   GccEnt_noqualifier if the tangency argument is a point, or
    	-- -   GccEnt_unqualified in certain limit cases where it
    	--   is impossible to qualify the solution as enclosed, enclosing or outside.
    	-- Exceptions
    	-- Standard_OutOfRange if Index is less than zero or
    	-- greater than the number of solutions computed by this algorithm.
    	-- StdFail_NotDone if the construction fails.
        
Tangency1(me                                     ;
          Index         : Integer   from Standard;
          ParSol,ParArg : out Real  from Standard;
          PntSol        : out Pnt2d from gp      )
raises OutOfRange, NotDone
is static;
    	---Purpose: Returns informations about the tangency point between the 
    	-- result number Index and the first argument.
    	-- ParSol is the intrinsic parameter of the point PntSol on the solution curv.
    	-- ParArg is the intrinsic parameter of the point PntSol on the argument curv.
    	-- OutOfRange is raised if Index is greater than the number of solutions.
    	-- notDone is raised if the construction algorithm did not succeed.

Tangency2(me                                     ;
          Index         : Integer   from Standard;
          ParSol,ParArg : out Real  from Standard;
          PntSol        : out Pnt2d from gp      )
raises OutOfRange, NotDone
is static;
    	---Purpose: Returns informations about the tangency point between the 
    	-- result number Index and the second argument.
    	-- ParSol is the intrinsic parameter of the point PntSol on the solution curv.
    	-- ParArg is the intrinsic parameter of the point PntSol on the argument curv.
    	-- OutOfRange is raised if Index is greater than the number of solutions.
    	-- notDone is raised if the construction algorithm did not succeed.

IsTheSame1(me                            ;
           Index : Integer  from Standard) returns Boolean from Standard
raises OutOfRange, NotDone
is static;
    	---Purpose: Returns true if the solution of index Index and,
    	-- respectively, the first or second argument of this
    	-- algorithm are the same (i.e. there are 2 identical circles).
    	-- If Rarg is the radius of the first or second argument,
    	-- Rsol is the radius of the solution and dist is the
    	-- distance between the two centers, we consider the two
    	-- circles to be identical if |Rarg - Rsol| and dist
    	-- are less than or equal to the tolerance criterion given at
    	-- the time of construction of this algorithm.
    	-- OutOfRange is raised if Index is greater than the number of solutions.
    	-- notDone is raised if the construction algorithm did not succeed.

IsTheSame2(me                            ;
           Index : Integer from Standard ) returns Boolean from Standard
raises OutOfRange, NotDone
is static;
      	---Purpose: Returns true if the solution of index Index and,
    	-- respectively, the first or second argument of this
    	-- algorithm are the same (i.e. there are 2 identical circles).
    	-- If Rarg is the radius of the first or second argument,
    	-- Rsol is the radius of the solution and dist is the
    	-- distance between the two centers, we consider the two
    	-- circles to be identical if |Rarg - Rsol| and dist
    	-- are less than or equal to the tolerance criterion given at
    	-- the time of construction of this algorithm.
    	-- OutOfRange is raised if Index is greater than the number of solutions.
    	-- notDone is raised if the construction algorithm did not succeed.

fields

    WellDone : Boolean from Standard;
    	---Purpose: Returns True if the algorithm succeeded.

    cirsol   : Array1OfCirc2d from TColgp;
    	---Purpose: TheSolution.

    NbrSol   : Integer from Standard;
    	---Purpose: Returns the number of solutions.

    qualifier1 : Array1OfPosition from GccEnt;
    	---Purpose: The qualifiers of the first argument.

    qualifier2 : Array1OfPosition from GccEnt;
    	---Purpose: The qualifiers of the second argument.

    TheSame1 : Array1OfInteger from TColStd;
    	---Purpose: Returns 1 if the solution and the first argument are the same (2 circles).
    	-- if R1 is the radius of the first argument and Rsol the radius 
    	-- of the solution and dist the distance between the two centers,
	-- we concider the two circles are identical if R1+dist-Rsol is less than Tolerance.
    	-- 0 in the other cases.

    TheSame2 : Array1OfInteger from TColStd;
    	---Purpose: 1 if the solution and the second argument are the same (2 circles).
    	-- if R2 is the radius of the second argument and Rsol the radius 
    	-- of the solution and dist the distance between the two centers,
    	-- we concider the two circles are identical if R2+dist-Rsol is less than Tolerance.
    	-- 0 in the other cases.

    pnttg1sol   : Array1OfPnt2d from TColgp;
    	---Purpose: The tangency point between the solution and the first argument on the solution.

    pnttg2sol   : Array1OfPnt2d from TColgp;
    	---Purpose: The tangency point between the solution and the second argument on the solution.

    par1sol   : Array1OfReal from TColStd;
    	---Purpose: The parameter of the tangency point between the solution and the first argument on the solution.

    par2sol   : Array1OfReal from TColStd;
    	---Purpose: The parameter of the tangency point between the solution and the second argument on the solution.

    pararg1   : Array1OfReal from TColStd;
    	---Purpose: The parameter of the tangency point between the solution and the first argument on the first argument.

    pararg2   : Array1OfReal from TColStd;
    	---Purpose: The parameter of the tangency point between the solution and the second argument on the second argument.

    Invert   : Boolean from Standard;
    
--    CircAna  : Circ2d2TanRad from GccAna;
--    CircGeo  : MyrCirc2d2TanRad from Geom2dGcc;
--    TypeAna  : Boolean;

end Circ2d2TanRad;

