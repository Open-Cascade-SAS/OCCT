-- Created on: 1993-09-07
-- Created by: Bruno DUMORTIER
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class ComputeApprox from ProjLib 


uses
     HCurve       from Adaptor3d,
     HSurface     from Adaptor3d,
     BSplineCurve from Geom2d,
     BezierCurve  from Geom2d
is

    Create(C   : HCurve   from Adaptor3d ; 
           S   : HSurface from Adaptor3d;
    	   Tol : Real     from Standard) 
    	---Purpose: <Tol>    is   the   tolerance   with  which    the
    	--          approximation is performed.
    returns ComputeApprox from ProjLib;
    
    BSpline(me) returns BSplineCurve from Geom2d ;

    Bezier(me)  returns BezierCurve  from Geom2d ;
    
    Tolerance(me) returns Real from Standard;
    	---Purpose: returns the reached Tolerance.
    
fields

    myTolerance : Real         from Standard;    
    myBSpline   : BSplineCurve from Geom2d ;
    myBezier    : BezierCurve  from Geom2d ;

end ComputeApprox;
