-- File:        PersonAndOrganizationRole.cdl
-- Created:     Mon Dec  4 12:02:28 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWPersonAndOrganizationRole from RWStepBasic

	---Purpose : Read & Write Module for PersonAndOrganizationRole

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     PersonAndOrganizationRole from StepBasic

is

	Create returns RWPersonAndOrganizationRole;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable PersonAndOrganizationRole from StepBasic);

	WriteStep (me; SW : in out StepWriter; ent : PersonAndOrganizationRole from StepBasic);

end RWPersonAndOrganizationRole;
