-- Created on: 1995-03-29
-- Created by: Frederic MAUPAS
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class TranslateEdgeLoop from StepToTopoDS
    inherits Root from StepToTopoDS
    
    ---Purpose:
    --         

uses

    FaceBound              from StepShape,
    Surface                from StepGeom,
    Tool                   from StepToTopoDS,
    TranslateEdgeLoopError from StepToTopoDS,
    Shape                  from TopoDS,
    Surface                from Geom,
    Face                   from TopoDS,
    NMTool                 from StepToTopoDS
    
raises NotDone from StdFail

is

    Create returns TranslateEdgeLoop;
    
    Create (FB     : FaceBound     from StepShape;
            F      : Face          from TopoDS;
            S      : Surface       from Geom;
            SS     : Surface       from StepGeom;
            ss     : Boolean       from Standard;
            T      : in out Tool   from StepToTopoDS;
            NMTool : in out NMTool from StepToTopoDS)
    	returns TranslateEdgeLoop;
	    
    Init (me     : in out;
          FB     : FaceBound     from StepShape;
          F      : Face          from TopoDS;
          S      : Surface       from Geom;
          SS     : Surface       from StepGeom;
          ss     : Boolean       from Standard;
          T      : in out Tool   from StepToTopoDS;
          NMTool : in out NMTool from StepToTopoDS);

    Value (me) returns Shape from TopoDS
    	raises NotDone
	is static;
	---C++: return const &

    Error (me) returns TranslateEdgeLoopError from StepToTopoDS;
    
fields

    myError  : TranslateEdgeLoopError  from StepToTopoDS;
    
    myResult : Shape               from TopoDS;
    
end TranslateEdgeLoop;
