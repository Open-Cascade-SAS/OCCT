-- Created on: 1997-11-06
-- Created by: Roman BORISOV
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

private  class PrjFunc from ProjLib inherits  FunctionSetWithDerivatives from math

	---Purpose: 

uses   
    Vector from math,  
    Matrix from math, 
    CurvePtr  from  Adaptor3d,
    SurfacePtr  from  Adaptor3d,
    Pnt2d  from  gp 

raises  ConstructionError

is
    Create  (C: CurvePtr  from  Adaptor3d; FixVal:  Real  from  Standard;  S:  SurfacePtr  from  Adaptor3d; Fix: Integer)   
    returns  PrjFunc 
    raises  ConstructionError;

    NbVariables(me)
    	---Purpose: returns the number of variables of the function.

    returns Integer;
    
    NbEquations(me)
    	---Purpose: returns the number of equations of the function.

    returns Integer;
    
    Value(me: in out; X: Vector  from  math; F: out Vector  from  math)
    	---Purpose: computes the values <F> of the Functions for the 
    	--          variable <X>.
    	--          Returns True if the computation was done successfully, 
    	--          False otherwise.

    returns Boolean;
    
    Derivatives(me: in out; X: Vector  from  math; D: out Matrix  from  math)
    	---Purpose: returns the values <D> of the derivatives for the 
    	--          variable <X>.
    	--          Returns True if the computation was done successfully, 
    	--          False otherwise.

    returns Boolean;
    
    Values(me: in out; X: Vector  from  math; F: out Vector  from  math; D: out Matrix  from  math)
    	---Purpose: returns the values <F> of the functions and the derivatives
    	--          <D> for the variable <X>.
    	--          Returns True if the computation was done successfully, 
    	--          False otherwise.

    returns Boolean;
  
    Solution(me)  returns  Pnt2d  from  gp; 
    	---Purpose:  returns  point  on  surface

fields 

    myCurve      :  CurvePtr    from  Adaptor3d; 
    mySurface    :  SurfacePtr  from  Adaptor3d; 
    myt          :  Real        from  Standard;
    myU,  myV    :  Real        from  Standard;	
    myFix        :  Integer     from  Standard; 
    myNorm       :  Real        from  Standard;     
end PrjFunc;
