-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class RationalBSplineCurve from StepGeom 

inherits BSplineCurve from StepGeom 

uses

	HArray1OfReal from TColStd, 
	Real from Standard, 
	HAsciiString from TCollection, 
	Integer from Standard, 
	HArray1OfCartesianPoint from StepGeom, 
	BSplineCurveForm from StepGeom, 
	Logical from StepData
is

	Create returns mutable RationalBSplineCurve;
	---Purpose: Returns a RationalBSplineCurve


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aDegree : Integer from Standard;
	      aControlPointsList : mutable HArray1OfCartesianPoint from StepGeom;
	      aCurveForm : BSplineCurveForm from StepGeom;
	      aClosedCurve : Logical from StepData;
	      aSelfIntersect : Logical from StepData) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aDegree : Integer from Standard;
	      aControlPointsList : mutable HArray1OfCartesianPoint from StepGeom;
	      aCurveForm : BSplineCurveForm from StepGeom;
	      aClosedCurve : Logical from StepData;
	      aSelfIntersect : Logical from StepData;
	      aWeightsData : mutable HArray1OfReal from TColStd) is virtual;

	-- Specific Methods for Field Data Access --

	SetWeightsData(me : mutable; aWeightsData : mutable HArray1OfReal);
	WeightsData (me) returns mutable HArray1OfReal;
	WeightsDataValue (me; num : Integer) returns Real;
	NbWeightsData (me) returns Integer;

fields

	weightsData : HArray1OfReal from TColStd;

end RationalBSplineCurve;
