-- Created on: 1997-04-21
-- Created by: Prestataire Mary FABIEN
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Filter from TopOpeBRepDS 

---Purpose: 

uses

    Shape       from TopoDS,
    Edge        from TopoDS,
    ListOfShape from TopTools,
    IndexedMapOfShape from TopTools,
    
    Config                           from TopOpeBRepDS,    
    Interference                     from TopOpeBRepDS,
    ListOfInterference               from TopOpeBRepDS,
    ListIteratorOfListOfInterference from TopOpeBRepDS,
    ListOfShapeOn1State from TopOpeBRepDS,
    DataMapOfShapeListOfShapeOn1State from TopOpeBRepDS,
    HDataStructure from TopOpeBRepDS,
    PShapeClassifier from TopOpeBRepTool

is

    Create(HDS : HDataStructure from TopOpeBRepDS;
           pClassif: PShapeClassifier from TopOpeBRepTool = 0) returns Filter;

    ProcessInterferences(me : in out); -- oldies
    
    ProcessFaceInterferences(me : in out;
    	    	    	     MEsp : DataMapOfShapeListOfShapeOn1State from TopOpeBRepDS);
    ProcessFaceInterferences(me : in out; I : Integer;
	    		     MEsp : DataMapOfShapeListOfShapeOn1State from TopOpeBRepDS);

    ProcessEdgeInterferences(me : in out);
    ProcessEdgeInterferences(me : in out; I : Integer);

    ProcessCurveInterferences(me: in out);
    ProcessCurveInterferences(me: in out; I : Integer);


fields

    myHDS : HDataStructure from TopOpeBRepDS;
    myPShapeClassif: PShapeClassifier from TopOpeBRepTool;
    
end Filter from TopOpeBRepDS;
