-- Created on: 1993-06-17
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class PaveClassifier from TopOpeBRepBuild 
    inherits LoopClassifier from TopOpeBRepBuild 

---Purpose: 
-- This class compares vertices on an edge. 
-- 
-- A vertex V1 is inside a vertex V2 if V1 is on the
-- part of the curve defined by V2.
-- 
-- If V2 is FORWARD V1 must be after V2 on the curve.
-- If V2 is REVERSED V1 must be before V2 on the curve.
-- If V2 is INTERNAL V1 is always inside.
-- If V2 is EXTERNAL V1 is never inside.

uses

    ShapeEnum from TopAbs,
    State from TopAbs,
    Shape from TopoDS,
    Edge from TopoDS,
    Orientation from TopAbs,
    Loop from TopOpeBRepBuild
    
is

    Create(E : Shape from TopoDS) returns PaveClassifier;
    ---Purpose: Create a Pave classifier to compare vertices on edge <E>.

    Compare(me : in out; L1,L2 : Loop from TopOpeBRepBuild)  
    returns State from TopAbs;
    ---Purpose: Returns state of vertex <L1> compared with <L2>.

    SetFirstParameter(me : in out; P : Real from Standard) 
    is static;
    ClosedVertices(me : in out; B : Boolean from Standard)
    is static;

    AdjustCase(myclass;p1:Real;o:Orientation;
    	    	       first,period:Real;tol:Real;
    	    	       cas:out Integer) returns Real;

    CompareOnNonPeriodic(me : in out) returns State from TopAbs 
    is static private;
    CompareOnPeriodic(me : in out) returns State from TopAbs 
    is static private;
    AdjustOnPeriodic(me : in out) 
    is static private;
    ToAdjustOnPeriodic(me) returns Boolean from Standard 
    is static private;

fields

    myEdge : Edge from TopoDS;
    myEdgePeriodic : Boolean from Standard;
    myFirst  : Real from Standard;
    myPeriod : Real from Standard;
    mySameParameters : Boolean from Standard;
    myClosedVertices : Boolean from Standard;

    myP1 : Real from Standard;
    myP2 : Real from Standard;
    myO1 : Orientation from TopAbs;
    myO2 : Orientation from TopAbs;

    myCas1 : Integer from Standard;  -- debug
    myCas2 : Integer from Standard;  -- debug

end PaveClassifier from TopOpeBRepBuild;
