-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Organization from StepBasic 

inherits TShared from MMgt

uses

	HAsciiString from TCollection, 
	Boolean from Standard
is

	Create returns mutable Organization;
	---Purpose: Returns a Organization

	Init (me : mutable;
	      hasAid : Boolean from Standard;
	      aId : mutable HAsciiString from TCollection;
	      aName : mutable HAsciiString from TCollection;
	      aDescription : mutable HAsciiString from TCollection) is virtual;

	-- Specific Methods for Field Data Access --

	SetId(me : mutable; aId : mutable HAsciiString);
	UnSetId (me:mutable);
	Id (me) returns mutable HAsciiString;
	HasId (me) returns Boolean;
	SetName(me : mutable; aName : mutable HAsciiString);
	Name (me) returns mutable HAsciiString;
	SetDescription(me : mutable; aDescription : mutable HAsciiString);
	Description (me) returns mutable HAsciiString;

fields

	id : HAsciiString from TCollection;   -- OPTIONAL can be NULL
	name : HAsciiString from TCollection;
	description : HAsciiString from TCollection;
	hasId : Boolean from Standard;

end Organization;
