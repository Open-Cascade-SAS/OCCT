-- File:	IGESAppli_ToolFlow.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolFlow  from IGESAppli

    ---Purpose : Tool to work on a Flow. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses Flow from IGESAppli,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolFlow;
    ---Purpose : Returns a ToolFlow, ready to work


    ReadOwnParams (me; ent : mutable Flow;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : Flow;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : Flow;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a Flow <ent>, from
    --           its specific (own) parameters

    OwnCorrect (me; ent : mutable Flow) returns Boolean  is static;
    ---Purpose : Sets automatic unambiguous Correction on a Flow
    --           (NbContextFlags forced to 2)

    DirChecker (me; ent : Flow) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : Flow;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : Flow; entto : mutable Flow;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : Flow;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolFlow;
