-- Created on: 1995-03-03
-- Created by: Jean-Louis Frenkel
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


private class RectangularGraphicGrid from V2d inherits Primitive from Graphic2d


uses
	Drawer          from Graphic2d,
	GraphicObject	from Graphic2d,
	Length          from Quantity,
        GridDrawMode    from Aspect,
	FStream         from Aspect 
is

	Create (aGraphicObject: GraphicObject from Graphic2d;
		X, Y, alpha, beta, xo ,yo: Real from Standard;
                aTenthColorIndex: Integer from Standard)
	returns mutable RectangularGraphicGrid from V2d;

	SetDrawMode(me: mutable; aDrawMode: GridDrawMode from Aspect)
	is static;
	
	Draw (me: mutable; aDrawer: Drawer from Graphic2d)
	is redefined static protected;
	---Level: Internal
	---Purpose: Draws the grid

	Pick (me: mutable; X, Y: ShortReal from Standard;
		aPrecision: ShortReal from Standard;
		aDrawer: Drawer from Graphic2d)
	returns Boolean from Standard is redefined static protected;
	---Level: Internal
	---Purpose: Returns Standard_True if the infinite line <me> is picked,
	--	    Standard_False if not.

        DrawNetwork(me; aDrawer: Drawer from Graphic2d; 
                        alpha,step:ShortReal from Standard;
                        xfrom,yfrom, sizefrom: ShortReal from Standard )
	is static private;

        DrawPoints(me;  aDrawer: Drawer from Graphic2d; 
                        xfrom,yfrom, sizefrom: ShortReal from Standard )
	is static private;

	Save( me; aFStream: in out FStream from Aspect ) is virtual;

fields
	StepX, StepY,a1,a2,OX,OY: ShortReal from Standard;
        DrawMode: GridDrawMode from Aspect;
	myTenthColorIndex: Integer from Standard;
end RectangularGraphicGrid from V2d;

