-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class OrientedPath from StepShape 

inherits Path from StepShape 

uses

	Boolean from Standard, 
	HArray1OfOrientedEdge from StepShape, 
	OrientedEdge from StepShape, 
	HAsciiString from TCollection,
	EdgeLoop from StepShape
is

	Create returns OrientedPath;
	---Purpose: Returns a OrientedPath


	Init (me : mutable;
	      aName : HAsciiString from TCollection;
	      aEdgeList : HArray1OfOrientedEdge from StepShape) is redefined;

	Init (me : mutable;
	      aName : HAsciiString from TCollection;
	      aPathElement : EdgeLoop from StepShape;
	      aOrientation : Boolean from Standard) is virtual;

	-- Specific Methods for Field Data Access --

	SetPathElement(me : mutable; aPathElement : EdgeLoop);
	PathElement (me) returns EdgeLoop;
	SetOrientation(me : mutable; aOrientation : Boolean);
	Orientation (me) returns Boolean;
	SetEdgeList(me : mutable; aEdgeList : HArray1OfOrientedEdge) is redefined;
	EdgeList (me) returns HArray1OfOrientedEdge is redefined;
	EdgeListValue (me; num : Integer) returns OrientedEdge is redefined;
	NbEdgeList (me) returns Integer is redefined;

fields

	pathElement : EdgeLoop from StepShape;
	orientation : Boolean from Standard;

 -- 
 -- NB : field <edge_list> inherited from classe <EdgeLoop> is redeclared.
 --      it shall appears in a physical file as a *.
 --

end OrientedPath;
