-- Created by: Peter KURNEV
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


package BOPAlgo 
---Purpose: 

uses
    gp, 
    TopAbs, 
    Geom,  
    GeomAPI, 
    BRepClass3d,
    TopoDS, 
    TopTools, 
    IntTools,
    IntSurf,
    --
    BOPDS, 
    BOPInt, 
    BOPCol, 
    BOPTools 
is   
    enumeration Operation is  
      COMMON, 
      FUSE, 
      CUT,    
      CUT21,
      SECTION, 
      UNKNOWN
    end Operation;   
     
    enumeration CheckStatus is
      CheckUnknown,
      BadType,
      SelfIntersect,
      TooSmallEdge,
      NonRecoverableFace,
      IncompatibilityOfVertex,
      IncompatibilityOfEdge,
      IncompatibilityOfFace, 
      OperationAborted,
      NotValid
    end CheckStatus;

    --
    -- classes 
    --   
    deferred class Algo; 
    deferred class BuilderShape; 
    class PaveFiller;
    class Builder; 
    class BOP; 
    --	
    deferred class BuilderArea;
    class BuilderFace;
    class WireEdgeSet;
    class WireSplitter; 
    class BuilderSolid; 
    class Tools; 
    class SectionAttribute; 
    class CheckerSI; 
    class ArgumentAnalyzer; 
    class CheckResult;
    --
    --  pointers
    --
    pointer PPaveFiller to PaveFiller from BOPAlgo; 
    pointer PWireEdgeSet to WireEdgeSet from BOPAlgo; 
    pointer PBOP to BOP from BOPAlgo;  
    pointer PBuilder to Builder from BOPAlgo;  
    pointer PArgumentAnalyzer to ArgumentAnalyzer from BOPAlgo;  
    -- 
    imported ListOfCheckResult; 
    
end BOPAlgo;
