-- File:	IntStart_ArcTool.cdl
-- Created:	Tue May  4 18:01:10 1993
-- Author:	Jacques GOUSSARD
--		<jag@topsn2>
---Copyright:	 Matra Datavision 1993


deferred generic class ArcTool from IntStart
    (TheArc as any )


    ---Purpose: Template class for a tool on the restriction of
    --          a surface.
    -- It is possible to implement this class with an instantiation
    -- of the class CurveTool from Adaptor3d..


is


    Resolution(myclass; A: TheArc; Tol3d: Real from Standard)

        ---Purpose :  Returns the parametric resolution corresponding
        --         to the space resolution Tol3d.

    	returns Real from Standard;


end ArcTool;



