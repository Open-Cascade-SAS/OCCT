-- Created on: 1993-06-14
-- Created by: Martine LANGLOIS
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class MakeAxis2Placement3d from GeomToStep inherits Root from GeomToStep

    ---Purpose: This class implements the mapping between classes 
    --          Axis2Placement from Geom and Ax2, Ax3 from gp, and the class
    --          Axis2Placement3d from StepGeom which describes an
    --          axis2_placement_3d from Prostep. 
   
uses Ax2 from gp,
     Ax3 from gp,
     Trsf from gp,
     Axis2Placement from Geom,
     Axis2Placement3d from StepGeom
     
raises NotDone from StdFail
     
is 

Create returns MakeAxis2Placement3d;
-- creates an identity (original axis)

Create ( A : Ax2 from gp ) returns MakeAxis2Placement3d;

Create ( A : Ax3 from gp ) returns MakeAxis2Placement3d;

Create ( T : Trsf from gp) returns MakeAxis2Placement3d;

Create ( A : Axis2Placement from Geom ) returns MakeAxis2Placement3d;

Value (me) returns Axis2Placement3d from StepGeom
    raises NotDone
    is static;
    ---C++: return const&

fields

    theAxis2Placement3d : Axis2Placement3d from StepGeom;
    	-- TheOP solution from StepGeom
    	
end MakeAxis2Placement3d;


