-- Created on: 2004-02-04
-- Created by: Sergey KUUL
-- Copyright (c) 2004-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class SplitCommonVertex from ShapeFix inherits Root from ShapeFix

	---Purpose: Two wires have common vertex - this case is valid in BRep model
        --          and isn't valid in STEP => before writing into STEP it is necessary
        --          to split this vertex (each wire must has one vertex)

uses
    Shape from TopoDS
    
is
    Create returns SplitCommonVertex;
    ---Purpose :

    Init(me: mutable; S : Shape from TopoDS); 
    ---Purpose :
    
    Perform(me:mutable);	
    ---Purpose :
    
    Shape(me : mutable) returns Shape from TopoDS;
    ---Purpose :

fields

    myShape    : Shape from TopoDS;
    myResult   : Shape from TopoDS;
    myStatus   : Integer; -- error status

end SplitCommonVertex;
