-- Created on: 1993-02-03
-- Created by: Gilles DEBARBOUILLE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class RealParameter from Dynamic

inherits

    Parameter from Dynamic
	---Purpose: This  inherited class from Parameter describes all
	--          the parameters, which  are characterized by a real
	--          value.

uses

    OStream from Standard,
    CString from Standard,
    Real    from Standard


is

    Create(aparameter : CString from Standard )
    
    ---Level: Public 
    
    ---Purpose: Creates a RealParameter with <aparameter> as name.
    
    returns mutable RealParameter from Dynamic;

    Create(aparameter : CString from Standard ; avalue : Real from Standard) 
    
    ---Level: Public 
    
    ---Purpose: With  the name  of the Parameter  <aparameter> and the
    --          real <avalue>, creates an instance of RealParameter.
    
    returns mutable RealParameter from Dynamic;
    
    Value(me) returns Real from Standard
    
    ---Level: Public 
    
    ---Purpose: Returns the value of the parameter which is a real.
    
    is static;

    Value (me : mutable ; avalue : Real from Standard)
    
    ---Level: Public 
    
    --- Purpose: Sets the real <avalue> in <me>.

    is static;
    
    Dump(me ; astream : in out OStream from Standard)
    
    ---Level: Internal 
    
    ---Purpose: Useful for debugging.

    is redefined;
    
fields

    thevalue : Real from Standard;

end RealParameter;
