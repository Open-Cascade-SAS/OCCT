-- Created on: 1996-12-16
-- Created by: Christian CAILLET
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SelectInt  from StepData    inherits SelectMember

    ---Purpose : A SelectInt is a SelectMember specialised for a basic integer
    --           type in a select which also accepts entities : this one has
    --           NO NAME.
    --           For a named select, see SelectNamed

uses CString, Logical

is

    Create returns SelectInt;

    Kind (me) returns Integer  is redefined;
    --  possible kind for Int : integer boolean logical enum(without text)

    SetKind  (me : mutable; kind : Integer)  is redefined;
    --  called by various Set*

    Int  (me) returns Integer  is redefined;

    SetInt (me : mutable; val : Integer)  is redefined;

fields

    thekind : Integer;
    theval  : Integer;

end SelectInt;
