-- Created on: 2008-01-20
-- Created by: Alexander A. BORODIN
-- Copyright (c) 2008-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


-- Updated:       


class FontMgr from OSD inherits TShared from MMgt

 ---Purpose: Structure for store of Font System Information

uses Path,
     SystemFont,
     NListOfSystemFont,
     AsciiString from TCollection
is
 GetInstance(myclass)
    returns FontMgr;
    ---Level: Public

 GetAvalableFonts(me)
    returns NListOfSystemFont;

--- Private methods

 Create returns FontMgr is private;
    ---Purpose: Creates empty font object
    ---Level: Private

 InitFontDataBase(me:mutable) is private;

fields

 MyListOfFonts:         NListOfSystemFont;

end FontMgr;