-- Created on: 1993-06-17
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class CurveIterator from TopOpeBRepDS 
    inherits InterferenceIterator from TopOpeBRepDS

uses

    State         from TopAbs,
    Orientation   from TopAbs,
    Interference  from TopOpeBRepDS,
    ListOfInterference  from TopOpeBRepDS,
    Curve         from Geom2d
    
is
    Create(L : ListOfInterference from TopOpeBRepDS) returns CurveIterator; 
    ---Purpose: Creates an  iterator on the  curves on surface
    --          described by the interferences in <L>.
    
    MatchInterference(me; I : Interference from TopOpeBRepDS) 
    returns Boolean from Standard
    ---Purpose: Returns  True if the Interference <I>  has a 
    --          GeometryType() TopOpeBRepDS_CURVE
    --          returns False else.
    is redefined;

    Current(me) returns Integer from Standard
    ---Purpose: Index of the curve in the data structure.
    is static;
    
    Orientation(me; S : State from TopAbs) returns Orientation from TopAbs
    is static;
    
    PCurve(me) returns Curve from Geom2d
    ---C++: return const &
    is static;
    
end CurveIterator from TopOpeBRepDS;
