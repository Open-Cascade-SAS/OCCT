-- Created on: 1994-10-07
-- Created by: Yves FRICAUD
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class LinkTopoBilo from BRepMAT2d 

	---Purpose:Constucts links between the Face of the explorer and
    	--         the BasicElts contained in the bisecting locus. 

uses
    Shape                            from TopoDS,
    Wire                             from TopoDS,	    
    Explorer                         from BRepMAT2d,
    DataMapOfShapeSequenceOfBasicElt from BRepMAT2d,
    DataMapOfBasicEltShape           from BRepMAT2d,
    BisectingLocus                   from BRepMAT2d,
    BasicElt                         from MAT

raises
    ConstructionError from Standard
    
is

    Create  returns LinkTopoBilo from BRepMAT2d;    

    Create( Explo : Explorer       from BRepMAT2d; 
    	    BiLo  : BisectingLocus from BRepMAT2d)	
    returns LinkTopoBilo from BRepMAT2d    
	---Purpose: Constructs the links Between S and BiLo.
	--          
    raises
    	ConstructionError from Standard;
	---Purpose: raises if <S> is not a face.
    
    
    Perform( me    : in out; 
	     Explo : Explorer       from BRepMAT2d; 
    	     BiLo  : BisectingLocus from BRepMAT2d)  
    	---Purpose: Constructs the links Between S and BiLo.
 	--     
    raises
    	ConstructionError from Standard
	---Purpose: raises if <S> is not a face or a wire.         
    is static;
    
    
    Init (me : in out; S : Shape from TopoDS)
    	---Purpose: Initialise the Iterator on <S>
    	--          <S> is an edge or a vertex of the initial
    	--          wire or face.
    raises
    	ConstructionError from Standard
	---Purpose: raises if <S> is not an edge or a vertex.
    is static;
    
    
    More (me : in out)	returns Boolean from Standard
    	---Purpose: Returns True if there  is a current  BasicElt.
    is static;
    
    
    Next (me : in out)    	
    	---Purpose: Proceed to the next BasicElt.
    is static;
    
    
    Value(me) returns BasicElt from MAT	
    	---Purpose: Returns the current BasicElt.
    is static;
    
    GeneratingShape (me ; aBE : BasicElt from MAT)
	---Purpose: Returns the Shape linked to <aBE>.
    returns Shape from TopoDS
    is static;
    
    LinkToWire (me           : in out; 
    	        W            : Wire           from TopoDS;
		Explo        : Explorer       from BRepMAT2d;    
                IndexContour : Integer        from Standard;
                BiLo         : BisectingLocus from BRepMAT2d) 
    is static private;
    

fields
    myMap      : DataMapOfShapeSequenceOfBasicElt from BRepMAT2d;
    myBEShape  : DataMapOfBasicEltShape           from BRepMAT2d;
    myKey      : Shape                            from TopoDS;
    current    : Integer                          from Standard; 
    isEmpty    : Boolean                          from Standard;
    
end ;



