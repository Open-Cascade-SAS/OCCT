-- Created on: 1992-08-13
-- Created by: Remi LEQUETTE
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




package TopBas 

	---Purpose: The  TopBas package  provides  data structure  for
	--          topological algorithms.   THe data  structures are
	--          used to store the intermediary dat and the results
	--          of the algorithms.
	--          
	--          *  Interference, List  :  An Interference  is  the
	--          topological    representation  of an intersection.
	--          The classes are generic in order to be independant
	--          of the data structure.

uses
    Standard,
    TCollection,
    TopAbs

is
    generic class Interference;
	---Purpose: The   Interference  is  the    description  of  an
	--          intersection on a Shape.

    class TestInterference instantiates Interference from TopBas
    	    	    	    (Real    from Standard,
    	    	    	     Integer from Standard);
			    
    class ListOfTestInterference instantiates 
    List from TCollection (TestInterference);

end TopBas;


