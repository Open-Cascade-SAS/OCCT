-- File:	StepDimTol_DatumReference.cdl
-- Created:	Wed Jun  4 13:34:35 2003 
-- Author:	Galina KULIKOVA
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class DatumReference from StepDimTol
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity DatumReference

uses
    Datum from StepDimTol

is
    Create returns DatumReference from StepDimTol;
	---Purpose: Empty constructor

    Init (me: mutable; aPrecedence: Integer;
                       aReferencedDatum: Datum from StepDimTol);
	---Purpose: Initialize all fields (own and inherited)

    Precedence (me) returns Integer;
	---Purpose: Returns field Precedence
    SetPrecedence (me: mutable; Precedence: Integer);
	---Purpose: Set field Precedence

    ReferencedDatum (me) returns Datum from StepDimTol;
	---Purpose: Returns field ReferencedDatum
    SetReferencedDatum (me: mutable; ReferencedDatum: Datum from StepDimTol);
	---Purpose: Set field ReferencedDatum

fields
    thePrecedence: Integer;
    theReferencedDatum: Datum from StepDimTol;

end DatumReference;
