-- Created on: 1997-08-26
-- Created by: SMO
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




package MPrsStd 

	---Purpose: Storage    and  Retrieval  drivers   for graphic
	--          attributes.   Transient  attributes are defined in
	--          package TPrsStd and persistent one are defined in
	--          package PPrsStd

uses TDF,
     PDF,
     MDF, 
     CDM

is

    	    ---Purpose: Storage drivers for graphic attributes from
    	    --          TPrsStd
    	    ---Category: StorageDriver

	class AISPresentationStorageDriver;
	class PositionStorageDriver;
	
    	    ---Purpose: Retrieval drivers for graphic attributes from
    	    --          PPrsStd
    	    ---Category: RetrievalDriver


        class AISPresentationRetrievalDriver;
        class AISPresentationRetrievalDriver_1;	
	class PositionRetrievalDriver;
	
    AddStorageDrivers(aDriverTable : ASDriverHSequence from MDF;theMessageDriver : MessageDriver from CDM);
	---Purpose: Adds the attribute storage drivers to <aDriverTable>.
    	---Category: StorageDriversTable


    AddRetrievalDrivers(aDriverTable : ARDriverHSequence from MDF;theMessageDriver : MessageDriver from CDM);
	---Purpose: Adds the attribute retrieval drivers to <aDriverTable>.
    	---Category: RetrievalDriversTable


end MPrsStd;



