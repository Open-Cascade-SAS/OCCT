-- Created on: 1991-02-27
-- Created by: Jean Claude Vauthier
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class UniformAbscissa from GCPnts 
  

    ---Purpose: This class allows to compute a uniform distribution of points
    --          on a curve (ie the points will all be equally distant).
uses 
    Curve        from Adaptor3d,
    Curve2d      from Adaptor2d,
    HArray1OfReal from TColStd

    
raises DomainError       from Standard, 
       ConstructionError from Standard,
       OutOfRange        from Standard,
       NotDone           from StdFail

is
        
    Create 
    	---Purpose: creation of a indefinite UniformAbscissa
    	returns UniformAbscissa from GCPnts;

    Create(C : in out Curve from Adaptor3d ; Abscissa : Real ; Toler : Real = -1)
        --- Purpose : Computes a uniform abscissa distribution of points on 
        --  the Curve <C>. Parameter Toler is equal Precision::Confusion by default.
	--  It Is used for more precise calculation of curve length
    	returns UniformAbscissa from GCPnts
     	raises ConstructionError;

    Create(C : in out Curve from Adaptor3d ; Abscissa, U1, U2 : Real ; 
               Toler : Real = -1)
        --- Purpose : Computes a Uniform abscissa distribution of points 
        --  on a part of the Curve <C>. Parameter Toler is equal Precision::Confusion by default.
	--  It Is used for more precise calculation of curve length
     	returns UniformAbscissa from GCPnts
     	raises ConstructionError,
               DomainError;

    Create(C : in out Curve from Adaptor3d ; NbPoints : Integer ; 
           Toler : Real = -1)
        --- Purpose : Computes a uniform abscissa distribution of points on 
        --  the Curve <C>. 
        --  <NbPoints> defines the nomber of desired points. 
	--  Parameter Toler is equal Precision::Confusion by default.
	--  It Is used for more precise calculation of curve length
    	returns UniformAbscissa from GCPnts
     	raises ConstructionError,
               DomainError;

    Create(C : in out Curve from Adaptor3d ; NbPoints : Integer; U1, U2 : Real ; 
           Toler : Real = -1)
        --- Purpose : Computes a Uniform abscissa distribution of points 
        --  on a part of the Curve <C>. 
	--  Parameter Toler is equal Precision::Confusion by default.
	--  It Is used for more precise calculation of curve length
     	returns UniformAbscissa from GCPnts
     	raises ConstructionError,
               DomainError;

    Initialize(me : in out; C : in out Curve from Adaptor3d ; Abscissa : Real ;
                            Toler : Real = -1)
    	---Purpose: Initialize the algoritms with <C>, <Abscissa>, <Toler>
     	raises ConstructionError
	is static;

    Initialize(me : in out; C : in out Curve from Adaptor3d ; Abscissa, U1, U2 : Real ; 
                            Toler : Real = -1)
    	---Purpose: Initialize the algoritms with <C>, <Abscissa>, <U1>,
    	--          <U2>, <Toler>
     	raises ConstructionError,
               DomainError
	is static;

  
    Initialize(me : in out; C : in out Curve from Adaptor3d ; NbPoints : Integer ; 
                            Toler : Real = -1)
    	---Purpose: Initialize the algoritms with <C>, <NbPoints>, <Toler> and 
     	raises ConstructionError
	is static;


    Initialize(me : in out; C : in out Curve from Adaptor3d ; NbPoints : Integer; U1, U2 : Real ; 
                            Toler : Real = -1)
    	---Purpose: Initialize the algoritms with <C>, <Abscissa>, <U1>,
    	--          <U2>, <Toler>.
     	raises ConstructionError,
               DomainError
	is static;

    Create(C : in out Curve2d from Adaptor2d ; Abscissa : Real ; Toler : Real = -1)
        --- Purpose : Computes a uniform abscissa distribution of points on 
        --  the Curve2d <C>. 
        --  Parameter Toler is equal Precision::Confusion by default.
	--  It Is used for more precise calculation of curve length
    	returns UniformAbscissa from GCPnts
     	raises ConstructionError;

    Create(C : in out Curve2d from Adaptor2d ; Abscissa, U1, U2 : Real ; Toler : Real = -1)
        --- Purpose : Computes a Uniform abscissa distribution of points 
        --  on a part of the Curve2d <C>. 
	--  Parameter Toler is equal Precision::Confusion by default.
	--  It Is used for more precise calculation of curve length
     	returns UniformAbscissa from GCPnts
     	raises ConstructionError,
               DomainError;

    Create(C : in out Curve2d from Adaptor2d ; NbPoints : Integer ; 
               Toler : Real = -1)
        --- Purpose : Computes a uniform abscissa distribution of points on 
        --  the Curve2d <C>. 
        --  <NbPoints> defines the nomber of desired points. 
	--  Parameter Toler is equal Precision::Confusion by default.
	--  It Is used for more precise calculation of curve length
    	returns UniformAbscissa from GCPnts
     	raises ConstructionError,
               DomainError;

    Create(C : in out Curve2d from Adaptor2d ; NbPoints : Integer; U1, U2 : Real ; 
               Toler : Real = -1)
        --- Purpose : Computes a Uniform abscissa distribution of points 
        --  on a part of the Curve2d <C>. 
	--  Parameter Toler is equal Precision::Confusion by default.
	--  It Is used for more precise calculation of curve length
     	returns UniformAbscissa from GCPnts
     	raises ConstructionError,
               DomainError;

    Initialize(me : in out; C : in out Curve2d from Adaptor2d ; Abscissa : Real ; Toler : Real = -1)
    	---Purpose: Initialize the algoritms with <C>, <Abscissa>, <Toler>
     	raises ConstructionError
	is static;

    Initialize(me : in out; C : in out Curve2d from Adaptor2d ; Abscissa, U1, U2 : Real ; 
                            Toler : Real = -1)
    	---Purpose: Initialize the algoritms with <C>, <Abscissa>, <U1>,
    	--          <U2>, <Toler>
     	raises ConstructionError,
               DomainError
	is static;

  
    Initialize(me : in out; C : in out Curve2d from Adaptor2d ; NbPoints : Integer ; 
                            Toler : Real = -1)
    	---Purpose: Initialize the algoritms with <C>, <NbPoints>, <Toler> and 
     	raises ConstructionError
	is static;


    Initialize(me : in out; C : in out Curve2d from Adaptor2d ; NbPoints : Integer; U1, U2 : Real ;
                            Toler : Real = -1)
    	---Purpose: Initialize the algoritms with <C>, <Abscissa>, <U1>,
    	--          <U2>, <Toler>.
     	raises ConstructionError,
               DomainError
	is static;

	       
    IsDone(me) returns Boolean 
	---C++: inline
    	is static;

	       
    NbPoints(me) returns Integer
	---C++: inline
    	 is static;
  
    Parameter(me; Index : Integer) returns Real 
        ---Purpose : returns the computed Parameter of index <Index>.
	---C++: inline
    	is static;
   
    Abscissa(me) returns Real
      	---Purpose : returne the current abscissa
      	-- ie the distance between two consecutive points
	---C++: inline
	is static;

fields

    myDone       : Boolean;
    myNbPoints   : Integer ;
    -- stores the number of points computed with the 
    -- requested Abscissa else stores the requested
    -- number of points 
    myAbscissa   : Real;
    myParams     : HArray1OfReal from TColStd ;
    -- the size of this array will be be bigger than myNbPoints
    --  by one or two 
    
    

end UniformAbscissa;
