-- Created on: 1994-08-31
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class EdgeInfo from Draft

	---Purpose: 

uses Curve   from Geom,
     Curve   from Geom2d,
     Pnt     from gp,
     Face    from TopoDS

raises DomainError from Standard

is


    Create
    
    	returns EdgeInfo from Draft;


    Create(HasNewGeometry: Boolean from Standard)
    
    	returns EdgeInfo from Draft;


    Add(me: in out; F: Face from TopoDS)
    
    	is static;


    RootFace(me: in out; F: Face from TopoDS)
    
    	is static;


    Tangent(me: in out; P: Pnt from gp)
    
    	is static;


    IsTangent(me; P: out Pnt from gp)
    
    	returns Boolean from Standard
	is static;


    NewGeometry(me)
    
    	returns Boolean from Standard
	is static;

    SetNewGeometry(me: in out; NewGeom : Boolean from Standard)
    
	is static;


    Geometry(me)

    	returns Curve from Geom
	is static;
	---C++: return const&


    FirstFace(me)
    
    	returns Face from TopoDS
	is static;
	 ---C++: return const&


    SecondFace(me)
    
    	returns Face from TopoDS
	is static;
	 ---C++: return const&

    FirstPC(me)
    
    	returns Curve from Geom2d
	is static;
	 ---C++: return const&


    SecondPC(me)
    
    	returns Curve from Geom2d
	is static;
	 ---C++: return const&


    ChangeGeometry(me: in out)
    
    	returns Curve from Geom
	is static;
	---C++: return &


    ChangeFirstPC(me: in out)
    
    	returns Curve from Geom2d
	is static;
	---C++: return &


    ChangeSecondPC(me: in out)
    
    	returns Curve from Geom2d
	is static;
	---C++: return &


    RootFace(me)
    
	---C++: return const&
    	returns Face from TopoDS
	is static;

    Tolerance(me: in out; tol: Real from Standard)
	is static;

    Tolerance(me)
    
    	returns Real from Standard
	is static;

fields

    myNewGeom : Boolean from Standard;
    myGeom    : Curve   from Geom;
    myFirstF  : Face    from TopoDS;
    mySeconF  : Face    from TopoDS;
    myFirstPC : Curve   from Geom2d;
    mySeconPC : Curve   from Geom2d;
    myRootFace: Face    from TopoDS;
    myTgt     : Boolean from Standard;
    myPt      : Pnt     from gp;
    myTol     : Real    from Standard;

end EdgeInfo;




