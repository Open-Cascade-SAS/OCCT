-- Created on: 1993-01-09
-- Created by: CKY / Contract Toubro-Larsen ( Arun MENON )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class BasicDimension from IGESDimen   inherits IGESEntity
     
    ---Purpose: Defines IGES Basic Dimension, Type 406, Form 31,
    --          in package IGESDimen
    --          The basic Dimension Property indicates that the referencing 
    --          dimension entity is to be displayed with a box around text. 

uses

        Pnt2d       from gp,
        XY          from gp

is

        Create returns mutable BasicDimension;

            -- --specific-- --

        Init(me                    : mutable; 
             nbPropVal             : Integer;
             lowerLeft, lowerRight : XY;
             upperRight, upperLeft : XY); 
        -- This method is used to set the fields of the
        -- class BasicDimension
        --       - nbPropVal  : Number of property values
        --       - lowerLeft  : Coordinates of lower left corner
        --       - lowerRight : Coordinates of lower right corner
        --       - upperRight : Coordinates of upper right corner
        --       - upperLeft  : Coordinates of upper left corner

        NbPropertyValues(me) returns Integer;
        ---Purpose : returns the number of properties = 8

        LowerLeft(me) returns Pnt2d;
        ---Purpose : returns coordinates of lower left corner

        LowerRight(me) returns Pnt2d;
        ---Purpose : returns coordinates of lower right corner

        UpperRight(me) returns Pnt2d;
        ---Purpose : returns coordinates of upper right corner

        UpperLeft(me) returns Pnt2d;
        ---Purpose : returns coordinates of upper left corner

fields

--
-- Class    : IGESDimen_BasicDimension
-- 
-- Purpose  : Declaration of variables specific to the definition
--            of the Class BasicDimension.
--
-- Reminder : A BasicDimension instance is defined by :
--                - The number of property values, always 8
--                - Coordinates of lower left corner
--                - Coordinates of lower right corner
--                - Coordinates of upper right corner
--                - Coordinates of upper left corner
--
--

        theNbPropertyValues : Integer;
        theLowerLeft        : XY;
        theLowerRight       : XY;
        theUpperRight       : XY;
        theUpperLeft        : XY;

end BasicDimension;
