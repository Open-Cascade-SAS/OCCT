-- Created on: 1993-02-05
-- Created by: Gilles DEBARBOUILLE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DynamicDerivedClass from Dynamic 


inherits

    DynamicClass from Dynamic
    
	---Purpose: The object of  this class is  to allow, as in  the
	--          C++ language,    the  possibility  to   define   a
	--          DynamicDerivedClass  which  inherits from   one or
	--          more DynamicClass.

uses

    CString from Standard,
    Method            from Dynamic,
    DynamicInstance   from Dynamic,
    SequenceOfClasses from Dynamic

is

    Create(aname : CString from Standard) returns mutable DynamicDerivedClass from Dynamic;
    
    ---Level: Public 
    
    ---Purpose: Creates a new instance of this class with <aname> as name.
    
    AddClass(me : mutable ; aclass : any DynamicClass from Dynamic)
    
    ---Level: Public 
    
    ---Purpose: Adds another class <aclass> to the sequence of derived
    --          classes.
    
    is static;
    
    Method(me ; amethod : CString from Standard) returns any Method from Dynamic
    
    ---Level: Public 
    
    ---Purpose: Starting with  the name of  a method,  this  redefined
    --          method searches for   the  right method object  in the
    --          sequence of methods  of  the derived class and  in all
    --          the inherited classes.

    is redefined;
    
    Instance(me) returns mutable DynamicInstance from Dynamic
    
    ---Level: Public 
    
    ---Purpose: Defines an instance of this class definition.

    is redefined;

fields

    thesequenceofclasses : SequenceOfClasses from Dynamic;

end DynamicDerivedClass;
