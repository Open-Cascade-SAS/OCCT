-- Created on: 1993-10-29
-- Created by: Christophe MARION
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PolyHidingData from HLRAlgo
  ---Purpose: Data structure of a set of Hiding Triangles.

uses
    Address from Standard,
    Integer from Standard,
    Real    from Standard

is
    Create returns PolyHidingData from HLRAlgo;
    	---C++: inline

    Set(me : in  out;
	Index,Minim,Maxim : Integer from Standard;
	A,B,C,D           : Real    from Standard)
    	---C++: inline
    is static;
    
    IndexAndMinMax(me) returns Address from Standard
    	---C++: inline
    is static;
    
    Plan(me) returns Address from Standard
    	---C++: inline
    is static;
    
fields
    myMinMax : Integer from Standard[3];
    myPlan   : Real    from Standard[4];
end PolyHidingData;
