-- Created on: 1993-01-09
-- Created by: CKY / Contract Toubro-Larsen ( Anand NATRAJAN )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ExternalRefFileIndex from IGESBasic  inherits IGESEntity

        ---Purpose: defines ExternalRefFileIndex, Type <402> Form <12>
        --          in package IGESBasic
        --          Contains a list of the symbolic names used by the
        --          referencing files and the DE pointers to the
        --          corresponding definitions within the referenced file

uses

        HAsciiString from TCollection,
        HArray1OfHAsciiString     from Interface,
        HArray1OfIGESEntity from IGESData

raises DimensionMismatch, OutOfRange

is

        Create returns mutable ExternalRefFileIndex;

        -- Specific Methods pertaining to the class

        Init (me : mutable; aNameArray : HArray1OfHAsciiString;
              allEntities : HArray1OfIGESEntity)
        raises DimensionMismatch;
        ---Purpose : This method is used to set the fields of the class
        --           ExternalRefFileIndex
        --       - aNameArray  : External Reference Entity symbolic names
        --       - allEntities : External Reference Entities
        -- raises exception if array lengths are not equal
        -- if size of aNameArray is not equal to size of allEntities

        NbEntries (me) returns Integer;
        ---Purpose : returns number of index entries

        Name (me; Index : Integer) returns HAsciiString from TCollection
        raises OutOfRange;
        ---Purpose : returns the External Reference Entity symbolic name
        -- raises exception if Index <= 0 or Index > NbEntries()

        Entity (me; Index : Integer) returns IGESEntity
        raises OutOfRange;
        ---Purpose : returns the internal entity
        -- raises exception if Index <= 0 or Index > NbEntries()

fields

--
-- Class    : IGESBasic_ExternalRefFileIndex
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class ExternalRefFileIndex.
--
-- Reminder : A ExternalRefFileIndex instance is defined by :
--            - External Reference Entity symbolic names
--            - External Reference Entities

        theNames    : HArray1OfHAsciiString;
        theEntities : HArray1OfIGESEntity;

end ExternalRefFileIndex;
