-- File:        ProductDefinitionWithAssociatedDocuments.cdl
-- Created:     Mon Dec  4 12:02:29 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWProductDefinitionWithAssociatedDocuments from RWStepBasic

	---Purpose : Read & Write Module for ProductDefinitionWithAssociatedDocuments

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     ProductDefinitionWithAssociatedDocuments from StepBasic,
     EntityIterator from Interface

is

	Create returns RWProductDefinitionWithAssociatedDocuments;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable ProductDefinitionWithAssociatedDocuments from StepBasic);

	WriteStep (me; SW : in out StepWriter; ent : ProductDefinitionWithAssociatedDocuments from StepBasic);

	Share(me; ent : ProductDefinitionWithAssociatedDocuments from StepBasic; iter : in out EntityIterator);

end RWProductDefinitionWithAssociatedDocuments;
