-- Created on: 1998-06-03
-- Created by: data exchange team
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package ShapeBuild 

    ---Purpose: This package provides basic building tools for other packages in ShapeHealing.
    -- These tools are rather internal for ShapeHealing .

uses
    gp,
    Geom,
    Geom2d,
    TopAbs,
    TopLoc,
    TopoDS,
    TopTools,
    BRep,
    ShapeExtend,
    BRepTools

is

    class Vertex;
    	---Purpose: Provides low-level functions used for constructing vertices
	
    class Edge;
    	---Purpose: Provides low-level functions used for rebuilding edge
	
    class ReShape;
    	---Purpose: Rebuilds a shape with substitution of some components

    PlaneXOY returns Plane from Geom;
    	---Purpose: Returns a Geom_Surface which is the Plane XOY (Z positive)
    	--          This allows to consider an UV space homologous to a 3D space,
    	--          with this support surface

end ShapeBuild;
