-- Created on: 1997-03-26
-- Created by: Christian CAILLET
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DerivedUnit  from StepBasic    inherits TShared

    ---Purpose : Added from StepBasic Rev2 to Rev4

uses
     DerivedUnitElement from StepBasic,
     HArray1OfDerivedUnitElement from StepBasic

is

    Create returns mutable DerivedUnit;

    Init (me : mutable; elements : HArray1OfDerivedUnitElement from StepBasic);

    SetElements (me : mutable; elements : HArray1OfDerivedUnitElement from StepBasic);
    Elements    (me) returns HArray1OfDerivedUnitElement from StepBasic;
    NbElements  (me) returns Integer;
    ElementsValue (me; num : Integer) returns DerivedUnitElement from StepBasic;

fields

    theElements : HArray1OfDerivedUnitElement from StepBasic;

end DerivedUnit;
