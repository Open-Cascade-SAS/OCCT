-- Created on: 1991-05-13
-- Created by: Laurent Painnot
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class FunctionWithDerivative from math
    	 ---Purpose:
    	 -- This abstract class describes the virtual functions associated with
    	 -- a function of a single variable for which the first derivative is
    	 -- available.

inherits Function

is

    Delete(me:out) is virtual;
    	---C++: alias "Standard_EXPORT virtual ~math_FunctionWithDerivative(){Delete();}"
    
    Value(me: in out; X: Real; F: out Real)
        ---Purpose: Computes the value <F>of the function for the variable <X>.
    	--          Returns True if the calculation were successfully done, 
    	--          False otherwise.

    returns Boolean
    is deferred;
 
    Derivative(me: in out; X: Real; D: out Real)
        ---Purpose: Computes the derivative <D> of the function 
        --          for the variable <X>.
    	--           Returns True if the calculation were successfully done, 
    	--           False otherwise.

    returns Boolean
    is deferred;    

    Values(me: in out; X: Real; F, D: out Real)
    	---Purpose: Computes the value <F> and the derivative <D> of the 
    	--          function for the variable <X>.
    	--          Returns True if the calculation were successfully done,
    	--          False otherwise.

    returns Boolean
    is deferred;
    
end FunctionWithDerivative;
