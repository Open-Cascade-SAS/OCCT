-- Created on: 1992-01-17
-- Created by: GG
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Modified:	GG 23/11/00 Add Display(),Erase(),IsDisplayed() methods


class Plane from V3d

inherits

	TShared
	---Purpose: Defines the services of Plane type objects. Only
	--	    the creation and editing of the functions is dealt
	--	    with here.
	-- Warning: The representation of the clipping plane must be
	--	    calculated by the application by means of Graphic3d.
	--	    Editing of this representation must be coherent with
	--	    respect to the position of the plane.

uses

	View from V3d,
	ClipPlane from Visual3d,
	Structure from Graphic3d,
	Parameter from Quantity,
	Color from Quantity


raises

        BadValue from V3d

is

        --
        -- The methods :
        --

	Create (A: Parameter = 0.0;
	        B: Parameter = 0.0;
	        C: Parameter = 1.0;
	        D: Parameter = 0.0
	)  returns mutable Plane
	---Level : Public
        ---Purpose: Creates a clipping plane using the equation :
        --          <A>*X + <B>*Y + <C>*Z + <D> = 0.0
	raises BadValue from V3d;
	---Purpose:  Warning! raises BadValue from V3d
	--          if the norm of the plane is NULL.

        --------------------------------------------------------
        ---Category: Methods to modify the Attributs of the Plane
        --------------------------------------------------------

	SetPlane( me : mutable; A,B,C,D : Parameter)
	---Level : Public
	---Purpose: Modifies the plane equation.
	raises BadValue from V3d
	---Purpose:  Warning! raises BadValue from V3d
	--          if the norm of the plane is NULL.
	--	If the norm of the plane is NULL.
        is static;

        Display(me: mutable; aView: View from V3d;
			     aColor: Color from Quantity= Quantity_NOC_GRAY)
	---Level : Public
	---Purpose: Display the plane representation
        --          in the choosen view.
        is virtual;

        Erase(me: mutable) is static;
        ---Level: Public
        ---Purpose: Erase the plane representation.

        ---------------------------------------------------
        ---Category: Inquire methods
        ---------------------------------------------------

	Plane( me ; A,B,C,D : out Parameter )  is static;
	---Level : Public
	---Purpose: Returns the parameters of the plane .

	IsDisplayed( me ) returns Boolean from Standard is static;
	---Level : Public
	---Purpose: Returns TRUE when the plane representation is displayed

        -----------------------------------------
        ---Category: Private or Protected methods
        -----------------------------------------

        Plane( me) returns mutable ClipPlane from Visual3d is static private ;
	---Level : Internal
        ---Purpose: Returns the associated plane from Visual3d.

	Update( me : mutable ) is static private;
	---Level : Internal
	---Purpose: Updates the the plane representation.


fields

	MyPlane:	ClipPlane from Visual3d ;
	MyGraphicStructure:     Structure from Graphic3d is protected;

friends

        SetPlaneOn from class View from V3d ( me : mutable ),
        SetPlaneOn from class View from V3d
                                ( me : mutable ; Plane : Plane from V3d ),
        SetPlaneOff from class View from V3d ( me : mutable ),
        SetPlaneOff from class View from V3d
                                ( me : mutable ; Plane : Plane from V3d )

end Plane;
