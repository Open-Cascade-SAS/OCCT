-- Created on: 1999-11-26
-- Created by: Andrey BETENEV
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0

class CurveBoundedSurface from StepGeom
inherits BoundedSurface from StepGeom

    ---Purpose: Representation of STEP entity CurveBoundedSurface

uses
    HAsciiString from TCollection,
    Surface from StepGeom,
    HArray1OfSurfaceBoundary from StepGeom

is
    Create returns CurveBoundedSurface from StepGeom;
	---Purpose: Empty constructor

    Init (me: mutable; aRepresentationItem_Name: HAsciiString from TCollection;
                       aBasisSurface: Surface from StepGeom;
                       aBoundaries: HArray1OfSurfaceBoundary from StepGeom;
                       aImplicitOuter: Boolean);
	---Purpose: Initialize all fields (own and inherited)

    BasisSurface (me) returns Surface from StepGeom;
	---Purpose: Returns field BasisSurface
    SetBasisSurface (me: mutable; BasisSurface: Surface from StepGeom);
	---Purpose: Set field BasisSurface

    Boundaries (me) returns HArray1OfSurfaceBoundary from StepGeom;
	---Purpose: Returns field Boundaries
    SetBoundaries (me: mutable; Boundaries: HArray1OfSurfaceBoundary from StepGeom);
	---Purpose: Set field Boundaries

    ImplicitOuter (me) returns Boolean;
	---Purpose: Returns field ImplicitOuter
    SetImplicitOuter (me: mutable; ImplicitOuter: Boolean);
	---Purpose: Set field ImplicitOuter

fields
    theBasisSurface: Surface from StepGeom;
    theBoundaries: HArray1OfSurfaceBoundary from StepGeom;
    theImplicitOuter: Boolean;

end CurveBoundedSurface;
