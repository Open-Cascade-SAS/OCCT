-- Created on: 2000-05-10
-- Created by: Andrey BETENEV
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1

class RoleAssociation from StepBasic
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity RoleAssociation

uses
    ObjectRole from StepBasic,
    RoleSelect from StepBasic

is
    Create returns RoleAssociation from StepBasic;
	---Purpose: Empty constructor

    Init (me: mutable; aRole: ObjectRole from StepBasic;
                       aItemWithRole: RoleSelect from StepBasic);
	---Purpose: Initialize all fields (own and inherited)

    Role (me) returns ObjectRole from StepBasic;
	---Purpose: Returns field Role
    SetRole (me: mutable; Role: ObjectRole from StepBasic);
	---Purpose: Set field Role

    ItemWithRole (me) returns RoleSelect from StepBasic;
	---Purpose: Returns field ItemWithRole
    SetItemWithRole (me: mutable; ItemWithRole: RoleSelect from StepBasic);
	---Purpose: Set field ItemWithRole

fields
    theRole: ObjectRole from StepBasic;
    theItemWithRole: RoleSelect from StepBasic;

end RoleAssociation;
