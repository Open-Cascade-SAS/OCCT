-- File:	StepToGeom_MakeCircle.cdl
-- Created:	Mon Jun 14 15:18:28 1993
-- Author:	Martine LANGLOIS
---Copyright:	 Matra Datavision 1993

class MakeCircle from StepToGeom

    ---Purpose: This class implements the mapping between classes 
    --          Circle from StepGeom which describes a circle from
    --          Prostep and Circle from Geom.
  
uses 
     Circle from Geom,
     Circle from StepGeom
     
is 

    Convert ( myclass; SC : Circle from StepGeom;
                       CC : out Circle from Geom )
    returns Boolean from Standard;

end MakeCircle;
