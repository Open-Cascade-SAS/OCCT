-- Created on: 2001-07-06
-- Created by: Michael KLOKOV
-- Copyright (c) 2001-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class BeanBeanIntersector from IntTools

    ---Purpose: The class BeanBeanIntersector computes ranges of parameters on
    ---         the curve of a first bean (part of edge) that bounds the parts of bean which
    ---	        are on the other bean according to tolerance of edges.

uses
    SequenceOfRoots     from IntTools,
    MarkedRangeSet      from IntTools,
    SequenceOfRanges    from IntTools,
    Range               from IntTools,
    ExtCC               from Extrema,
    ProjectPointOnCurve from GeomAPI,
    Edge                from TopoDS,
    Curve               from BRepAdaptor,
    Curve               from Geom


is
    Create returns BeanBeanIntersector from IntTools;
    
    Create(theEdge1: Edge from TopoDS;
    	   theEdge2: Edge from TopoDS)
	   returns BeanBeanIntersector from IntTools;
    	---Purpose: 
    	--- Initializes the algorithm
	---

    Create(theCurve1        : Curve   from BRepAdaptor;
    	   theCurve2        : Curve from BRepAdaptor;
    	   theBeanTolerance1: Real from Standard;
    	   theBeanTolerance2: Real from Standard)
	   returns BeanBeanIntersector from IntTools;
    	---Purpose: 
    	--- Initializes the algorithm
	---

    Create(theCurve1          : Curve   from BRepAdaptor;
    	   theCurve2          : Curve   from BRepAdaptor;
	   theFirstParOnCurve1: Real from Standard;
	   theLastParOnCurve1 : Real from Standard;
    	   theFirstParOnCurve2: Real from Standard;
	   theLastParOnCurve2 : Real from Standard;
    	   theBeanTolerance1  : Real from Standard;
    	   theBeanTolerance2  : Real from Standard)
	   returns BeanBeanIntersector from IntTools;
    	---Purpose: 
    	--- Initializes the algorithm
	---

    Init(me: in out;theEdge1: Edge from TopoDS;
    	            theEdge2: Edge from TopoDS);
    	---Purpose: 
    	--- Initializes the algorithm
	---



    Init(me: in out;theCurve1        : Curve   from BRepAdaptor;
	    	    theCurve2        : Curve from BRepAdaptor;
    	    	    theBeanTolerance1: Real from Standard;
    	    	    theBeanTolerance2: Real from Standard);
    	---Purpose: 
    	--- Initializes the algorithm
	---

    Init(me: in out;theCurve1          : Curve   from BRepAdaptor;
    	    	    theCurve2          : Curve   from BRepAdaptor;
	    	    theFirstParOnCurve1: Real from Standard;
	    	    theLastParOnCurve1 : Real from Standard;
    	    	    theFirstParOnCurve2: Real from Standard;
	    	    theLastParOnCurve2 : Real from Standard;
    	    	    theBeanTolerance1  : Real from Standard;
    	    	    theBeanTolerance2  : Real from Standard);
    	---Purpose: 
    	--- Initializes the algorithm
	---

    SetBeanParameters(me: in out;IsFirstBean       : Boolean from Standard;
    	    	    	    	 theFirstParOnCurve: Real from Standard;
	    	    	    	 theLastParOnCurve : Real from Standard);
    	---Purpose: 
    	--- Sets bounding parameters for first bean if IsFirstBean is true
	--- and for second bean if IsFirstBean is false
	---


    Perform(me: in out);
    	---Purpose: 
    	--- Launches the algorithm
	--- 

    IsDone(me) returns Boolean from Standard;
    	---C++: inline
	---Purpose: 
    	--- Returns true if the computations was successfull
	--- otherwise returns false

    Result(me)
	returns SequenceOfRanges from IntTools;
	---C++: return const &

    Result(me; theResults: out SequenceOfRanges from IntTools);


    -- private

    ComputeRoughIntersection(me: in out)
    	is private;

    FastComputeIntersection(me: in out)
    	returns Boolean from Standard is private;
    
    ComputeUsingExtrema(me: in out; theRange2: Range from IntTools)
    	is private;
    
    ComputeNearRangeBoundaries(me: in out; theRange2: Range from IntTools)
    	is private;
    
    ComputeRangeFromStartPoint(me: in out; ToIncreaseParameter : Boolean from Standard;
    	    	   			   theParameter        : Real from Standard;
					   theIndex            : Integer from Standard;
					   theParameter2       : Real from Standard;
    	    	    	    	    	   theRange2           : Range from IntTools)
    	is private;

    Distance(me: in out; theArg           : Real from Standard;
    	    	    	 theArgOnOtherBean: out Real from Standard)
    	returns Real from Standard
    	is private;

fields

    -- sources    
    myCurve1          : Curve   from BRepAdaptor;
    myCurve2          : Curve   from BRepAdaptor;
    myTrsfCurve1      : Curve from Geom;
    myTrsfCurve2      : Curve from Geom;

    myFirstParameter1 : Real from Standard;
    myLastParameter1  : Real from Standard;
    myFirstParameter2 : Real from Standard;
    myLastParameter2  : Real from Standard;

    myBeanTolerance1  : Real from Standard;
    myBeanTolerance2  : Real from Standard;
    
    myCurveResolution1: Real from Standard;
    myCriteria        : Real from Standard;

    -- tools
    myProjector      : ProjectPointOnCurve from GeomAPI;
    myRangeManager   : MarkedRangeSet from IntTools;    
    myDeflection     : Real from Standard;

    -- results
    myResults        : SequenceOfRanges from IntTools;

    myIsDone         : Boolean from Standard;

end BeanBeanIntersector from IntTools;
