-- Created on: 2000-10-20
-- Created by: Julia DOROVSKIKH
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class MidPointPresentation from DsgPrs

uses
    Presentation from Prs3d,
    Drawer       from Prs3d,
    Pnt   from gp,
    Lin   from gp,
    Circ  from gp,
    Elips from gp,
    Ax2   from gp

is
    Add( myclass; aPresentation: Presentation from Prs3d;
    	    	  aDrawer      : Drawer from Prs3d;
		  theAxe       : Ax2 from gp;
		  MidPoint     : Pnt from gp;
	          Position     : Pnt from gp;
	       	  AttachPoint  : Pnt from gp;
    	    	  first        : Boolean from Standard);
	           ---Purpose: draws the representation of a MidPoint between
	           --          two vertices.

    Add( myclass; aPresentation: Presentation from Prs3d;
    	    	  aDrawer      : Drawer from Prs3d;
		  theAxe       : Ax2 from gp;
		  MidPoint     : Pnt from gp;
		  Position     : Pnt from gp;
	       	  AttachPoint  : Pnt from gp;
	       	  Point1       : Pnt from gp;
		  Point2       : Pnt from gp;
    	    	  first        : Boolean from Standard);
		   ---Purpose: draws the representation of a MidPoint between
		   --          two lines or linear segments.

    Add( myclass; aPresentation: Presentation from Prs3d;
    	    	  aDrawer      : Drawer from Prs3d;
		  aCircle      : Circ from gp;
		  MidPoint     : Pnt from gp;
		  Position     : Pnt from gp;
	       	  AttachPoint  : Pnt from gp;
	       	  Point1       : Pnt from gp;
		  Point2       : Pnt from gp;
    	    	  first        : Boolean from Standard);
		   ---Purpose: draws the representation of a MidPoint between
		   --          two entire circles or two circular arcs.

    Add( myclass; aPresentation: Presentation from Prs3d;
    	    	  aDrawer      : Drawer from Prs3d;
		  anElips      : Elips from gp;
		  MidPoint     : Pnt from gp;
		  Position     : Pnt from gp;
	       	  AttachPoint  : Pnt from gp;
	       	  Point1       : Pnt from gp;
		  Point2       : Pnt from gp;
    	    	  first        : Boolean from Standard);
		   ---Purpose: draws the representation of a MidPoint between
		   --          two entire ellipses or two elliptic arcs.

end MidPointPresentation;
