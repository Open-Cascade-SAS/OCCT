-- Created on: 2003-12-11
-- Created by: Alexander SOLOVYOV
-- Copyright (c) 2003-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class DeformedDataSource from MeshVS inherits DataSource from MeshVS

	---Purpose: The class provides default class which helps to represent node displacements by deformed mesh
        --    This class has an internal handle to canonical non-deformed mesh data source and
        -- map of displacement vectors. The displacement can be magnified to useful size.
        -- All methods is implemented with calling the corresponding methods of non-deformed data source.

uses
  Integer from Standard,
  Real    from Standard,
  Boolean from Standard,
  Address from Standard,

  Vec from gp,

  Array1OfReal               from TColStd,
  Array1OfInteger            from TColStd,
  PackedMapOfInteger         from TColStd,

  DataMapOfIntegerVector     from MeshVS,
  EntityType                 from MeshVS,
  HArray1OfSequenceOfInteger from MeshVS

is

  Create ( theNonDeformDS : DataSource from MeshVS;
           theMagnify     : Real ) returns mutable DeformedDataSource from MeshVS;
	---Purpose:  Constructor
        -- theNonDeformDS is canonical non-deformed data source, by which we are able to calculate
        --   deformed mesh geometry
        -- theMagnify is coefficient of displacement magnify

  GetGeom ( me; ID     : Integer;
            IsElement  : Boolean;
            Coords     : out Array1OfReal from TColStd;
            NbNodes    : out Integer;
            Type       : out EntityType from MeshVS ) returns Boolean is redefined;

  GetGeomType ( me; ID     : Integer;
                IsElement  : Boolean;
                Type       : out EntityType from MeshVS ) returns Boolean is redefined;

  Get3DGeom( me; ID      : Integer;
                 NbNodes : out Integer;
                 Data    : out HArray1OfSequenceOfInteger from MeshVS ) returns Boolean is redefined;

  GetAddr ( me; ID     : Integer;
            IsElement  : Boolean   ) returns Address is redefined;

  GetNodesByElement ( me; ID  : Integer;
		      NodeIDs : out Array1OfInteger from TColStd;
		      NbNodes : out Integer ) returns Boolean is redefined;

  GetAllNodes    ( me ) returns PackedMapOfInteger from TColStd is redefined;
	---C++: return const &

  GetAllElements ( me ) returns PackedMapOfInteger from TColStd is redefined;
	---C++: return const &

  GetVectors ( me ) returns DataMapOfIntegerVector from MeshVS;
	---C++: return const &
	---Purpose: This method returns map of nodal displacement vectors

  SetVectors ( me: mutable; Map : DataMapOfIntegerVector from MeshVS );
	---Purpose: This method sets map of nodal displacement vectors (Map).

  GetVector  ( me;          ID  : Integer; Vect : out Vec from gp ) returns Boolean;
	---Purpose: This method returns vector ( Vect ) assigned to node number ID.

  SetVector  ( me: mutable; ID  : Integer; Vect :     Vec from gp );
	---Purpose: This method sets vector ( Vect ) assigned to node number ID.

  SetNonDeformedDataSource ( me: mutable; theDS : DataSource from MeshVS );
  GetNonDeformedDataSource    ( me ) returns DataSource from MeshVS;
	---Purpose: With this methods you can read and change internal canonical data source

  SetMagnify ( me: mutable; theMagnify : Real );
  GetMagnify ( me ) returns Real;
	---Purpose: With this methods you can read and change magnify coefficient of nodal displacements

fields
  myNonDeformedDataSource : DataSource from MeshVS;
  myEmptyMap              : PackedMapOfInteger from TColStd;
  myVectors               : DataMapOfIntegerVector from MeshVS;
  myMagnify               : Real;

end DataSource;
