-- File:	TFace1.cdl
-- Created:	Mon Dec 17 11:18:44 1990
-- Author:	Remi Lequette
--		<rle@topsn3>
---Copyright:	 Matra Datavision 1990, 1992



class TFace1 from PTopoDS inherits TShape1 from PTopoDS

	---Purpose: A topological  Face1.

uses
    ShapeEnum from TopAbs

is
    Create returns mutable TFace1 from PTopoDS;
	---Purpose: the new TFace1 covers the whole 2D space.
    ---Level: Internal 
    	
    ShapeType(me) returns ShapeEnum from TopAbs;
    ---Level: Internal 

end TFace1;
