-- Created on: 1992-04-07
-- Created by: Christian CAILLET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



deferred class TransfEntity  from IGESData  inherits IGESEntity

    ---Purpose : defines required type for Transf in directory part
    --           an effective Transf entity must inherits it

uses GTrsf

is

    Value (me) returns GTrsf  is deferred;
    ---Purpose : gives value of the transformation, as a GTrsf
    --           To be defined by an effective class of Transformation Entity
    --  Warning : Must take in account Composition : if a TransfEntity has in
    --           its Directory Part, a Transf, this means that it is Compound,
    --           Value must return the global result

end TransfEntity;
