-- Created on: 1993-01-09
-- Created by: CKY / Contract Toubro-Larsen ( SIVA )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Sphere from IGESSolid  inherits IGESEntity

        ---Purpose: defines Sphere, Type <158> Form Number <0>
        --          in package IGESSolid
        --          This defines a sphere with a center and radius

uses

        Pnt             from gp,
        XYZ             from gp

is

        Create returns mutable Sphere;

        -- Specific Methods pertaining to the class

        Init (me      : mutable;
              aRadius : Real;
              aCenter : XYZ);
        ---Purpose : This method is used to set the fields of the class Sphere
        --       - aRadius : the radius of the sphere
        --       - aCenter : the center point coordinates (default (0,0,0))

        Radius (me) returns Real;
        ---Purpose : returns the radius of the sphere

        Center (me) returns Pnt;
        ---Purpose : returns the center of the sphere

        TransformedCenter (me) returns Pnt;
        ---Purpose : returns the center of the sphere after applying 
        -- TransformationMatrix

fields

--
-- Class    : IGESSolid_Sphere
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class Sphere.
--
-- Reminder : A Sphere instance is defined by :
--            its center (X1,Y1,Z1) and a radius (Radius) > 0
--

        theRadius : Real;
            -- the radius of the sphere

        theCenter : XYZ;
            -- the center point coordinates

end Sphere;
