-- Created on: 1995-12-04
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.





package RWStepRepr 

uses

	StepData, Interface, TCollection, TColStd, StepRepr

is


--class ReadWriteModule;

--class GeneralModule;

class RWDefinitionalRepresentation;
class RWDescriptiveRepresentationItem;
class RWFunctionallyDefinedTransformation;
class RWGlobalUncertaintyAssignedContext;
class RWGlobalUnitAssignedContext;
class RWItemDefinedTransformation;
--moved to StepBasic: class RWGroup;
--moved to StepBasic: class RWGroupRelationship;
class RWMappedItem;
class RWParametricRepresentationContext;
class RWProductDefinitionShape;
class RWPropertyDefinition;
class RWPropertyDefinitionRepresentation;
--moved to StepAP214: class RWRepItemGroup;
class RWRepresentation;
class RWRepresentationContext;
class RWRepresentationItem;
class RWRepresentationMap;
class RWRepresentationRelationship;

class RWShapeAspect;
class RWShapeAspectRelationship;
class RWShapeAspectTransition;
-- class RWShapeDefinitionRepresentation;  moved to StepShape

    	-- Added from AP214 CC1 to CC2

class RWMakeFromUsageOption;
class RWAssemblyComponentUsage;
class RWQuantifiedAssemblyComponentUsage;
class RWSpecifiedHigherUsageOccurrence;

class RWAssemblyComponentUsageSubstitute;

class RWRepresentationRelationshipWithTransformation;
class RWShapeRepresentationRelationshipWithTransformation;

class RWMaterialDesignation;

-- ABV added for CAX TRJ 2 validation properties
class RWMeasureRepresentationItem;

    -- Added for AP203
    class RWConfigurationDesign;
    class RWConfigurationEffectivity;
    class RWConfigurationItem;
    class RWProductConcept;

    -- Added for Dimensional Tolerancing (CKY 25 APR 2001 for TR7J)
    class RWCompoundRepresentationItem;

	---Package Method ---

--- added for AP209
    class RWDataEnvironment;
    class RWMaterialPropertyRepresentation;
    class RWPropertyDefinitionRelationship;
    class RWMaterialProperty;
    class RWStructuralResponseProperty;
    class RWStructuralResponsePropertyDefinitionRepresentation;

--- added for TR12J (GD&T) 
    class RWCompositeShapeAspect;
    class RWDerivedShapeAspect;
    class RWExtension;
    class RWShapeAspectDerivingRelationship;
    class RWReprItemAndLengthMeasureWithUnit;
    
--	Init;
	---Purpose: enforced the initialisation of the  libraries

end RWStepRepr;
