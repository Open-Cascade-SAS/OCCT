-- Created on: 1993-07-06
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




package BRepPrimAPI 

	---Purpose: The  BRepBuilderAPI  package   provides  an   Application
	--          Programming Interface  for the BRep  topology data
	--          structure.
	--          
	--          The API is a set of classes aiming to provide :
	--          
	--          * High level and simple calls  for the most common
	--          operations. 
	--          
	--          *    Keeping   an   access  on    the    low-level
	--          implementation of high-level calls.
	--          
	--          * Examples  of programming of high-level operations
	--          from low-level operations.
	--          
	--          * A complete coverage of modelling :
	--          
	--             - Creating vertices ,edges, faces, solids.
	--             
	--             - Sweeping operations.
	--             
	--             - Boolean operations.
	--             
	--             - Global properties computation.
	--
	-- 	    
	-- 	    The API provides  classes to  build  objects:
	-- 	    
	-- 	    * The  constructors  of the classes  provides  the
	-- 	    different constructions methods.
	-- 	    
	-- 	    * The  class keeps as fields the   different tools
	-- 	    used to build the object.
	-- 	    
	-- 	    *   The class  provides  a  casting  method to get
	-- 	    automatically the  result  with  a   function-like
	-- 	    call. 
	-- 	    
	-- 	    For example to make a  vertex <V> from a point <P>
	-- 	    one can writes :
	-- 	    
	-- 	    V = BRepBuilderAPI_MakeVertex(P);
	-- 	    
	-- 	    or
	-- 	    
	-- 	    BRepBuilderAPI_MakeVertex MV(P);
	-- 	    V = MV.Vertex();
	-- 	    
	-- 	    
	-- 	    For tolerances  a default precision is  used which
	-- 	    can    be   changed    by    the   packahe  method
	-- 	    BRepBuilderAPI::Precision. 
	-- 	    
	-- 	    For error handling the BRepBuilderAPI commands raise only
	-- 	    the NotDone error. When Done is false on a command
	-- 	    the error description can be asked to the command.
	-- 	    
	-- 	    In  theory  the  comands can be    called with any
	-- 	    arguments, argument  checking  is performed by the
	-- 	    command.
	
	

uses
    StdFail,
    gp,
    TColgp,
    Geom2d,
    Geom,
    GeomAbs,
    TopAbs,
    TopoDS,
    TopTools,
    TopLoc,
    BRep,
    BRepLib,
    BRepTools,
    BRepPrim,
    BRepBuilderAPI, 
    BRepSweep

is
    
    --
    --  Primitives
    --  
    
    class MakeHalfSpace;           ---  inherits MakeShape from BRepBuilderAPI

    class MakeBox;                 ---  inherits MakeShape from BRepBuilderAPI
    
    class MakeWedge;               ---  inherits MakeShape from BRepBuilderAPI
    
    deferred class MakeOneAxis;    ---  inherits MakeShape from BRepBuilderAPI
	---Purpose: Root class for rotational primitives.
    
    class MakeCylinder;            ---  inherits MakeShape from BRepBuilderAPI
    
    class MakeCone;                ---  inherits MakeShape from BRepBuilderAPI
    
    class MakeSphere;              ---  inherits MakeOneAxis from BRepPrimAPI 
    
    class MakeTorus;               ---  inherits MakeOneAxis from BRepPrimAPI
    
    class MakeRevolution;          ---  inherits MakeOneAxis from BRepPrimAPI

    --
    -- Sweeping
    -- 

    deferred class MakeSweep;      ---  inherits MakeShape from BRepBuilderAPI

    class MakePrism;               ---  inherits MakeSweep from BRepPrimAPI
    
    class MakeRevol;               ---  inherits MakeSweep from BRepPrimAPI
    
 


end BRepPrimAPI;
