-- File:	MeshDS_Mesh2d.cdl
-- Created:	Wed Mar 17 11:20:52 1993
-- Author:	Didier PIFFAULT
--		<dpf@phylox>
---Copyright:	 Matra Datavision 1993


generic class Mesh2d from MeshDS
    	    	(Node as any;       -- Signature of Node from MeshDS
    	    	 Link as any;       -- Signature of Link from MeshDS
    	    	 Element as any)    -- Signature of Element2d from MeshDS
     inherits TShared from MMgt

	---Purpose: Describes  the data structure  necessary  for  the
	--          mesh  algorithms  in  two  dimensions  plane or on
	--          surface by meshing in UV space.


uses        Integer from Standard,
    	    ListOfInteger from MeshDS,
      	    MapOfInteger from MeshDS,
	    PairOfIndex from MeshDS,
	    Box from Bnd,
	    BoundSortBox from Bnd,
	    BaseAllocator from MeshDS

    	    class NodeHasher instantiates MapHasher(Node);
    	    class LinkHasher instantiates MapHasher(Link);
    	    class ElemHasher instantiates MapHasher(Element);

	    class IDMapOfNode  instantiates IndexedDataMap from TCollection
    	    	    	    	       (Node,
    	    	    	    	    	ListOfInteger from MeshDS,
    	    	    	    	    	NodeHasher);


	    class IDMapOfLink  instantiates IndexedDataMap from TCollection
    	    	    	    	       (Link,
    	    	    	    	    	PairOfIndex from MeshDS,
    	    	    	    	    	LinkHasher);


	    class IMapOfElement instantiates IndexedMap from TCollection
    	    	    	    	       (Element,
    	    	    	    	    	ElemHasher);

            
    	    class Selector from MeshDS 

    	    	---Purpose: Describes a selector and  an Iterator on a
    	    	--          selector of components of a Mesh.

    	    uses    Integer from Standard,
	            Box from Bnd,
		    MapOfInteger from MeshDS

    	    is	    Create returns Selector from MeshDS;

	    	    Create      (theMesh     : Mesh2d from MeshDS)
    	    	    	returns Selector from MeshDS;

	    	    Initialize  (me          : in out;
    	    	    	         theMesh     : Mesh2d from MeshDS) 
    	    	    	is static;


		    NeighboursOf(me          : in out;
		    	    	 theNode     : in Node) 
    	    	    	is static;

		    NeighboursOfNode(me          : in out;
		    	    	     indexNode   : in Integer from Standard) 
    	    	    	is static;


		    NeighboursOf(me          : in out;
		    	    	 theLink     : in Link) 
    	    	    	is static;

		    NeighboursOfLink(me          : in out;
		    	    	     indexLink   : in Integer from Standard) 
    	    	    	is static;


		    NeighboursOf(me          : in out;
		       	       	 theElem     : in Element) 
    	    	    	is static;

		    NeighboursOfElement(me        : in out;
		    	    	        indexElem : in Integer from Standard) 
			---Purpose: All Neighbours  Of the Element. By
			--          edge or by vertices.
    	    	    	is static;


		    NeighboursByEdgeOf (me        : in out;
		    	    	    	theElem   : in Element) 
			---Purpose: Neighbours by edge Of the Element.
    	    	    	is static;


		    NeighboursOf(me          : in out;
		       	       	 theSelector : in Selector from MeshDS) 
			---Purpose: Adds a level of Neighbours by edge
			--          to the selector <theSelector>.
    	    	    	is static;


		    AddNeighbours(me       : in out)
			---Purpose: Adds a level of Neighbours by edge
			--          to the selector <me>.
    	    	    	is static;


		    Nodes       (me) 
			---C++: return const &
    	    	    	returns  MapOfInteger from MeshDS is static;

		    Links       (me) 
			---C++: return const &
    	    	    	returns  MapOfInteger from MeshDS is static;

		    Elements    (me) 
			---C++: return const &
    	    	    	returns  MapOfInteger from MeshDS is static;

		    FrontierLinks(me) 
			---Purpose: Gives the  list  of links  incices
			--          frontier  of  the  selector  <me>.
			---C++: return const &
    	    	    	returns  MapOfInteger from MeshDS is static;


    	    fields  myMesh      : Mesh2d from MeshDS;
    	    	    myNodes     : MapOfInteger from MeshDS;
    	    	    myLinks     : MapOfInteger from MeshDS;
    	    	    myElements  : MapOfInteger from MeshDS;
	    	    myFrontier  : MapOfInteger from MeshDS;

    	    end Selector;



is          Create     (theAllocator: BaseAllocator from MeshDS;
    	    	    	NodeNumber : Integer from Standard = 100)
	    ---Purpose: <NodeNumber>   is just  an   evaluation of the
	    --          presumed  number of nodes  in this mesh.   The
	    --          Mesh   data  structure will   be automatically
	    --          redimensioned if necessary.
       	    	returns mutable Mesh2d from MeshDS;

    	    AddNode    (me      : mutable ;
    	    	    	theNode : Node) 
    	    	returns Integer from Standard
	    ---Purpose: Adds a node to the  mesh  if  the node is  not
	    --          already in the Mesh.  Returns the index of the
	    --          node in the structure.
		is static;

    	    GetNode    (me      : mutable; 
    	    	    	Index   : Integer from Standard)
    	    	returns any Node 
	    ---Purpose: Get the value of node <Index>.
	    ---C++:  return const &
	    ---C++:  alias operator ()
		is static;

    	    GetNodeList    (me      : mutable; 
    	    	    	    Index   : Integer from Standard)
    	    	returns ListOfInteger from MeshDS
	    ---Purpose: Get the list of node <Index>.
	    ---C++:  return const &
		is static;

    	    ForceRemoveNode (me    : mutable;
	    	    	     Index : Integer from Standard) 
	    ---Purpose: Removes the node of index <index> from the mesh.
	    is static;

    	    ForceRemoveLink (me    : mutable;
  	    	    	     Index : Integer from Standard) 
	    ---Purpose: Removes the link of index <index> from the mesh.
	    is static;

    	    ReplaceNodes (me       : mutable;
  	    	    	  NewNodes : IDMapOfNode from MeshDS) 
	    ---Purpose: Removes the all nodes and sets new map of 
            -- nodes from the mesh.
	    -- For internal use only.
	    is static;

    	    RemoveNode (me      : mutable;
	    	    	Index   : Integer from Standard) 
	    ---Purpose: Removes the node of index <index> from the mesh.
	    is static;

    	    MoveNode   (me      : mutable ;
	    	    	Index   : Integer from Standard;
    	    	    	newNode : Node) 
	    ---Purpose: Changes the UV  value of node of index <Index>  by
	    --          <newNode>. Returns false if <newnode> is already in
	    --          the structure.
	    returns Boolean from Standard is static;

    	    NbNodes        (me)
    	    	    	    returns Integer from Standard
    	    ---Purpose: Gives the number of nodes in this mesh.
	    is static;


    	    AddLink    (me      : mutable;
    	    	    	theLink : Link) 
    	    	returns Integer from Standard
	    ---Purpose: Adds a Link  to the  mesh if  the Link is  not
	    --          already in the structure. Returns the index of
	    --          the link in the structure.
	    is static;

    	    GetLink    (me    : mutable; 
    	    	    	Index : Integer from Standard)
    	    	returns any Link 
	    ---Purpose: Get the value of Link <Index>.
	    ---C++: return const &
		is static;

    	    RemoveLink (me      : mutable;
	    	    	Index   : Integer from Standard) 
	    ---Purpose: Removes the Link of  index  <Index> from the
	    --          mesh.
	    is static;

    	    SubstituteLink (me      : mutable ;
	    	    	    Index   : Integer from Standard;
    	    	    	    newLink : Link) 
	    ---Purpose: Substitutes  the  Link  of  index  <Index>  by
	    --          <newLink> clear the connectivity.
	    returns Boolean from Standard is static;

    	    NbLinks        (me)
    	    	    	    returns Integer from Standard
    	    ---Purpose: Gives the number of elements in this mesh.
	    is static;


    	    AddElement     (me         : mutable;
    	    	    	    theElement : Element) 
    	    	returns Integer from Standard
	    ---Purpose: Adds an element  to  the mesh  if it    is not
	    --          already in the  Mesh. Returns the index of the
	    --          element in the structure.
	    is static;

    	    GetElement     (me    : mutable; 
    	    	    	    Index : Integer from Standard)
    	    	returns any Element
	    ---Purpose: Get the value of Element <Index>.
	    ---C++: return const &
	    is static;

    	    RemoveElement  (me      : mutable;
	    	    	    Index   : Integer from Standard) 
	    ---Purpose: Removes the element of index <Index> in the mesh.
	    is static;

    	    SubstituteElement  (me         : mutable ;
	    	    	    	Index      : Integer from Standard;
    	    	    	    	newElement : Element) 
	    ---Purpose: Substitutes  the  element   of  index  <Index>  by
	    --          <newElement>. The links connectivity is updated.
	    returns Boolean from Standard is static;

    	    NbElements     (me)
    	    	returns Integer from Standard
    	    ---Purpose: Gives the number of elements in this mesh.
	    is static;


    	    ClearDomain        (me         : mutable) 
	    ---Purpose:  Removes all elements
	    is static;


    	    IndexOf        (me;
	    	    	    aNode : Node)
    	    ---Purpose: Finds the index of the node.  Returns 0 if the
    	    --          node is not in the mesh.
	    	returns Integer from Standard;

    	    IndexOf        (me;
	    	    	    aLink : Link)
    	    ---Purpose: Finds the index of the Link.  Returns 0 if the
    	    --          Link is not in the mesh.
	    	returns Integer from Standard;

    	    IndexOf        (me;
	    	    	    anElement : Element)
    	    ---Purpose: Finds the index  of the Element.  Returns 0 if
    	    --          the Element is not in the mesh.
	    	returns Integer from Standard;


    	    LinkNeighboursOf (me;
    	    	    	      theNode         : in Integer from Standard)
	    	returns ListOfInteger from MeshDS
	    ---C++: return const &
    	    ---Purpose: Gives the list of  Link's indices handling the
    	    --          node <theNode>.
	    is static;

    
    	    ElemConnectedTo (me;
    	    	    	     theLink     : in Integer from Standard)
	    	returns PairOfIndex from MeshDS
	    ---C++: return const &
    	    ---Purpose: Gives the element's indices conected
    	    --          to <theLink>.
	    is static;
    
    	    ElemOfDomain     (me)
	    	returns MapOfInteger from MeshDS
	    ---C++: return const &
    	    ---Purpose: Gives  the  list  of element's indices
	    is static;


    	    LinkOfDomain     (me)
	    	returns MapOfInteger from MeshDS
	    ---C++: return const &
    	    ---Purpose: Gives  the  list  of link's indices
	    is static;


    	    ClearDeleted     (me : mutable)
    	    ---Purpose: This method  substitute the deleted  items  by
    	    --          the last in  Indexed Data  Maps  to  have only
    	    --          non-deleted  elements, links  or  nodes in the
    	    --          structure.
	    is static;


-- Internal methods :

    	    ClearElement   (me      : mutable;
	    	    	    Index   : Integer from Standard;
	    	    	    theElem : Element) 
	    ---Purpose: Deletes  the element of  index <Index> in
	    --          the mesh. Used by RemoveElement.
	    is static private;

    	    Statistics     (me;
	    	    	    flot  : in out OStream from Standard) 
	    ---Purpose: Give informations on map.
	    is static;
	    
	    Allocator (me) returns BaseAllocator from MeshDS;
	    	---C++: return const&

    
fields      myNodes        : IDMapOfNode   from MeshDS;
    	    myDelNodes     : ListOfInteger from MeshDS;
    	    myLinks        : IDMapOfLink   from MeshDS;
    	    myDelLinks     : ListOfInteger from MeshDS;
    	    myElements     : IMapOfElement from MeshDS;
    	    --myDelElements  : ListOfInteger from MeshDS;
	    myElemOfDomain : MapOfInteger  from MeshDS;
	    myLinkOfDomain : MapOfInteger  from MeshDS;
	    myAllocator    : BaseAllocator from MeshDS;
end Mesh2d;
