-- Created on: 1997-02-28
-- Created by: Christophe LEYNADIER
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

private class TypedCallBack from Storage 

inherits TShared from MMgt

uses CallBack from Storage,
     AsciiString from TCollection
     
is
    Create returns TypedCallBack from Storage;

    Create(aTypeName : AsciiString from TCollection; aCallBack : CallBack from Storage)
    	returns TypedCallBack from Storage;

    SetType(me : mutable; aType : AsciiString from TCollection);
    Type(me) returns AsciiString from TCollection;
    
    SetCallBack(me : mutable; aCallBack : CallBack from Storage);
    CallBack(me) returns CallBack from Storage;

    SetIndex(me : mutable; anIndex : Integer from Standard);
    Index(me) returns Integer from Standard;
    
    fields
    
    	myType     : AsciiString from TCollection;
	myCallBack : CallBack from Storage;
    	myIndex    : Integer from Standard;
	
end;
