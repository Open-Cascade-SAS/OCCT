-- Created on: 1997-09-11
-- Created by: Philippe MANGIN
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



deferred class SmoothCriterion from AppParCurves
inherits  TShared  from MMgt

	---Purpose: defined criterion to smooth  points in  curve
                             

uses
   Vector  from  math, 
   Matrix  from  math, 
   Curve   from  FEmTool, 
   HAssemblyTable    from  FEmTool,  
   HArray2OfInteger  from TColStd, 
   HArray1OfReal    from TColStd,
   Array1OfReal    from TColStd 
    
raises 
  NotImplemented,   
  DomainError 
   
 

is 
    SetParameters(me  :  mutable;  Parameters  : HArray1OfReal) 
    is  deferred; 

    SetCurve(me  :  mutable;  C  :Curve from FEmTool) 
    is  deferred; 
     
    GetCurve(me;  C  :  out  Curve  from FEmTool) 
    is  deferred; 
     
    SetEstimation(me  :  mutable;  E1,  E2,  E3  :  Real)   
    is  deferred; 
     
    EstLength(me  :  mutable)   
    ---C++: return &
    returns  Real  is  deferred;     
     
    GetEstimation(me;  E1,  E2,  E3  : out Real)   
    is  deferred; 
     
    AssemblyTable(me)  
    returns HAssemblyTable  from  FEmTool   
    is  deferred; 
     
    DependenceTable(me)  
    returns  HArray2OfInteger  from TColStd   
    is  deferred;  
    
    QualityValues  (me : mutable; J1min,  J2min,  J3min  :  Real; 
    	    	    	    	  J1,  J2,  J3  :  out  Real)
    returns  Integer  is  deferred;
     
    ErrorValues(me  :  mutable;   
                MaxError,  QuadraticError,  AverageError  :  out  Real) 
    is  deferred;
     
    Hessian(me  :  mutable ;  
            Element    :  Integer; 
	    Dimension1  :  Integer; 
	    Dimension2  :  Integer;
            H  :  out  Matrix  from  math)  
     raises  DomainError -- If DependenceTable(Dimension1,Dimension2) is False 
     is  deferred;  
   
    
    Gradient(me  :  mutable;  
             Element  :  Integer; 
	     Dimension  :  Integer;
             G  :  out  Vector  from  math) 
    is  deferred; 
    
    InputVector(me  :  mutable;  X : Vector from math;   
                                 AssTable  :  HAssemblyTable  from  FEmTool)  
    ---Purpose: Convert the assembly Vector in an Curve;
    --          
    raises  DomainError  is  deferred; 
     
    SetWeight(me:  mutable;  
              QuadraticWeight,  QualityWeight  :  Real; 
	      percentJ1,  percentJ2,  percentJ3  :  Real) 
    is  deferred;  
     
    GetWeight(me;  QuadraticWeight,  QualityWeight  :  out  Real)  
    is  deferred;  
     
    SetWeight(me:  mutable;  
              Weight  :  Array1OfReal)
    is  deferred;
          
end SmoothCriterion;












