-- Created on: 2000-11-21
-- Created by: Peter KURNEV
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class ShapeShapeInterference from BOPTools 

	---Purpose: 
	--  Root class for storing  an  Interference        
	--  between a couple BRep shapes  
is
    Create 
    	returns ShapeShapeInterference from BOPTools;  
    	---Purpose:  
    	--- Empty constructor 
    	---
    Create (anIndex1:  Integer from Standard;  
    	    anIndex2:  Integer from Standard)
    	returns ShapeShapeInterference from BOPTools;  
    	---Purpose:   
    	--- Constructor 
    	---
    SetIndex1(me:out; anIndex1:Integer from Standard);  
    	---Purpose:  
    	--- Modifier  
    	--- Sets DS-index for the first shape from the  couple 
    	---
    SetIndex2(me:out; anIndex2:Integer from Standard);   
    	---Purpose:  
    	--- Modifier 
    	--- Sets DS-index for the second shape from the  couple  
    	---
    SetNewShape(me:out; anIndex:Integer from Standard);   
    	---Purpose:  
    	--- Modifier   
    	--- Sets DS-index for the new shape 
    	---
    Index1(me) 
    	returns Integer from Standard;
    	---Purpose:  
    	--- Selector  
    	---
    Index2(me) 
    	returns Integer from Standard;
    	---Purpose:  
    	--- Selector  
    	---
    Indices(me; 
    	    anIndex1:out Integer from Standard;	      
    	    anIndex2:out Integer from Standard); 
    	---Purpose:  
    	--- Selector  
    	---
    OppositeIndex(me; 
    	     anIndex:Integer from Standard) 
    	returns Integer from Standard; 		     
    	---Purpose:  
    	--- Selector  
    	--- Gets the value of index 
    	--- if  anIndex==myIndex1 it returns myIndex2; 
    	--- if  anIndex==myIndex2 it returns myIndex1; 
    	--- otherwise it returns 0; 
    	---
    NewShape(me) 
    	returns Integer from Standard; 
     	---Purpose:  
    	--- Selector  
    	---

fields
    myIndex1  : Integer from Standard; 
    myIndex2  : Integer from Standard; 
    myNewShape: Integer from Standard; 
    
end ShapeShapeInterference;
