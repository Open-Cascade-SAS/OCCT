-- Created on: 1992-05-06
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package IntPatch 

	---Purpose: Intersection between two patches.
	--          The class PatchIntersection implements the algorithmes
	--          of intersection.
	--          The classes IntPoint, PointOnDomain, Line, ILin, a.s.o...
	--          describe the results of the algorithmes.

        ---Level: Internal
        --
        -- All the methods of the classes of this package are Internal.
	--

uses Standard, MMgt, StdFail, GeomAbs, TopAbs, TCollection, TColStd, math, 
     gp, TColgp, IntAna,IntSurf, IntImp, IntStart, IntWalk, Bnd, Intf,  
     Adaptor2d,Adaptor3d, Geom2d, Geom, Precision

is

    class ALineToWLine;

    class Point;

    deferred class Line;
    
    	class GLine;      -- inherits Line from IntPatch

    	class ALine;      -- inherits Line from IntPatch
    
    	class WLine;      -- inherits Line from IntPatch
    
    	class RLine;      -- inherits Line from IntPatch

    class ArcFunction;

-- implicite/implicite

    class ImpImpIntersection;


-- commun implicite/parametree et parametree/parametree

    deferred class Polygo;
      
    	class PolyLine;    -- inherits Polygo from IntPatch

        class PolyArc;     -- inherits Polygo from IntPatch

    class RstInt;


-- implicite/parametre

    class ImpPrmIntersection;


-- parametre/parametre

    class Polyhedron;

    class PolyhedronTool;
    
    class PrmPrmIntersection_T3Bits;

    class PrmPrmIntersection;


-- algorithme general

    enumeration IType is
    -- type of the line of intersection

    	Lin,       -- pour conflit avec deferred class Line
    	Circle,
    	Ellipse,
    	Parabola,
    	Hyperbola,
    	Analytic,
        Walking,
    	Restriction
    end IType;

    class HInterTool;

    class HCurve2dTool;

    class LineConstructor;

    class Intersection;


    class SequenceOfPoint instantiates Sequence from TCollection (Point from IntPatch);

    class SequenceOfLine instantiates Sequence from TCollection (Line from IntPatch);

    class TheSurfFunction instantiates ZerImpFunc from IntImp
        (HSurface     from Adaptor3d,
         HSurfaceTool from Adaptor3d,
         Quadric      from IntSurf,
         QuadricTool  from IntSurf);

    class TheIWalking instantiates IWalking from IntWalk
        (PathPoint               from IntSurf, 
         PathPointTool           from IntSurf,
         SequenceOfPathPoint     from IntSurf,
         InteriorPoint           from IntSurf,
         InteriorPointTool       from IntSurf,
         SequenceOfInteriorPoint from IntSurf,
         HSurface                from Adaptor3d,
         HSurfaceTool            from Adaptor3d,
         TheSurfFunction         from IntPatch);

    class TheSearchInside instantiates SearchInside from IntStart
        (HSurface        from Adaptor3d,
         HSurfaceTool    from Adaptor3d,
         TopolTool       from Adaptor3d,
         HInterTool      from IntPatch,
         TheSurfFunction from IntPatch);

    class TheSOnBounds instantiates SearchOnBoundaries from IntStart(
         HVertex from Adaptor3d,
         HCurve2d from Adaptor2d,
         HCurve2dTool from IntPatch,
         HInterTool from IntPatch,
         TopolTool from Adaptor3d,
         ArcFunction from IntPatch);

    class TheInterfPolyhedron instantiates InterferencePolyhedron from Intf(
              Polyhedron from IntPatch,
              PolyhedronTool from IntPatch,
              Polyhedron from IntPatch,
              PolyhedronTool from IntPatch);

    class ThePWalkingInter instantiates PWalking from IntWalk(
              HSurface     from Adaptor3d,
              HSurfaceTool from Adaptor3d);

    alias SearchPnt is InterferencePolygon2d from Intf;

    class CSFunction instantiates ZerCOnSSParFunc from IntImp
    	(HSurface from Adaptor3d,
         HSurfaceTool from Adaptor3d,
         HCurve2d from Adaptor2d,
         HCurve2dTool from IntPatch);

    class CurvIntSurf instantiates IntCS from IntImp
    	(HSurface from Adaptor3d,
         HSurfaceTool from Adaptor3d,
         HCurve2d from Adaptor2d,
         HCurve2dTool from IntPatch,
         CSFunction from IntPatch);

end IntPatch;
