-- File:	PGeom2d_AxisPlacement.cdl
-- Created:	Tue Apr  6 16:31:20 1993
-- Author:	Philippe DAUTRY
--		<fid@mastox>
-- Copyright:	 Matra Datavision 1993


class AxisPlacement from PGeom2d inherits Geometry from PGeom2d

        ---Purpose :   An  axis  placement  defines a  local cartesian
        --         coordinate  system and   can be used to  locate  an
        --         entity in 3D space.
        --  

uses Ax2d from gp

is


    Create returns mutable AxisPlacement from PGeom2d;
	---Purpose: Initializes the field(s) with default value(s).
	---Level: Internal 


    Create(aAxis: Ax2d from gp) returns mutable AxisPlacement from PGeom2d;
	---Purpose: Initializes the field axis with <aAxis>.
	---Level: Internal 


  Axis (me : mutable; aAxis : Ax2d from gp);
        --- Purpose : Set the field axis with <aAxis>.
	---Level: Internal 


  Axis (me)  returns Ax2d from gp;
        --- Purpose : Returns the value of the field axis.
	---Level: Internal 


fields

  axis : Ax2d from gp;

end;
