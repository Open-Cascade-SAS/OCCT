-- File:	FuncExtPS.cdl
-- Created:	Wed Jul 24 14:31:49 1991
-- Author:	Michel CHAUVAT
--		<mca@topsn3>
---Copyright:	 Matra Datavision 1991

-- Modified by skv - Thu Sep 30 15:19:59 2004 OCC593


private class FuncExtPS from Extrema

 inherits FunctionSetWithDerivatives from math
    ---Purpose: Function to find the extrema of the 
    --          distance between a point and a surface.

uses    POnSurf           from Extrema,
	SequenceOfPOnSurf from Extrema,
	SequenceOfReal    from TColStd,
	Pnt               from gp,
	Vector            from math,
	Matrix            from math,
	Surface           from Adaptor3d,
    	SurfacePtr        from Adaptor3d

raises  OutOfRange from Standard

is
    Create returns FuncExtPS;

    Create (P: Pnt; S: Surface from Adaptor3d) returns FuncExtPS;
    	---Purpose:

    Initialize(me: in out; S: Surface from Adaptor3d)
    	---Purpose: sets the field mysurf of the function.
    is static;
    
    SetPoint(me: in out; P: Pnt)
    	---Purpose: sets the field mysurf of the function.
    is static;

    ------------------------------------------------------------
    -- In all next methods, an exception is raised if the fields 
    -- were not initialized.

    NbVariables (me) returns Integer;

    NbEquations (me) returns Integer;

    Value (me: in out; UV: Vector; F: out Vector) returns Boolean;
    	---Purpose: Calculate Fi(U,V).

    Derivatives (me: in out; UV: Vector; DF: out Matrix)
    	returns Boolean;
    	---Purpose: Calculate Fi'(U,V).

    Values (me: in out; UV: Vector; F: out Vector; DF: out Matrix)
    	returns Boolean;
    	---Purpose: Calculate Fi(U,V) and Fi'(U,V).

    GetStateNumber (me: in out) returns Integer
    	---Purpose: Save the found extremum.
    	is redefined;

    NbExt (me) returns Integer;
    	---Purpose: Return the number of found extrema.

    SquareDistance (me; N: Integer) returns Real
    	---Purpose: Return the value of the Nth distance.
    	raises  OutOfRange;
	    	-- if N < 1 or N > NbExt(me).

    Point (me; N: Integer) returns POnSurf
    	---Purpose: Returns the Nth extremum.
    	raises  OutOfRange;
	    	-- if N < 1 or N > NbExt(me).

-- Modified by skv - Thu Sep 30 15:19:59 2004 OCC593 Begin
    HasDegIso(me) returns Boolean from Standard;
-- Modified by skv - Thu Sep 30 15:19:59 2004 OCC593 End

    Bidon(me) returns SurfacePtr from Adaptor3d
    is static private;
 
fields
    myP    : Pnt from gp;
    myS    : SurfacePtr from Adaptor3d;

    myU    : Real;          -- current value of U
    myV    : Real;          -- current value of V
    myPs   : Pnt from gp;   -- current point

    mySqDist: SequenceOfReal    from TColStd;
    myPoint: SequenceOfPOnSurf from Extrema;
    myPinit: Boolean;
    mySinit: Boolean;
    myUIsoIsDeg: Boolean;
    myVIsoIsDeg: Boolean;

end FuncExtPS;
