-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class VectorOrDirection from StepGeom inherits SelectType from StepData

	-- <VectorOrDirection> is an EXPRESS Select Type construct translation.
	-- it gathers : Vector, Direction

uses

	Vector,
	Direction
is

	Create returns VectorOrDirection;
	---Purpose : Returns a VectorOrDirection SelectType

	CaseNum (me; ent : Transient) returns Integer;
	---Purpose: Recognizes a VectorOrDirection Kind Entity that is :
	--        1 -> Vector
	--        2 -> Direction
	--        0 else

	Vector (me) returns any Vector;
	---Purpose : returns Value as a Vector (Null if another type)

	Direction (me) returns any Direction;
	---Purpose : returns Value as a Direction (Null if another type)


end VectorOrDirection;

