-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


package XmlMDataStd 

        ---Purpose: Storage and Retrieval drivers for modelling attributes.
        --          Transient attributes are defined in package TDataStd.

uses XmlMDF,
     XmlObjMgt,
     TDF,
     CDM

is
        ---Purpose: Storage/Retrieval drivers for TDataStd attributes
        --          =======================================

        class NameDriver;

        class IntegerDriver;
        
        class RealDriver;
        
        class IntegerArrayDriver;
        
        class RealArrayDriver;
        
        class ExtStringArrayDriver;
        
        class UAttributeDriver;
        
        class DirectoryDriver;
        
        class CommentDriver;
        
        class VariableDriver;
        
        class ExpressionDriver;
        
        class RelationDriver;
        
        class NoteBookDriver;
        
        class TreeNodeDriver;  
	
	-- Extension	 
        class TickDriver;

        -- Lists:
       class IntegerListDriver; 
       class RealListDriver;
       class ExtStringListDriver;
       class BooleanListDriver;
       class ReferenceListDriver;
    
       -- Arrays:
       class BooleanArrayDriver;
       class ReferenceArrayDriver;
       class ByteArrayDriver;


       class NamedDataDriver;  
       class AsciiStringDriver;
       class IntPackedMapDriver; 

    AddDrivers (aDriverTable : ADriverTable  from XmlMDF;
                anMsgDrv     : MessageDriver from CDM);
        ---Purpose: Adds the attribute drivers to <aDriverTable>.  
	
    SetDocumentVersion (DocVersion  : Integer from Standard); 
    
    DocumentVersion returns Integer from Standard; 	

end XmlMDataStd;
