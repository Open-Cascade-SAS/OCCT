-- Created on: 1996-09-16
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class BuildShape from LocOpe

	---Purpose: 

uses Shape       from TopoDS,
     ListOfShape from TopTools


is

    Create
    	returns BuildShape from LocOpe;
	---C++: inline


    Create(L: ListOfShape from TopTools)
	---Purpose: Builds shape(s) from  the list <L>.  Uses only the
	--          faces of <L>.
	---C++: inline
    
    	returns BuildShape from LocOpe;


    Perform(me: in out; L: ListOfShape from TopTools)
	---Purpose: Builds shape(s) from  the list <L>.  Uses only the
	--          faces of <L>.
    
    	is static;

    Shape(me)
    
	---C++: inline
	---C++: return const&
    	returns Shape from TopoDS
	is static;


fields

    myRes : Shape from TopoDS;

end BuildShape;
