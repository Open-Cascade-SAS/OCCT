-- Created on: 1992-10-22
-- Created by: Gilles DEBARBOUILLE
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Material from Materials 

	---Purpose: This  class describes  the facilities available to
	--          create and manipulate materials.

inherits

    FuzzyInstance from Materials
    
uses

    HAsciiString from TCollection,
    AsciiString from TCollection

--raises

is

    Create(amaterial : CString from Standard)
    
    ---Level: Internal 
    
    ---Purpose: Creates the material <amaterial>.
    
    returns mutable Material from Materials;
    
    Name(me) returns AsciiString from TCollection
    
    ---Level: Public 
    
    ---Purpose: Returns the name of the material.
    
    is static;
    
    Dump(me ; astream : in out OStream)
    
    ---Level: Internal 
    
    ---Purpose: Useful for debugging.
    
    is redefined;
    
fields

    thematerial      : HAsciiString from TCollection;

end Material;
