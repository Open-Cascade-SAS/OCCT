-- Created on: 1991-09-02
-- Created by: NW,JPB,CAL
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class AspectMarker from Aspect

inherits

	TShared

	---Purpose: This class allows the definition of a group
	--	    of attributes for the primitive MARKER.
	--	    the attributes are:
	--		* Colour
	--		* Type
	--		* Scale factor
	--	    When any value of the group is modified
	--	    all graphic objects using the group are modified

uses

	Color		from Quantity,

	TypeOfMarker 	from Aspect

raises

	AspectMarkerDefinitionError 	from Aspect

is

	Initialize;
	---Level: Public
	---Purpose: Initialise the constructor for Graphic3d_AspectMarker3d.
	--
	-- defaults values :
	--
	--	Color	= Quantity_NOC_YELLOW;
	--	Type	= Aspect_TOM_X;
	--	Scale	= 1.0;

	Initialize ( AColor	: Color from Quantity;
		     AType	: TypeOfMarker from Aspect;
		     AScale	: Real from Standard )
	---Level: Public
	---Purpose: Initialise the values for the
	--	    constructor of Graphic3d_AspectMarker3d.
	--  Warning: Raises AspectMarkerDefinitionError if the
	--	    scale is a negative value.
	raises AspectMarkerDefinitionError from Aspect;

	---------------------------------------------------
	-- Category: Methods to modify the class definition
	---------------------------------------------------

	SetColor ( me		: mutable;
		   AColor	: Color from Quantity );
	---Level: Public
	---Purpose: Modifies the colour of <me>.
	---Category: Methods to modify the class definition

	SetScale ( me		: mutable;
		   AScale	: Real from Standard )
	---Level: Public
	---Purpose: Modifies the scale factor of <me>.
	--	    Marker type Aspect_TOM_POINT is not affected
	--	    by the marker size scale factor. It is always
	--	    the smallest displayable dot.
	--  Warning: Raises AspectMarkerDefinitionError if the
	--	    scale is a negative value.
	raises AspectMarkerDefinitionError from Aspect;

	SetType ( me	: mutable;
		  AType	: TypeOfMarker from Aspect );
	---Level: Public
	---Purpose: Modifies the type of marker <me>.
	---Category: Methods to modify the class definition

	----------------------------
	-- Category: Inquire methods
	----------------------------

	Values ( me;
		 AColor	: out Color from Quantity;
		 AType	: out TypeOfMarker from Aspect;
		 AScale	: out Real from Standard );
	---Level: Public
	---Purpose: Returns the current values of the group <me>.
	---Category: Inquire methods

--

fields

--
-- Class	:	Aspect_AspectMarker
--
-- Purpose	:	Declaration of variables specific to the context of
--			drawing markers
--
-- Reminder	:	A drawing context for markers is defined by :
--			- the colour
--			- the type
--			- the scale
--

	-- the colour
	MyColor	:	Color from Quantity;

	-- the type
	MyType	:	TypeOfMarker from Aspect;

	-- the scale
	MyScale	:	Real from Standard;

end AspectMarker;
