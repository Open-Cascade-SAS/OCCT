-- File:	StepShape_LimitsAndFits.cdl
-- Created:	Tue Apr 24 13:48:52 2001
-- Author:	Atelier IED
--		<ied@photox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 2001

class LimitsAndFits  from StepShape    inherits TShared

    ---Purpose : Added for Dimensional Tolerances

uses
    HAsciiString from TCollection

is

    Create returns mutable LimitsAndFits;

    Init (me : mutable; form_variance, zone_variance, grade, source :
    	    	        HAsciiString from TCollection);

    FormVariance (me) returns HAsciiString from TCollection;
    SetFormVariance (me : mutable; form_variance : HAsciiString from TCollection);

    ZoneVariance (me) returns HAsciiString from TCollection;
    SetZoneVariance (me : mutable; zone_variance : HAsciiString from TCollection);

    Grade (me) returns HAsciiString from TCollection;
    SetGrade (me : mutable; grade : HAsciiString from TCollection);

    Source (me) returns HAsciiString from TCollection;
    SetSource (me : mutable; source : HAsciiString from TCollection);

fields

    theFormVariance : HAsciiString from TCollection;
    theZoneVariance : HAsciiString from TCollection;
    theGrade  : HAsciiString from TCollection;
    theSource : HAsciiString from TCollection;

end LimitsAndFits;
