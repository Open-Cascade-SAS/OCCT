-- Created on: 1992-09-18
-- Created by: Odile Olivier
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Drawer from AIS inherits Drawer from Prs3d

	---Purpose: 
    	-- A framework to manage display attributes of interactive objects.
    	-- An interactive object can have a certain number of
    	-- display attributes specific to it. These include
    	-- visualization mode, color, material
    	-- and so on. To deal with this information, the
    	-- interactive context has a Drawer attribute manager
    	-- which is valid by default for the objects it
    	-- controls.   When an interactive object is visualized, the
    	-- required graphic display attributes are first taken from
    	-- its own Drawer if it has the ones required, or from the
    	-- context drawer for those it does not have them.
    	-- The set of display attributes of an interactive object is
    	-- stocked in an AIS_Drawer, which is, in fact, a
    	-- Prs3d_Drawer with the possibility of a link to another
    	-- display attribute manager. This drawer then manages
    	-- the stocked graphic display attributes by specifying
    	-- how the presentation algorithms compute the
    	-- presentation of a specific kind of object. These
    	-- factors involved include color, width and type of line,
    	-- and maximal chordal deviation. The Drawer includes
    	-- instances of the aspect classes providing the default
    	-- values for them.
    	-- Prs3d_Drawer completes   AIS_Drawer by adding
    	-- functions for setting deviation angle and deviation
    	-- coefficient in presentations using hidden line removal.
        
uses
    Drawer from Prs3d,
    DatumAspect from Prs3d,
    LineAspect from Prs3d,
    TextAspect from Prs3d,
    PointAspect from Prs3d,
    ShadingAspect from Prs3d,
    IsoAspect from Prs3d,
    DimensionAspect from Prs3d,
    PlaneAspect from Prs3d,
    ArrowAspect from Prs3d,
    TypeOfDeflection from Aspect,
    NameOfColor from Quantity,
    PlaneAngle from Quantity,
    Length from Quantity,
    DimensionUnits from Prs3d,
    VertexDrawMode from Prs3d,
    AsciiString from TCollection,
    TypeOfHLR from Prs3d,
    Ax2 from gp

is
    Create returns Drawer from AIS;
    	 ---Purpose:
    	 -- Constructs an empty attribute management framework.   
    TypeOfDeflection(me) returns TypeOfDeflection from Aspect
    is redefined static;
    	 --- Purpose:
    	 -- Returns the type of chordal deflection: relative to the
    	 -- size of the object or absolute.  
    
    MaximalChordialDeviation (me) returns Length from Quantity
	 ---Purpose: Returns the maximal chordal deviation. The default
    	 -- value is 0.1. Drawings of curves or patches are
    	 -- made with respect to an absolute maximal chordal deviation.
    is redefined static;
	    

------------------------------------------------------------                                                               
    SetDeviationCoefficient(me: mutable) ;
	 ---Purpose: Sets the hasOwnDeviationCoefficient flag to Standard_False 
	 ---C++: inline

    SetHLRDeviationCoefficient(me: mutable) ;
	 ---Purpose: Sets the deviation coefficient aCoefficient for
 	 -- removal of hidden lines created by different
	 -- viewpoints in different presentations. The Default value is 0.02.
	 ---C++: inline
         
    SetDeviationAngle(me: mutable) ;
	 ---Purpose: Sets the hasOwnDeviationAngle flag to Standard_False 
	 ---C++: inline

    SetHLRAngle(me: mutable) ;
	 ---Purpose: Sets the angle of maximum chordal deviation for
    	 -- removal of hidden lines created by different viewpoints 
    	 -- in different presentations. The default value is 20*PI/180.
	 ---C++: inline
		    
    SetDeviationCoefficient(me: mutable; aCoefficient: Real from Standard )   
	 ---Purpose: Sets the hasOwnDeviationCoefficient flag to Standard_True,
    	 --          sets myOwnDeviationCoefficient and  myPreviousDeviationCoefficient
    is redefined static;
    
    SetHLRDeviationCoefficient(me: mutable; aCoefficient: Real from Standard )   
	 ---Purpose: Sets the hasOwnHLRDeviationCoefficient flag to Standard_True,
	 --          sets myOwnHLRDeviationCoefficient and  myPreviousHLRDeviationCoefficient
    is redefined static;
        
    SetDeviationAngle(me: mutable; anAngle: Real from Standard )  is redefined ;
	 ---Purpose: Sets the hasOwnDeviationAngle flag to Standard_True,
	 --          sets myOwnDeviationAngle and  myPreviousDeviationAngle
    	
    SetHLRAngle(me: mutable; anAngle: Real from Standard )   
	 ---Purpose: Sets the hasOwnHLRDeviationAngle flag to Standard_True,
	 --          sets myOwnHLRDeviationAngle and  myPreviousHLRDeviationAngle
    is redefined static;

    SetTypeOfHLR(me: mutable; theTypeOfHLR: TypeOfHLR from Prs3d)
    is redefined;
    ---Purpose: Sets the type of HLR algorithm
    --          used by drawer's interactive objects
    ---C++: inline
    
    TypeOfHLR(me) returns TypeOfHLR from Prs3d
    is redefined;
    ---Purpose: Returns the type of HLR algorithm currently in use.
    ---C++: inline

    DeviationCoefficient(me) returns Real from Standard
     	 ---Purpose: Drawings of curves or patches are made with respect
    	 -- to a maximal chordal deviation. A Deviation coefficient
    	 -- is used in the shading display mode. The shape is
    	 -- seen decomposed into triangles. These are used to
    	 -- calculate reflection of light from the surface of the
    	 -- object. The triangles are formed from chords of the
    	 -- curves in the shape. The deviation coefficient gives
    	 -- the highest value of the angle with which a chord can
    	 -- deviate from a tangent to a   curve. If this limit is
    	 -- reached, a new triangle is begun.
    	 -- This deviation is absolute and is set through the
    	 -- method: SetMaximalChordialDeviation. The default value is 0.001.
    	 -- In drawing shapes, however, you are allowed to ask
    	 -- for a relative deviation. This deviation will be:
    	 -- SizeOfObject * DeviationCoefficient.
    is redefined static;
    
    HLRDeviationCoefficient(me) returns Real from Standard
        ---Purpose: Returns the real number value of the HLR deviation
    	-- coefficient in this framework, if the flag
    	-- hasOwnHLRDeviationCoefficient is true.
    	-- If hasOwnHLRDeviationCoefficient is false, the
    	-- shape's HLR deviation coefficient is used.
    	-- A Deviation coefficient is used in the shading display
    	-- mode. The shape is seen decomposed into triangles.
    	-- These are used to calculate reflection of light from the
    	-- surface of the object.
    	-- The triangles are formed from chords of the curves in
    	-- the shape. The deviation coefficient give the highest
    	-- value of the angle with which a chord can deviate
    	-- from a tangent to a curve. If this limit is reached, a
    	-- new triangle is begun.
    	-- To find the hidden lines, hidden line display mode
    	-- entails recalculation of the view at each different
    	-- projector perspective.
    	-- Since hidden lines entail calculations of more than
    	-- usual complexity to decompose them into these
    	-- triangles, a deviation coefficient allowing greater
    	-- tolerance is used. This increases efficiency in calculation.
    	-- The Default value is 0.02.
    is redefined static;   
    
    
    DeviationAngle(me) returns Real from Standard
	---Purpose: Returns myOwnDeviationAngle if hasOwnDeviationAngle is True
	--          else gets myDeviationAngle field from Prs3d_Drawer 
    is redefined;
      		
    HLRAngle(me) returns Real from Standard
	---Purpose: Returns the real number value of the deviation angle
    	-- in hidden line removal views. The default value is 20*PI/180.
        is redefined static;              
    
    
    PreviousDeviationCoefficient(me) returns Real from Standard
	---Purpose: Saves the previous value used for the chordal
	-- deviation coefficient. The default value is 0.1.
	---C++: inline
    is static;          
  
    PreviousHLRDeviationCoefficient(me) returns Real from Standard
	---Purpose: returns myPreviousHLRDeviationCoefficient
	---C++: inline
    is static;

    PreviousDeviationAngle(me) returns Real from Standard
	---Purpose: returns myPreviousDeviationAngle
	---C++: inline
    is  static;

    PreviousHLRDeviationAngle(me) returns Real from Standard
	---Purpose: returns myPreviousHLRDeviationAngle
	---C++: inline 
    is  static;
    
    IsOwnDeviationCoefficient(me) returns Boolean from Standard;
    	---Purpose: Returns true if the there is a local setting for deviation
    	-- coefficient in this framework for a specific interactive object.
        ---C++: inline
             
    IsOwnHLRDeviationCoefficient(me) returns Boolean from Standard;
    	---Purpose: Returns true if the there is a setting for HLR deviation
    	-- coefficient in this framework for a specific interactive object.
        ---C++: inline
     							       
    IsOwnDeviationAngle(me) returns Boolean from Standard;
     	---Purpose: Returns true if the there is a local setting for deviation
    	-- angle in this framework for a specific interactive object.
        ---C++: inline

    IsOwnHLRDeviationAngle(me) returns Boolean from Standard;
    	---Purpose: Returns true if the there is a setting for HLR deviation
    	-- angle in this framework for a specific interactive object.
    	---C++: inline

    Discretisation(me) returns Integer from Standard
    is redefined static;
    	---Purpose: Draws algorithms using discretisation, a default
    	-- number of points has been set to 17. You can use the
    	-- method Prs3d_Drawer_SetDiscretisation to change this value. 
    
    MaximalParameterValue(me) returns Real from Standard
    is redefined static;
    	---Purpose:
    	-- Sets the maximum value allowed for the first and last
    	-- parameters of an infinite curve. By default, this value is 500000.
    
    IsoOnPlane(me) returns Boolean from Standard 
	---Purpose: returns True if the drawing of isos on planes is enabled.
    is redefined static;


-- 
-- Attributes for the U Isoparametric lines of patches.
--    
    UIsoAspect (me:mutable) returns IsoAspect from Prs3d
	 ---Purpose: Defines the attributes which are used when drawing an 
	 --          U isoparametric curve of a face. Defines the number
	 --          of U isoparametric curves to be drawn for a single face.
	 --          The LineAspect for U isoparametric lines can be edited
	 --          (methods SetColor, SetTypeOfLine, SetWidth, SetNumber)
	 --          The default values are:
	 --          COLOR       : Quantity_NOC_GRAY75
         --          TYPE OF LINE: Aspect_TOL_SOLID
   	 --          WIDTH       : 0.5
    	 -- These attributes are used by the following algorithms:
	 --          Prs3d_WFDeflectionSurface 
	 --          Prs3d_WFDeflectionRestrictedFace


    is redefined static;    
    
    HasUIsoAspect (me) returns Boolean from Standard 
	 ---Purpose: Returns true if the Drawer has a UIso aspect setting active.
	 ---C++: inline
   is static;

-- Attributes for the V Isoparametric line of patches.


    VIsoAspect (me:mutable) returns IsoAspect from Prs3d
	 ---Purpose: Defines the attributes which are used when drawing an 
	 --          V isoparametric curve of a face. Defines the number
	 --          of V isoparametric curves to be drawn for a single face.
	 --          The LineAspect for V isoparametric lines can be edited
	 --          (methods SetColor, SetTypeOfLine, SetWidth, SetNumber)
	 --          The default values are:
	 --          COLOR       : Quantity_NOC_GRAY82
	 --          TYPE OF LINE: Aspect_TOL_SOLID
	 --          WIDTH       : 0.5
	 --          These attributes are used by the following algorithms:
	 --          Prs3d_WFDeflectionSurface 
	 --          Prs3d_WFDeflectionRestrictedFace
    is redefined static;    

    HasVIsoAspect (me) returns Boolean from Standard 
	 ---Purpose: Returns true if the Drawer has a VIso aspect setting active.
	 ---C++: inline
   is static;    

-- Attributes for the free boundaries

    FreeBoundaryAspect (me:mutable) returns LineAspect from Prs3d
	 ---Purpose: Returns a link with
    	 -- Prs3d_Drawer_FreeBoundaryAspect. Stores the
    	 -- values for presentation of free boundaries, in other
    	 -- words, boundaries which are not shared . The
    	 -- LineAspect for the free boundaries can be edited. The
    	 -- default values are: Color: Quantity_NOC_GREEN
     	 -- Type of line: Aspect_TOL_SOLID Width: 1.
    	 -- These attributes are used by Prs3d_WFShape.
    is redefined static;

    HasFreeBoundaryAspect (me) returns Boolean from Standard
    ---Purpose: Returns true if the Drawer has a free boundary aspect setting active.
    ---C++: inline
    is static;

    FreeBoundaryDraw(me) returns Boolean from Standard 
	 ---Purpose: returns True if the drawing of the free boundaries is enabled.
    is redefined static;
    

-- Attributes for the wires

    WireAspect (me:mutable) returns LineAspect from Prs3d
	 ---Purpose: Returns a link with Prs3d_Drawer_WireAspect.
    	 -- This method provides wire aspect settings.
    	 -- The LineAspect for wires can be edited. The default values are:
	 --          Color: Quantity_NOC_RED
    	 --          Type of line: Aspect_TOL_SOLID
    	 --          Width: 1.
    	 --          These attributes are used by the following algorithms:
	 --          Prs3d_WFShape
    is redefined static;    

    HasLineAspect (me) returns Boolean from Standard 
	 ---Purpose: Returns true if the Interactive Object has a line
	 -- visualization aspect.
	 ---C++: inline 
  is static;      

    HasWireAspect (me) returns Boolean from Standard 
     	 ---Purpose: Returns true if the Drawer has a wire aspect setting active.
     	 ---C++: inline 
    is static;      

    WireDraw(me) returns Boolean from Standard 
   	 ---Purpose: Returns a link   with Prs3d_Drawer_WireDraw. This
    	 -- method returns true if drawing of wires is enabled.
    	 -- The default setting is true.
    is redefined static;
    

-- Attributes for the unfree boundaries

    UnFreeBoundaryAspect (me:mutable) returns LineAspect from Prs3d
    	 ---Purpose: Returns a link with
    	 -- Prs3d_Drawer_UnFreeBoundaryAspect, which
    	 -- provides settings for shared boundary line aspects.
    	 -- The LineAspect for shared boundaries can be edited.
    	 -- The default values are:
    	 --          Color: Quantity_NOC_YELLOW
    	 --          Type of line: Aspect_TOL_SOLID
    	 --          Width: 1.
	 --          These attributes are used by the following algorithms:
	 --          Prs3d_WFShape
    is redefined static;

    HasUnFreeBoundaryAspect (me) returns Boolean from Standard
    ---Purpose: Returns true if the Drawer has an unfree boundary aspect setting active.
    ---C++: inline
    is static;

    UnFreeBoundaryDraw(me) returns Boolean from Standard 
    	 ---Purpose: Returns True if the drawing of the shared boundaries
    	 -- is enabled. True is the default setting.
    is redefined static;
    

-- 
--  Attributes for the lines.
-- 

    LineAspect(me:mutable) returns LineAspect from Prs3d
    	---Purpose:  Returns a link with Prs3d_Drawer_LineAspect,
    	-- which provides settings for line aspects. These
    	-- settings can be edited. The default values are:         
    	--          Color: Quantity_NOC_YELLOW
    	--          Type of line: Aspect_TOL_SOLID
    	--          Width: 1.
    	-- These attributes are used by the following algorithms:
    	--          Prs3d_Curve
    	--          Prs3d_Line
    	--          Prs3d_HLRShape

    is redefined static;
    
  

    HasTextAspect(me) returns Boolean from Standard
    is static;      
    	---C++: inline     
    TextAspect(me:mutable) returns TextAspect from Prs3d
    --          
    --          Color: Quantity_NOC_YELLOW
    is redefined static;    			    

    LineArrowDraw(me) returns Boolean from Standard 
    	---Purpose: Returns True if the drawing of an arrow at the end of
    	-- each line is enabled. The default setting is False.
    is redefined static;
    
    ArrowAspect(me:mutable) returns ArrowAspect from Prs3d 
    is redefined static;
    
    
-- -- 
--  Attributes for the points
-- 
    PointAspect(me:mutable) returns PointAspect from Prs3d
    	---Purpose:  Returns the point aspect setting. The default values
    	-- are:        Color: Quantity_NOC_YELLOW
	--          Type of marker: Aspect_TOM_PLUS
	--          Scale: 1.
	--          These attributes are used by the following algorithms:
	--          Prs3d_Point
    is redefined static;

    HasPointAspect (me) returns Boolean from Standard 
	---Purpose: Returns true if the Drawer has a point aspect setting active. 
    is static;      
	---C++: inline

    SetVertexDrawMode(me: mutable; theMode: VertexDrawMode from Prs3d)
      ---Purpose: Sets the mode of visualization of vertices by AIS_Shape and helper algorithms.
      -- By default, only isolated vertices not belonging to any face are drawn,
      -- that corresponds to <b>Prs3d_VDM_Isolated</b> mode.
      -- Switching to <b>Prs3d_VDM_Isolated</b> mode makes all shape's vertices visible.
      -- To inherit this parameter from the global drawer instance ("the link") when it is present,
      -- <b>Prs3d_VDM_Inherited</b> value should be used.
    is redefined static;

    VertexDrawMode(me) returns VertexDrawMode from Prs3d
      ---Purpose: Returns the current mode of visualization of vertices of a TopoDS_Shape instance.
    is redefined static;
    
    IsOwnVertexDrawMode(me) returns Boolean from Standard;
      ---Purpose: Returns true if the vertex draw mode is not equal to <b>Prs3d_VDM_Inherited</b>.
      -- This means that individual vertex draw mode value (i.e. not inherited from the global
      -- drawer) is used for a specific interactive object.
      ---C++: inline

--  Attributes for the faces:
--  
    ShadingAspect (me:mutable) returns ShadingAspect from Prs3d
    	---Purpose:
    	-- Returns a link with Prs3d_Drawer_ShadingAspect,
    	-- which provides settings for shading aspects.
    	-- These settings can be edited. The default values are:
	--    Color: Quantity_NOC_YELLOW
    	--          Material: Graphic3d_NOM_BRASS
    	-- hading aspect is obtained through decomposition of
    	-- 3D faces into triangles, each side of each triangle
    	-- being a chord of the corresponding curved edge in
    	-- the face. Reflection of light in each projector
    	-- perspective is then calculated for each of the
    	-- resultant triangular planes.
    is redefined static;

    HasShadingAspect (me) returns Boolean from Standard 
        ---C++: inline 
    	---Purpose: Returns True if the   Drawer has shading aspect active.
    is static;      
        
    ShadingAspectGlobal(me) returns Boolean from Standard
    is redefined static;  
    	---Purpose: Provides the attributes for hidden line removal.


    DrawHiddenLine(me) returns Boolean from Standard 
	---Purpose: Returns Standard_True if the hidden lines are to be drawn.
	--          By default the hidden lines are not drawn.
    is redefined static;
    
    HiddenLineAspect(me:mutable) returns LineAspect from Prs3d
	---Purpose: Returns a link with
    	-- Prs3d_Drawer_HiddenLineAspect, which provides
    	-- settings for hidden line aspects.
    	-- These settings can be edited. The default values are:
    	--          Color: Quantity_NOC_YELLOW
    	--          Type of line: Aspect_TOL_DASH
    	--          Width: 1.
    is redefined static;

    
    SeenLineAspect(me:mutable) returns LineAspect from Prs3d
    	---Purpose: Returns a link with
    	-- Prs3d_Drawer_SeenLineAspect, which provides
    	-- settings for seen line aspects.
    	-- These settings can be edited. The default values are:
    	--          Color: Quantity_NOC_YELLOW
    	--          Type of line: Aspect_TOL_SOLID
    	--          Width: 1.
    is redefined static;
    
  
    HasPlaneAspect(me) returns Boolean from Standard;
    	---C++: inline

    PlaneAspect(me:mutable) returns PlaneAspect from Prs3d
    is redefined static;
    	---Purpose:
    	-- Returns a link with Prs3d_Drawer_PlaneAspect.
    	-- This method provides settings for the appearance of planes.


    VectorAspect(me:mutable) returns LineAspect from Prs3d
    	---Purpose: Returns a link with Prs3d_Drawer_VectorAspect,
    	-- which provides settings for the appearance of vectors.
    	-- These settings can be edited. The default values are:
    	--          Color: Quantity_NOC_SKYBLUE
    	--          Type of line: Aspect_TOL_SOLID Width: 1.
    is redefined static;
    
    SetFaceBoundaryDraw (me           : mutable;
                         theIsEnabled : Boolean from Standard)
    is redefined static;
        ---Purpose: Enables or disables drawing of face boundaries for shading presentations.
        -- The method sets drawing flag owned by the drawer that will be used during
        -- visualization instead of the one set in link.
        -- theIsEnabled is a boolean flag indicating whether the face boundaries should be
        -- drawn or not.

    IsFaceBoundaryDraw (me) returns Boolean from Standard
    is redefined static;
        ---Purpose: Checks whether the drawing of face boundaries is enabled or not.

    SetFaceBoundaryAspect (me        : mutable;
                           theAspect : LineAspect from Prs3d)
    is redefined static;
        ---Purpose: Sets line aspect for face boundaries.
        -- The method sets line aspect owned by the drawer that will be used during
        -- visualization instead of the one set in link.
        -- theAspect is the line aspect that determines the look of the face boundaries.

    FaceBoundaryAspect (me : mutable) returns LineAspect from Prs3d
    is redefined static;
        ---Purpose: Returns line aspect of face boundaries.

    IsOwnFaceBoundaryDraw (me) returns Boolean from Standard
    is static;
        ---Purpose: Returns true if the drawer has its own attribute for 
        -- "draw face boundaries" flag that overrides the one in the link.
        ---C++: inline

    IsOwnFaceBoundaryAspect (me) returns Boolean from Standard
    is static;
        ---Purpose: Returns true if the drawer has its own attribute for 
        -- face boundaries aspect that overrides the one in the link.
        ---C++: inline
--
--  Attributes for the presentation of a Datum.
--  

    HasDatumAspect(me) returns Boolean from Standard;
    	---C++: inline 

    DatumAspect(me:mutable) returns DatumAspect from Prs3d
    	---Purpose: Returns a link with Prs3d_Drawer_DatumAspect,
    	-- which provides settings for the appearance of datums.
    	-- These settings can be edited. The default values for
    	-- the three axes are:
    	--          Color: Quantity_NOC_PEACHPUFF
    	--          Type of line: Aspect_TOL_SOLID Width: 1.
    is redefined static;

--
--  Attributes for the presentation of a dimensions.
--  

    DimensionAspect (me : mutable) returns DimensionAspect from Prs3d is redefined static;
    ---Purpose: Returns a link with Prs3d_Drawer_DimensionAspect,
    -- which provides settings for the appearance of dimensions.

    HasDimensionAspect (me) returns Boolean from Standard is static;
    ---C++: inline
    -- Purpose: Returns true if the Drawer has a dimension aspect setting active.

    SetDimLengthModelUnits (me: mutable; theUnits : AsciiString from TCollection) is redefined static;
    ---Purpose: Sets dimension length model units for computing of dimension presentation.

    SetDimAngleModelUnits (me: mutable; theUnits : AsciiString from TCollection) is redefined static;
    ---Purpose: Sets dimension angle model units for computing of dimension presentation.

    DimAngleModelUnits (me) returns AsciiString from TCollection is redefined static;
    ---Purpose: Returns angle model units for the dimension presentation.
    ---C++: return const &

    DimLengthModelUnits (me) returns AsciiString from TCollection is redefined static;
    ---Purpose: Returns length model units for the dimension presentation.
    ---C++: return const &

    SetDimLengthDisplayUnits (me: mutable; theUnits : AsciiString from TCollection) is redefined static;
    ---Purpose: Sets length units in which value for dimension presentation is displayed.

    SetDimAngleDisplayUnits (me: mutable; theUnits : AsciiString from TCollection) is redefined static;
    ---Purpose: Sets angle units in which value for dimension presentation is displayed.

    DimLengthDisplayUnits (me) returns AsciiString from TCollection is redefined static;
    ---Purpose: Returns length units in which dimension presentation is displayed.
    ---C++: return const &

    DimAngleDisplayUnits (me) returns AsciiString from TCollection is redefined static;
    ---Purpose: Returns angle units in which dimension presentation is displayed.
    ---C++: return const &

-- Attributes for the sections

    SectionAspect (me:mutable) returns LineAspect from Prs3d
    	---Purpose: Returns a link with Prs3d_Drawer_SectionAspect,
    	-- which provides settings for wires which highlight sections.
    	-- The LineAspect for the wire can be edited.
    	-- The default values are:
    	-- Color: Quantity_NOC_ORANGE
    	-- Type of line: Aspect_TOL_SOLID
    	-- Width: 1.
	-- These attributes are used by the following algorithms:
	-- Prs3d_WFShape
    is redefined static;    

    Link(me:mutable) returns any Drawer from Prs3d
    is static;
	---C++: return const&

    HasLink(me) returns Boolean from Standard
    is static;
 	---C++: inline

    Link (me:mutable; aDrawer: Drawer from Prs3d)     
    is static;
    	---C++: inline

    
    ClearLocalAttributes(me:mutable) is virtual;    
    	---Purpose: Removes attributes stored in a Local Context.    
    
    WasLastLocal(me) returns Boolean from Standard;
        ---C++: inline
    	---Purpose: Returns true if the last called attribute was local; false if it was global.
    
    HasLocalAttributes(me) returns Boolean from Standard;
        ---C++: inline
    	---Purpose:
    	-- Returns true if a Local Context has stored attributes
    	-- for Interactive Objects.

fields

    myLink                           : Drawer from Prs3d;
    hasLocalAttributes               : Boolean from Standard;		

    myhasOwnDeviationCoefficient     : Boolean from Standard;
    myOwnDeviationCoefficient        : Real from Standard;
    myPreviousDeviationCoefficient   : Real from Standard;

    myhasOwnHLRDeviationCoefficient  : Boolean from Standard;
    myOwnHLRDeviationCoefficient     : Real from Standard;
    myPreviousHLRDeviationCoefficient: Real from Standard;

    myhasOwnDeviationAngle           : Boolean from Standard;
    myOwnDeviationAngle              : Real from Standard;
    myPreviousDeviationAngle         : Real from Standard;

    myhasOwnHLRDeviationAngle        : Boolean from Standard;
    myOwnHLRDeviationAngle           : Real from Standard; 
    myPreviousHLRDeviationAngle      : Real from Standard;
    myHasOwnFaceBoundaryDraw         : Boolean from Standard;

    myHasOwnDimLengthModelUnits      : Boolean from Standard;
    myHasOwnDimLengthDisplayUnits    : Boolean from Standard;
    myHasOwnDimAngleModelUnits      : Boolean from Standard;
    myHasOwnDimAngleDisplayUnits    : Boolean from Standard;

end Drawer;
 

