-- Created on: 1991-10-10
-- Created by: Jean Claude VAUTHIER
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class CircleToBSplineCurve    from Convert   inherits ConicToBSplineCurve

        --- Purpose :
        --  This algorithm converts a circle into a rational B-spline curve.
        --  The circle is a Circ2d from package gp and its parametrization is :
        --  P (U) = Loc + R * (Cos(U) * Xdir + Sin(U) * YDir) where Loc is the
        --  center of the circle Xdir and Ydir are the normalized directions
        --  of the local cartesian coordinate system of the circle.
        --  The parametrization range for the circle is U [0, 2Pi].
        --  
        --- Warnings :
        --  The parametrization range for the B-spline curve is not [0, 2Pi].
        --  
        --- KeyWords :
        --  Convert, Circle, BSplineCurve, 2D .


uses Circ2d               from gp,
     ParameterisationType from Convert 

raises DomainError from Standard

is

  Create (C : Circ2d;
          Parameterisation : ParameterisationType from Convert 
    	    = Convert_TgtThetaOver2) 
  returns CircleToBSplineCurve;
        --- Purpose :
        --  The equivalent B-spline curve has the same orientation
        --  as the circle C.


  Create (C : Circ2d; U1, U2 : Real ;
    Parameterisation : ParameterisationType from Convert 
    = Convert_TgtThetaOver2)     
    returns CircleToBSplineCurve 
        --- Purpose : 
        --  The circle C is limited between the parametric values U1, U2
        --  in radians. U1 and U2 [0.0, 2*Pi] .
        --  The equivalent B-spline curve is oriented from U1 to U2 and has
        --  the same orientation as the circle C.
     raises DomainError;
        --- Purpose :
        --  Raised if U1 = U2 or U1 = U2 + 2.0 * Pi


end CircleToBSplineCurve;
  
