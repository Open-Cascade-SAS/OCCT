-- Created on: 2002-12-12
-- Created by: data exchange team
-- Copyright (c) 2002-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class DataEnvironment from StepRepr
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity DataEnvironment

uses
    HAsciiString from TCollection,
    HArray1OfPropertyDefinitionRepresentation from StepRepr

is
    Create returns DataEnvironment from StepRepr;
	---Purpose: Empty constructor

    Init (me: mutable; aName: HAsciiString from TCollection;
                       aDescription: HAsciiString from TCollection;
                       aElements: HArray1OfPropertyDefinitionRepresentation from StepRepr);
	---Purpose: Initialize all fields (own and inherited)

    Name (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Name
    SetName (me: mutable; Name: HAsciiString from TCollection);
	---Purpose: Set field Name

    Description (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Description
    SetDescription (me: mutable; Description: HAsciiString from TCollection);
	---Purpose: Set field Description

    Elements (me) returns HArray1OfPropertyDefinitionRepresentation from StepRepr;
	---Purpose: Returns field Elements
    SetElements (me: mutable; Elements: HArray1OfPropertyDefinitionRepresentation from StepRepr);
	---Purpose: Set field Elements

fields
    theName: HAsciiString from TCollection;
    theDescription: HAsciiString from TCollection;
    theElements: HArray1OfPropertyDefinitionRepresentation from StepRepr;

end DataEnvironment;
