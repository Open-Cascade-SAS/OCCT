-- Created on: 2002-11-19
-- Created by: Vladimir ANIKIN
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ApplicationDelta from TDocStd inherits TShared from MMgt

uses

	SequenceOfDocument from TDocStd,
	ExtendedString from TCollection,
	OStream from Standard

is

	Create returns ApplicationDelta from TDocStd;

	GetDocuments(me : mutable)
	returns SequenceOfDocument from TDocStd;
	---C++: return &
	---C++: inline

	GetName(me)
	returns ExtendedString from TCollection;
	---C++: return const &
	---C++: inline

    	SetName(me : mutable;
	    	theName : ExtendedString from TCollection);
	---C++: inline

	Dump(me;
	     anOS : in out OStream from Standard);

fields

	myDocuments : SequenceOfDocument from TDocStd;
	myName      : ExtendedString from TCollection;

end ApplicationDelta;
