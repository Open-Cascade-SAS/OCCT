-- Created on: 1996-01-29
-- Created by: PLOTNIKOV Eugeny
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class FontMapEntry from WNT inherits TShared from MMgt

	---Purpose: Defines correspondence between FontMapEntry from
        --          Aspect and Windows NT font handle. Also, provides
        --          some optimizations due to rotation, italics & underlining
        --          of fonts. Each font can be reffered by its name which
        --          is a character string. The format of the string takes
        --          after format of font name of X window system but there
        --          are some differences. The font name string format is:
        --          "h-w-e-o-wgt-i-u-so-cs-op-cp-q-pf-face".
        --           ^ ^ ^ ^  ^  ^ ^ ^  ^  ^  ^  ^ ^   ^
        --           | | | |  |  | | |  |  |  |  | |   |
        --           | | | |  |  | | |  |  |  |  | |   +- name of the typeface
        --           | | | |  |  | | |  |  |  |  | |      (Courier, Arial ...)
        --           | | | |  |  | | |  |  |  |  | +- pitch and family
        --           | | | |  |  | | |  |  |  |  +- quality
        --           | | | |  |  | | |  |  |  +- clip precision
        --           | | | |  |  | | |  |  +- out precision
        --           | | | |  |  | | |  +- character set
        --           | | | |  |  | | +- strike out
        --           | | | |  |  | +- underline
        --           | | | |  |  +- italic
        --           | | | |  +- weight
        --           | | | +- orientation
        --           | | +- escapement
        --           | +- width
        --           +- height
        --           Wildcarding is allowed by specifying '*' sign. This means
        --           a default value for parameter.
        --  Example: "13-8-*-*-400-*-*-*-255-1-2-*-25-courier".
        --          For more detail information see Microsoft Windows manual.
        --  Warning: Windows can output rotated text only if the selected for
        --          drawing font is True Type.
 uses

    Handle     from Aspect,
    LogFont    from WNT,
    Dword      from WNT,
    Factor     from Quantity,
    PlaneAngle from Quantity

 raises

    FontMapEntryDefinitionError from WNT

 is

    Create ( aFontName : CString from Standard )
     returns mutable FontMapEntry from WNT
    	---Purpose: Creates a class and loads font.
        --  Warning: Windows finds the real font that most closely matches
        --          the request. In doing so, it uses a
        --          "font-mapping-algorythm". So it is possible that loaded
        --          font differs from font in the request.
    	--  Trigger: Raises if font loading failed.
     raises FontMapEntryDefinitionError from WNT;

    Destroy ( me : mutable ) is virtual;
	---Level:   Public
	---Purpose: Destroys all ressources attached to the FontMapEntry
    	---C++:     alias ~

    HFont ( me ) returns Handle from Aspect;
	---Level:   Public
	---Purpose: Returns handle of the font.

    SetAttrib (
     me     : mutable;
     aFlags : Dword   from WNT;
     aData  : Address from Standard;
     aRepl  : Boolean from Standard = Standard_False
    ) returns Handle from Aspect is static;
	---Level:   Internal
	---Purpose: Sets certain attributes ( italics etc. ) for font.
        --  Warning: If <aRepl> is True then creates a new handle for font.
        --          In this case calling routine MUST DELETE THE FONT ITSELF
        --          WHEN THE FONT BECOME NO LONGER NEEDED.

    SetSlant ( me : mutable; aSlant : PlaneAngle from Quantity )
     returns PlaneAngle from Quantity is static;
     	---Level:   Internal
    	---Purpose: Sets the font's slant and returns a previous one.
    	---C++:     inline

    SetScale ( me : mutable; aScale : Factor from Quantity )
     returns Factor from Quantity is static; 
    	---Level:   Internal
    	---Purpose: Sets the font's scale and returns a previous one.
    	---C++:     inline

    Slant ( me )
     returns PlaneAngle from Quantity is static;
     	---Level:   Internal
     	---Purpose: Returns value of the font's slant.
     	---C++:     inline

    Scale ( me )
     returns Factor from Quantity is static;
     	---Level:   Internal
     	---Purpose: Returns value of the font's scale.
     	---C++:     inline

    LogFont ( me )
     returns Address from Standard is static;
     	---Level:   Internal
     	---Purpose: Returns pointer to LogFont structure.
     	---C++:     inline

 fields

    myLogFont : LogFont    from WNT      is protected;
    myHandle  : Handle     from Aspect   is protected;
    myScale   : Factor     from Quantity is protected;
    mySlant   : PlaneAngle from Quantity is protected;

 friends
 
    class WDriver from WNT,
    class DDriver from WNT

end FontMapEntry;
