-- Created on: 1999-06-30
-- Created by: Sergey ZARITCHNY
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

private class Translator from TNaming

	---Purpose: 

uses
    Shape  from  TopoDS, 
    DataMapOfShapeShape from  TopTools, 
    IndexedDataMapOfTransientTransient  from TColStd

is
 
    Create  returns  Translator  from  TNaming; 
     
    Add(me  : in  out;  aShape  :  Shape  from  TopoDS); 
     
    Perform (me  :  in  out); 
     
    IsDone(me) 
    	returns  Boolean  from  Standard;
     
    Copied(me;  aShape  :  Shape  from  TopoDS)   
    returns  Shape   from  TopoDS;  
    ---Purpose: returns copied  shape
    ---C++  :  return  const 
     
    Copied(me)   
    returns  DataMapOfShapeShape   from  TopTools; 
     ---C++  :  return  const&
     ---Purpose: returns  DataMap  of  results;  (shape <-> copied  shape)
    DumpMap(me;  isWrite  :  Boolean  from  Standard  =  Standard_False); 
    
fields  

    myIsDone           : Boolean       from Standard;
    myMap              : IndexedDataMapOfTransientTransient  from TColStd;  
    myDataMapOfResults : DataMapOfShapeShape  from  TopTools;
--    myListOfShape    : ListOfShape   from  TopTools;
--    myListOfResult   : ListOfShape   from  TopTools;
    
end Translator;
