-- Created on: 1997-02-06
-- Created by: Denis PASCAL
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Integer from TDataStd inherits Attribute from TDF

	---Purpose:  The basis to define an integer attribute.

uses Attribute       from TDF,
     Label           from TDF,
     GUID            from Standard,
     Integer         from Standard,
     RelocationTable from TDF

is 

    ---Purpose: class methods
    --          =============

    GetID (myclass)   
        ---C++: return const & 
	---Purpose: Returns the GUID for integers.  
    returns GUID from Standard;

    Set (myclass; label : Label from TDF; value : Integer from Standard)
    ---Purpose: Finds, or creates, an Integer attribute and sets <value>
    --          the Integer  attribute is returned.
    returns Integer from TDataStd;

    ---Purpose: Integer methods
    --          ===============
    
    Set (me : mutable; V : Integer from Standard);
    
    Get (me)
    returns Integer from Standard;
    ---Purpose: Returns the integer value contained in the attribute.
    IsCaptured(me) returns Boolean;
	---Purpose: Returns True if there is a reference on the same label

    ---Category: methodes de TDF_Attribute
    --           =========================
    
    ID (me)
    	---C++: return const & 
    returns GUID from Standard;

    Restore (me: mutable; With : Attribute from TDF);

    NewEmpty (me)
    returns Attribute from TDF;

    Paste (me; Into : Attribute from TDF;
	       RT   : RelocationTable from TDF);    

    Dump(me; anOS : in out OStream from Standard)
    	returns OStream from Standard
    	is redefined;
	---C++: return &


    Create
    returns Integer from TDataStd;    


fields

    myValue : Integer from Standard;

end Integer;
