-- Created on: 1995-09-18
-- Created by: Bruno DUMORTIER
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MakeOffset from BRepOffsetAPI inherits MakeShape from BRepBuilderAPI

	---Purpose: Describes algorithms for offsetting wires from a set of
    	-- wires contained in a planar face.
    	-- A MakeOffset object provides a framework for:
    	-- - defining the construction of an offset,
    	-- - implementing the construction algorithm, and
    	-- - consulting the result. 

uses
    Shape             from TopoDS,
    Wire              from TopoDS,
    Face              from TopoDS,
    ListOfShape       from TopTools,
    OffsetWire        from BRepFill, 
    ListOfOffsetWire  from BRepFill,
    JoinType          from GeomAbs
    
    
raises
    NotDone from StdFail
    
is
    Create returns MakeOffset from BRepOffsetAPI;
    	---Purpose: Constructs an algorithm for creating an empty offset
    Create( Spine : Face from TopoDS;
    	    Join  : JoinType from GeomAbs = GeomAbs_Arc)
    returns MakeOffset from BRepOffsetAPI;
    	---Purpose: Constructs an algorithm for creating an algorithm
    	-- to build parallels to the spine Spine   
    Init( me    : in out;
    	  Spine : Face     from TopoDS; 
    	  Join  : JoinType from GeomAbs  =  GeomAbs_Arc)
	---Purpose: Initializes the algorithm to construct parallels to the spine Spine.
    	-- Join defines the type of parallel generated by the
    	-- salient vertices of the spine. The default type is
    	-- GeomAbs_Arc where the vertices generate sections
    	-- of a circle. At present, this is the only construction type implemented.
    is static;
    
    Create( Spine : Wire from TopoDS;
    	    Join  : JoinType from GeomAbs = GeomAbs_Arc)
    returns MakeOffset from BRepOffsetAPI;
    
    Init( me    : in out;
    	  Join  : JoinType from GeomAbs  =  GeomAbs_Arc)
	---Purpose: Initialize the evaluation of Offseting.
    is static;

    AddWire (me : in out;
    	     Spine : Wire from TopoDS)
        ---Purpose: Initializes the algorithm to construct parallels to the wire Spine.
    is static;

    Perform (me : in out; 
    	     Offset : Real from Standard;
    	     Alt    : Real from Standard = 0.0)
	---Purpose:  Computes a parallel to the spine at distance Offset and
    	-- at an altitude Alt from the plane of the spine in relation
    	-- to the normal to the spine.
    	-- Exceptions: StdFail_NotDone if the offset is not built.
    raises
    	NotDone from StdFail
    is static;

	
    Build(me : in out)
    is redefined;
	---Purpose: Builds the resulting shape (redefined from MakeShape).
	---Level: Public    

    Generated  (me: in out; S : Shape from TopoDS)
    	---Purpose: returns a list of the created shapes
    	--          from the shape <S>.
    	---C++:     return const &
	---Level: Public
    returns ListOfShape from TopTools
    is redefined;


fields

    myIsInitialized : Boolean          from Standard;
    myLastIsLeft    : Boolean          from Standard;
    myJoin          : JoinType         from GeomAbs;	
    myFace          : Face             from TopoDS;
    myWires         : ListOfShape      from TopTools;   
    myLeft          : ListOfOffsetWire from BRepFill;
    myRight         : ListOfOffsetWire from BRepFill;
    
end MakeOffset;
