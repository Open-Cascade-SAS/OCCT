-- Created on: 1993-10-27
-- Created by: Jean-Louis FRENKEL
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ToolShadedShape from StdPrs inherits ShapeTool from BRepMesh 

uses
    Shape         from TopoDS,
    Face          from TopoDS,
    Array1OfDir   from TColgp,
    Connect       from Poly,
    Triangulation from Poly,
    Location      from TopLoc
is

    IsClosed(myclass; aShape: Shape from TopoDS) returns Boolean from Standard; 
    
    Triangulation(myclass; aFace: Face from TopoDS;
    	    	    	   loc  : out Location from TopLoc) 
    returns Triangulation from Poly;
    
    Normal(myclass; aFace: Face            from TopoDS;
    	    	    PC   : in out Connect  from Poly;
		    Nor  : out Array1OfDir from TColgp);
    
end ToolShadedShape from StdPrs;
