-- Created on: 1997-08-06
-- Created by: Philippe MANGIN
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

private  class QuasiAngularConvertor from GeomFill 

	---Purpose: To convert circular section in QuasiAngular Bezier
 	--          form   

uses
    Matrix from math, 
    Vector from  math,
    Pnt from gp,
    Vec from gp,  
    Array1OfReal from  TColStd,
    Array1OfPnt  from TColgp,
    Array1OfVec  from TColgp

raises NotDone from StdFail

is
    Create returns QuasiAngularConvertor from GeomFill;
    
    Initialized(me) 
    ---Purpose: say if <me> is Initialized
    returns Boolean;
    
    Init(me: in out);
    
    Section(me  :  in  out;
    	    FirstPnt : Pnt from gp;
	    Center   : Pnt from gp;
	    Dir      : Vec from gp;
	    Angle    : Real from Standard;
            Poles    : out Array1OfPnt  from TColgp; 
            Weights  : out Array1OfReal from TColStd);
	    
    Section(me:  in  out;
    	    FirstPnt  : Pnt from gp;
	    DFirstPnt : Vec from gp;
	    Center    : Pnt from gp;
	    DCenter   : Vec from gp;
	    Dir       : Vec from gp;
	    DDir      : Vec from gp;
	    Angle     : Real from Standard;
	    DAngle    : Real from Standard;
            Poles     : out Array1OfPnt   from TColgp;
            DPoles    : out Array1OfVec   from TColgp; 
            Weights   : out Array1OfReal from TColStd; 
            DWeights  : out Array1OfReal from TColStd);
	    
     Section(me  :  in  out;
    	    FirstPnt  : Pnt from gp;
	    DFirstPnt : Vec from gp;
	    D2FirstPnt: Vec from gp;
	    Center    : Pnt from gp;
	    DCenter   : Vec from gp;
	    D2Center  : Vec from gp;
	    Dir       : Vec from gp;
	    DDir      : Vec from gp;
	    D2Dir     : Vec from gp;
	    Angle     : Real from Standard;
	    DAngle    : Real from Standard;
	    D2Angle   : Real from Standard;
            Poles     : out Array1OfPnt   from TColgp;
            DPoles    : out Array1OfVec   from TColgp;
            D2Poles   : out Array1OfVec   from TColgp; 
            Weights   : out Array1OfReal from TColStd; 
            DWeights  : out Array1OfReal from TColStd; 
            D2Weights : out Array1OfReal from TColStd);  	    
 
fields  
    myinit : Boolean from Standard;
    B       : Matrix from math;  
    Px,  Py,  W,  Vx,  Vy, Vw : Vector  from  math; 
end QuasiAngularConvertor;
