-- Created on: 1993-09-29
-- Created by: Isabelle GRIGNON
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class GeomTool from BRepMesh
       	---Purpose: 

uses 
     Pnt                  from gp,
     Vec                  from gp,
     Dir                  from gp,
     Pnt2d                from gp,
     IsoType              from GeomAbs,
     TangentialDeflection from GCPnts,
     Curve                from BRepAdaptor,
     HSurface             from BRepAdaptor
     


is

    Create (C : in out Curve from BRepAdaptor;
            Ufirst,Ulast,AngDefl, Deflection : Real;
            nbpointsmin: Integer = 2)
    	returns GeomTool;
    
    Create (S        : HSurface from BRepAdaptor;
            ParamIso : Real;
            Type     : IsoType  from GeomAbs;
    	    Ufirst,Ulast,AngDefl,Deflection : Real;
    	    nbpointsmin: Integer = 2) returns GeomTool;

    AddPoint(me : in out; thePnt : in Pnt from gp;
                          theParam : in Real;
                          theIsReplace : in Boolean = Standard_True)
    returns Integer from Standard;
    ---Purpose: Add point to already calculated points (or replace existing)
    --          Returns index of new added point
    --           or founded with parametric tolerance (replaced if theIsReplace is true)
	    
    NbPoints(me) returns Integer from Standard;
    
    Value(me; IsoParam : Real ; Index : Integer ; 
          W : out Real; P : out Pnt from gp; UV : out Pnt2d from gp);
	      
    Value(me;C : Curve from BRepAdaptor;
             S : HSurface from BRepAdaptor;
             Index : Integer from Standard; 
    	     W : out Real; P : out Pnt from gp; UV : out Pnt2d from gp);    
	
    D0(myclass; F : HSurface  from BRepAdaptor;U,V : Real; P : out Pnt);
	
    Normal(myclass; F : HSurface from BRepAdaptor;U,V : Real ; P : out Pnt from gp; 
    	    	    	    	    	   Nor : out  Dir from gp)
    returns Boolean from Standard;
    ---Purpose: return false if the normal can not be computed 

fields

pnts                : TangentialDeflection from GCPnts;
parametric          : IsoType           from GeomAbs;

end GeomTool;
