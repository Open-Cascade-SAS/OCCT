-- Created on: 1993-01-11
-- Created by: CKY / Contract Toubro-Larsen ( Arun MENON )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class RegionRestriction from IGESAppli  inherits IGESEntity

        ---Purpose: defines RegionRestriction, Type <406> Form <2>
        --          in package IGESAppli
        --          Defines regions to set an application's restriction
        --          over a region.

uses  Integer  -- no one specific type

is

        Create returns mutable RegionRestriction;

        -- Specific Methods pertaining to the class

        Init (me         : mutable;
              nbPropVal  : Integer;
              aViasRest  : Integer;
              aCompoRest : Integer;
              aCktRest   : Integer);
        ---Purpose : This method is used to set the fields of the class
        --           RegionRestriction
        --       - nbPropVal  : Number of property values, always = 3
        --       - aViasRest  : Electrical Vias restriction
        --       - aCompoRest : Electrical components restriction
        --       - aCktRest   : Electrical circuitry restriction

        NbPropertyValues (me) returns Integer;
        ---Purpose : is always 3

        ElectricalViasRestriction (me) returns Integer;
        ---Purpose : returns the Electrical vias restriction
        -- is 0, 1 or 2

        ElectricalComponentRestriction (me) returns Integer;
        ---Purpose : returns the Electrical components restriction
        -- is 0, 1 or 2

        ElectricalCktRestriction (me) returns Integer;
        ---Purpose : returns the Electrical circuitry restriction
        -- is 0, 1 or 2

fields

--
-- Class    : IGESAppli_RegionRestriction
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class RegionRestriction.
--
-- Reminder : A RegionRestriction instance is defined by :
--            - Number of property values (always = 3)
--            - Electrical vias restriction
--            - Electrical components restriction
--            - Electrical circuitry restriction

        theNbPropertyValues  : Integer;
        theElectViasRestrict : Integer;
        theElectCompRestrict : Integer;
        theElectCktRestrict  : Integer;

end RegionRestriction;
