-- Created on: 1993-01-09
-- Created by: CKY / Contract Toubro-Larsen ( SIVA )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class SphericalSurface from IGESSolid  inherits IGESEntity

        ---Purpose: defines SphericalSurface, Type <196> Form Number <0,1>
        --          in package IGESSolid
        --          Spherical surface is defined by a center and radius.
        --          In case of parametrised surface an axis and a
        --          reference direction is provided.

uses

        Point           from IGESGeom,
        Direction       from IGESGeom,
        Pnt             from gp

is

        Create returns mutable SphericalSurface;

        -- Specific Methods pertaining to the class

        Init (me      : mutable;
              aCenter : Point;
              aRadius : Real;
              anAxis  : Direction;
              aRefdir : Direction);
        ---Purpose : This method is used to set the fields of the class
        --           SphericalSurface
        --       - aCenter : the coordinates of the center point
        --       - aRadius : value of radius
        --       - anAxis  : the direction of the axis
        --                   Null in case of Unparametrised surface
        --       - aRefdir : the reference direction
        --                   Null in case of Unparametrised surface

        Center(me) returns Point;
        ---Purpose : returns the center of the spherical surface

        TransformedCenter(me) returns Pnt;
        ---Purpose : returns the center of the spherical surface after applying
        -- TransformationMatrix

        Radius(me) returns Real;
        ---Purpose : returns the radius of the spherical surface

        Axis(me) returns Direction;
        ---Purpose : returns the direction of the axis (Parametrised surface)
        -- Null is returned if the surface is not parametrised

        ReferenceDir(me) returns Direction;
        ---Purpose : returns the reference direction (Parametrised surface)
        -- Null is returned if the surface is not parametrised

        IsParametrised(me) returns Boolean;
        ---Purpose : Returns True if the surface is parametrised, else False

fields

--
-- Class    : IGESSolid_SphericalSurface
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class SphericalSurface.
--
-- Reminder : A SphericalSurface instance is defined by :
--            the center point coordinates (Center), a radius (Radius).
--            In case of Parametrised surface, the direction of the axis
--            (Axis) and a reference direction (RefDir) is given.
--

        theCenter  : Point;
            --  the center of the spherical surface

        theRadius  : Real;
            --  the radius of the spherical surface

        theAxis    : Direction;
            -- the direction of the axis (Parametrised surface)

        theRefDir  : Direction;
            -- the reference direction (Parametrised surface)

end SphericalSurface;
