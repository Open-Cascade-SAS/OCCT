-- Created on: 2008-10-31
-- Created by: EPA
-- Copyright (c) 2008-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class FaceAttribute from BRepMesh inherits TShared from MMgt

    ---Purpose: auxiliary class for FastDiscret and FastDiscretFace classes

uses    
    Real          from Standard,
    Address       from Standard,
    ClassifierPtr from BRepMesh

is 

    Create returns mutable FaceAttribute from BRepMesh;

    GetDefFace(me:mutable) returns Real;
       ---C++: return &
       ---C++: inline    

    GetUMin(me:mutable) returns Real;
       ---C++: return &
       ---C++: inline

    GetVMin(me:mutable) returns Real;
       ---C++: return &
       ---C++: inline

    GetUMax(me:mutable) returns Real;
       ---C++: return &
       ---C++: inline

    GetVMax(me:mutable) returns Real;
       ---C++: return &
       ---C++: inline

    GetDeltaX(me:mutable) returns Real;
       ---C++: return &
       ---C++: inline

    GetDeltaY(me:mutable) returns Real;
       ---C++: return &
       ---C++: inline

    GetMinX(me:mutable) returns Real;
       ---C++: return &
       ---C++: inline

    GetMinY(me:mutable) returns Real;
       ---C++: return &
       ---C++: inline
       
    GetClassifier(me:mutable) returns ClassifierPtr from BRepMesh;
       ---C++: return &
       ---C++: inline

fields  
    mydefface   : Real          from Standard;
    myumin      : Real          from Standard;
    myumax      : Real          from Standard;
    myvmin      : Real          from Standard;
    myvmax      : Real          from Standard;
    mydeltaX    : Real          from Standard;
    mydeltaY    : Real          from Standard;
    myminX      : Real          from Standard;
    myminY      : Real          from Standard;
    myclassifier: ClassifierPtr from BRepMesh;

end FaceAttribute;
