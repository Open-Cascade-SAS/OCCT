-- File:	StepFEA_FeaParametricPoint.cdl
-- Created:	Thu Dec 12 17:51:06 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class FeaParametricPoint from StepFEA
inherits Point from StepGeom

    ---Purpose: Representation of STEP entity FeaParametricPoint

uses
    HAsciiString from TCollection,
    HArray1OfReal from TColStd

is
    Create returns FeaParametricPoint from StepFEA;
	---Purpose: Empty constructor

    Init (me: mutable; aRepresentationItem_Name: HAsciiString from TCollection;
                       aCoordinates: HArray1OfReal from TColStd);
	---Purpose: Initialize all fields (own and inherited)

    Coordinates (me) returns HArray1OfReal from TColStd;
	---Purpose: Returns field Coordinates
    SetCoordinates (me: mutable; Coordinates: HArray1OfReal from TColStd);
	---Purpose: Set field Coordinates

fields
    theCoordinates: HArray1OfReal from TColStd;

end FeaParametricPoint;
