-- File:        OrientedOpenShell.cdl
-- Created:     Mon Dec  4 12:02:28 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWOrientedOpenShell from RWStepShape

	---Purpose : Read & Write Module for OrientedOpenShell

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     OrientedOpenShell from StepShape,
     EntityIterator from Interface

is

	Create returns RWOrientedOpenShell;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable OrientedOpenShell from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : OrientedOpenShell from StepShape);

	Share(me; ent : OrientedOpenShell from StepShape; iter : in out EntityIterator);

end RWOrientedOpenShell;
