-- File:        Curve.cdl
-- Created:     Mon Dec  4 12:02:25 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWCurve from RWStepGeom

	---Purpose : Read & Write Module for Curve

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     Curve from StepGeom

is

	Create returns RWCurve;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable Curve from StepGeom);

	WriteStep (me; SW : in out StepWriter; ent : Curve from StepGeom);

end RWCurve;
