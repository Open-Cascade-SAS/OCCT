-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class CompositeCurveSegment from StepGeom 

inherits TShared from MMgt

uses

	TransitionCode from StepGeom, 
	Boolean from Standard, 
	Curve from StepGeom
is

	Create returns mutable CompositeCurveSegment;
	---Purpose: Returns a CompositeCurveSegment

	Init (me : mutable;
	      aTransition : TransitionCode from StepGeom;
	      aSameSense : Boolean from Standard;
	      aParentCurve : mutable Curve from StepGeom) is virtual;

	-- Specific Methods for Field Data Access --

	SetTransition(me : mutable; aTransition : TransitionCode);
	Transition (me) returns TransitionCode;
	SetSameSense(me : mutable; aSameSense : Boolean);
	SameSense (me) returns Boolean;
	SetParentCurve(me : mutable; aParentCurve : mutable Curve);
	ParentCurve (me) returns mutable Curve;

fields

	transition : TransitionCode from StepGeom; -- an Enumeration
	sameSense : Boolean from Standard;
	parentCurve : Curve from StepGeom;

end CompositeCurveSegment;
