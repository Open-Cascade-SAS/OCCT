-- Created on: 1993-01-09
-- Created by: CKY / Contract Toubro-Larsen (Kiran)
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class BoundedSurface from IGESGeom  inherits IGESEntity

        ---Purpose: defines BoundedSurface, Type <143> Form <0>
        --          in package IGESGeom
        --          A bounded surface is used to communicate trimmed
        --          surfaces. The surface and trimming curves are assumed
        --          to be represented parametrically.

uses

        Boundary            from IGESGeom,
        HArray1OfBoundary   from IGESGeom

raises OutOfRange

is

        Create returns mutable BoundedSurface;

        -- Specific Methods pertaining to the class

        Init (me        : mutable;
              aType     : Integer;
              aSurface  : IGESEntity;
              allBounds : HArray1OfBoundary);
        ---Purpose : This method is used to set the fields of the class
        --           BoundedSurface
        --       - aType     : Type of bounded surface representation
        --       - aSurface  : Surface entity to be bounded
        --       - allBounds : Array of boundary entities

        RepresentationType (me) returns Integer;
        ---Purpose : returns the type of Bounded surface representation
        -- 0 = The boundary entities may only reference model space curves
        -- 1 = The boundary entities may reference both model space curves
        --     and associated parameter space curve representations

        Surface (me) returns IGESEntity;
        ---Purpose : returns the bounded surface

        NbBoundaries (me) returns Integer;
        ---Purpose : returns the number of boundaries

        Boundary (me; Index : Integer) returns Boundary
        raises OutOfRange;
        ---Purpose : returns boundary entity
        -- raises exception if Index <= 0 or Index > NbBoundaries()

fields

--
-- Class    : IGESGeom_BoundedSurface
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class BoundedSurface.
--
-- Reminder : A BoundedSurface instance is defined by :
--            The type of bounded surface representation, the surface
--            entity bounded and a collection of boundary entities

        theType       : Integer;
        theSurface    : IGESEntity;
        theBoundaries : HArray1OfBoundary;

end BoundedSurface;
