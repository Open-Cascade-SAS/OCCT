-- Created on: 1999-11-26
-- Created by: Andrey BETENEV
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0

class ProductConceptContext from StepBasic
inherits ApplicationContextElement from StepBasic

    ---Purpose: Representation of STEP entity ProductConceptContext

uses
    HAsciiString from TCollection,
    ApplicationContext from StepBasic

is
    Create returns ProductConceptContext from StepBasic;
	---Purpose: Empty constructor

    Init (me: mutable; aApplicationContextElement_Name: HAsciiString from TCollection;
                       aApplicationContextElement_FrameOfReference: ApplicationContext from StepBasic;
                       aMarketSegmentType: HAsciiString from TCollection);
	---Purpose: Initialize all fields (own and inherited)

    MarketSegmentType (me) returns HAsciiString from TCollection;
	---Purpose: Returns field MarketSegmentType
    SetMarketSegmentType (me: mutable; MarketSegmentType: HAsciiString from TCollection);
	---Purpose: Set field MarketSegmentType

fields
    theMarketSegmentType: HAsciiString from TCollection;

end ProductConceptContext;
