-- Created on: 1993-02-03
-- Created by: Gilles DEBARBOUILLE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class InstanceParameter from Dynamic

inherits

    Parameter from Dynamic

	---Purpose: This class describes a parameter with a dynamic 
	--          fuzzy instance as value.

uses

    CString from Standard,
    OStream from Standard,
    DynamicInstance from Dynamic


is

    Create(aparameter : CString from Standard)
    
    ---Level: Public 
    
    ---Purpose: Creates an   InstanceParameter  with  <aparameter>  as
    --          identifier.
    
    returns mutable InstanceParameter from Dynamic;
    
    Create(aparameter : CString from Standard; avalue : DynamicInstance from Dynamic) 

    ---Level: Public 
    
    ---Purpose: Creates   an  InstanceParameter  with  <aparameter>  as
    --          identifier and <avalue> as initial value.

    returns mutable InstanceParameter from Dynamic;
    
    Value(me) returns DynamicInstance from Dynamic
    
    ---Level: Public 
    
    ---Purpose: Returns <thevalue>.
    
    is static;
    
    Value(me : mutable ; avalue : DynamicInstance from Dynamic)
    
    ---Level: Public 
    
    ---Purpose: Sets <avalue> to <thevalue>.
    
    is static;

    Dump(me ; astream : in out OStream from Standard)
    
    ---Level: Public 
    
    ---Purpose: Useful for debugging.
    
    is redefined;
    
fields

    thevalue : DynamicInstance from Dynamic;

end InstanceParameter;
