-- Created on: 1999-02-11
-- Created by: Pavel DURANDIN
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Counter from STEPSelections

	---Purpose: 

uses
   
    Graph from Interface,
    MapOfTransient from TColStd,
    ConnectedFaceSet from StepShape,
    CompositeCurve from StepGeom
  
is
    Create returns Counter from STEPSelections;
    
    Count(me: in out;graph: Graph from Interface;
    	            start: Transient);
	  
    Clear(me: in out);
    
    NbInstancesOfFaces(me)  returns Integer;
    	---C++: inline
    	---Purpose:
    
    POP(me)  returns Integer;
    	---C++: inline
    	---Purpose:
    
    POP2(me)  returns Integer
    	---C++: inline
	;
    	---Purpose:
    
    NbInstancesOfShells(me) returns Integer;
    	---C++: inline
    	---Purpose:
    
    NbInstancesOfSolids(me) returns Integer;
    	---C++: inline
    	---Purpose:
    
    NbInstancesOfEdges(me) returns Integer;
    	---C++: inline
	---Purpose:
    
    NbInstancesOfWires(me) returns Integer;
    	---C++: inline
	---Purpose:
	
    NbSourceFaces(me)  returns Integer;
    	---C++: inline
    	---Purpose:
    
    NbSourceShells(me) returns Integer;
    	---C++: inline
    	---Purpose:
    
    NbSourceSolids(me) returns Integer;
    	---C++: inline
    	---Purpose:
	
    NbSourceEdges(me) returns Integer;
    	---C++: inline
	---Purpose:
	
    NbSourceWires(me) returns Integer;
    	---C++: inline
	---Purpose:
	
   AddShell(me: in out; cfs: ConnectedFaceSet from StepShape) is private;
   
   AddCompositeCurve(me: in out; ccurve: CompositeCurve from StepGeom) is private;

fields

    myNbFaces : Integer;
    myNbShells: Integer;
    myNbSolids: Integer;
    myNbEdges : Integer;
    myNbWires : Integer;
    
    myMapOfFaces : MapOfTransient from TColStd;
    myMapOfShells: MapOfTransient from TColStd;
    myMapOfSolids: MapOfTransient from TColStd;  
    myMapOfEdges : MapOfTransient from TColStd;
    myMapOfWires : MapOfTransient from TColStd;

end Counter;
