-- File:	BSplineCurve.cdl<2>
-- Created:	Fri May 22 09:53:01 1992
-- Author:	Jean Claude VAUTHIER
--		<jcv@sdsun4>
---Copyright:	 Matra Datavision 1992


class BSplineCurve


from DrawTrSurf


inherits Curve from DrawTrSurf


uses BSplineCurve from Geom,
     Color from Draw,
     MarkerShape from Draw,
     Display from Draw,
     Drawable3D from Draw


is


  Create (C : BSplineCurve from Geom)
        --- Purpose :
        --  creates a drawable BSpline curve from a BSpline curve of 
        --  package Geom.
     returns mutable BSplineCurve from DrawTrSurf;



  Create (C : BSplineCurve from Geom;
          CurvColor, PolesColor, KnotsColor : Color from Draw;
          KnotsShape : MarkerShape from Draw; KnotsSize : Integer;
          ShowPoles, ShowKnots : Boolean; Discret : Integer; Deflection : Real;
          DrawMode : Integer)
        --- Purpose :
        --  creates a drawable BSpline curve from a BSpline curve of 
        --  package Geom.
     returns mutable BSplineCurve from DrawTrSurf;


  DrawOn (me; dis : in out Display from Draw)
     is redefined static;


  DrawOn (me; dis : in out Display from Draw;
          ShowPoles, ShowKnots : Boolean);


  DrawOn (me; 
          dis : in out Display from Draw; 
          U1, U2 : Real; 
          Pindex : Integer;
          ShowPoles : Boolean = Standard_True;
          ShowKnots : Boolean = Standard_True);


  ShowPoles (me : mutable)
     is static;


  ShowKnots (me : mutable)
     is static;
     

  ClearPoles (me : mutable)
     is static;
     
  
  ClearKnots (me : mutable)
     is static;
     

  FindPole(me; X,Y : Real; D : Display from Draw; Prec : Real; 
           Index : in out Integer)
        --- Purpose :
        --  Returns in <Index> the index of the first pole  of the
        --  curve projected by the Display <D> at a distance lower
        --  than <Prec> from <X,Y>. If no pole  is found  index is
        --  set to 0, else index is always  greater than the input
        --  value of index.
  is static;
  

  FindKnot(me; X,Y : Real; D : Display from Draw; Prec : Real; 
           Index : in out Integer)
  is static;
  

  SetPolesColor (me : mutable; aColor : Color from Draw)
        ---C++: inline
     is static;
     

  SetKnotsColor (me : mutable; aColor : Color from Draw)
        ---C++: inline
     is static;
     

  SetKnotsShape (me : mutable; Shape : MarkerShape from Draw)
        ---C++: inline
     is static;
     

  KnotsShape (me)  returns MarkerShape from Draw
        ---C++: inline
     is static;
     
  
  KnotsColor (me)  returns Color from Draw
        ---C++: inline
     is static;
     
  
  PolesColor (me)  returns Color from Draw
        ---C++: inline
     is static;
    
  Copy(me) returns mutable Drawable3D from Draw
	---Purpose: For variable copy.
  is redefined;	
    
    
fields

  drawPoles  : Boolean;
  drawKnots  : Boolean;
  knotsForm  : MarkerShape from Draw;
  knotsLook  : Color from Draw;
  knotsDim   : Integer;
  polesLook  : Color from Draw;
 
end BSplineCurve;

