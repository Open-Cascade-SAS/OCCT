-- File:	 CurveTool.cdl
-- Created:	 Wed Aug 26 15:32:21 1992
-- Author:       Jean-Claude Vauthier
---Copyright:	 Matra Datavision 1992





deferred generic class CurveTool from GProp (Curve as any)   

    --- Purpose :
    --  This template defines the minimum of methods required
    --  to compute the global properties of a C1 parametric
    --  curve in 3d space with the algorithmes of package GProp.
    --  To compute the global properties of your curves, you 
    --  have to define your own "CurveTool" using this template.  
    --
    --  Curve must be a bounded curve of continuity C1 defined in 3d
    --  space.

uses Pnt from gp,
     Vec from gp

is


  FirstParameter (myclass; C : Curve)   returns Real;
        --- Purpose :
        --  Returns the parametric value of the start point of
        --  the curve.  The curve is oriented from the start point
        --  to the end point.


  LastParameter (myclass; C : Curve)   returns Real;
        --- Purpose :
        --  Returns the parametric value of the end point of
        --  the curve.  The curve is oriented from the start point
        --  to the end point.


  IntegrationOrder (myclass; C : Curve)    returns Integer;
        --- Purpose :
        --  Returns the number of Gauss points required to do
        --  the integration with a good accuracy using the
        --  Gauss method.  For a polynomial curve of degree n
        --  the maxima of accuracy is obtained with an order
        --  of integration equal to 2*n-1.


  Value (myclass; C : Curve; U : Real)  returns Pnt;
    	--- Purpose : Returns the point of parameter U on the loaded curve.


  D1 (myclass; C : Curve; U: Real; P: out Pnt; V1: out Vec);
    	--- Purpose : 
    	--  Returns the point of parameter U and the first derivative
    	--  at this point.


end CurveTool;
