-- Created on: 1994-04-21
-- Created by: Christian CAILLET
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SelectSignature  from IFSelect    inherits SelectExtract

    ---Purpose : A SelectSignature sorts the Entities on a Signature Matching.
    --           The signature to match is given at creation time. Also, the
    --           required match is given at creation time : exact (IsEqual) or
    --           contains (the Type's Name must contain the criterium Text)
    --           
    --           Remark that no more interpretation is done, it is an
    --           alpha-numeric signature : for instance, DynamicType is matched
    --           as such, super-types are not considered
    --           
    --           Also, numeric (integer) comparisons are supported : an item
    --           can be <val ou <=val or >val or >=val , val being an Integer
    --           
    --           A SelectSignature may also be created from a SignCounter,
    --           which then just gives its LastValue as SignatureValue

uses CString, AsciiString from TCollection, Transient,
     SequenceOfAsciiString from TColStd,    SequenceOfInteger     from TColStd,
     InterfaceModel, Graph, Signature, SignCounter

is

    Create (matcher : Signature;
    	signtext : CString;
    	exact : Boolean = Standard_True)
    	returns SelectSignature;
    ---Purpose : Creates a SelectSignature with its Signature and its Text to
    --           Match.
    --           <exact> if True requires exact match,
    --           if False requires <signtext> to be contained in the Signature
    --           of the entity (default is "exact")

    Create (matcher : Signature;
    	    signtext : AsciiString from TCollection;
    	    exact : Boolean = Standard_True)
    	returns SelectSignature;
    ---Purpose : As above with an AsciiString

    Create (matcher : SignCounter;
    	signtext : CString;
    	exact : Boolean = Standard_True)
    	returns SelectSignature;
    ---Purpose : Creates a SelectSignature with a Counter, more precisely a
    --           SelectSignature. Which is used here to just give a Signature
    --           Value (by SignOnly Mode)
    --           Matching is the default provided by the class Signature

    Signature (me) returns Signature;
    ---Purpose : Returns the used Signature, then it is possible to access it,
    --           modify it as required. Can be null, hence see Counter

    Counter   (me) returns SignCounter;
    ---Purpose : Returns the used SignCounter. Can be used as alternative for
    --           Signature

    SortInGraph (me; rank : Integer; ent : Transient; G : Graph)
    	returns Boolean  is redefined;
    ---Purpose : Returns True for an Entity (model->Value(num)) of which the
    --           signature matches the text given as creation time
    --           May also work with a Counter from the Graph

    Sort (me; rank : Integer; ent : Transient; model : InterfaceModel)
    	returns Boolean;
    ---Purpose : Not called, defined only to remove a deferred method here

    SignatureText (me) returns AsciiString from TCollection;
    ---Purpose : Returns Text used to Sort Entity on its Signature or SignCounter
    ---C++ : return const &

    IsExact (me) returns Boolean;
    ---Purpose : Returns True if match must be exact

    ExtractLabel (me) returns AsciiString from TCollection;
    ---Purpose : Returns a text defining the criterium.
    --           (it refers to the text and exact flag to be matched, and is
    --           qualified by the Name provided by the Signature)

fields

    thematcher  : Signature;
    thecounter  : SignCounter;
    thesigntext : AsciiString from TCollection;
    theexact    : Integer;
    thesignlist : SequenceOfAsciiString from TColStd;
    thesignmode : SequenceOfInteger     from TColStd;

end SelectSignature;
