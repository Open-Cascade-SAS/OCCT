-- File:	StepToGeom_MakeBoundedCurve2d.cdl
-- Created:	Wed Aug  4 11:06:25 1993
-- Author:	Martine LANGLOIS
---Copyright:	 Matra Datavision 1993

class MakeBoundedCurve2d from StepToGeom

    ---Purpose: This class implements the mapping between classes 
    --          BoundedCurve from  
    --          StepGeom which describes a BoundedCurve from 
    --          prostep and BoundedCurve from  Geom2d.
    --          As BoundedCurve is an abstract BoundedCurve this class 
    --          is an access to the sub-class required.
  
uses BoundedCurve from Geom2d,
     BoundedCurve from StepGeom
     
is 

    Convert ( myclass; SC : BoundedCurve from StepGeom;
                       CC : out BoundedCurve from Geom2d )
    returns Boolean from Standard;

end MakeBoundedCurve2d;
