-- Created on: 1996-07-24
-- Created by: Herve LOUESSARD
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



package LocalAnalysis  

    ---Purpose:
    -- This package gives tools to check the local continuity 
    -- between two  points situated  on two curves or two surfaces. 

uses

    Standard,
    StdFail,
    LProp,
    GeomAbs,
    Geom,
    Geom2d,
    GeomLProp,
    gp
    
is


--  enumeration used to describe the  status error 
   
enumeration  StatusErrorType   is  NullFirstDerivative, NullSecondDerivative, 
                                 TangentNotDefined,NormalNotDefined,
                                 CurvatureNotDefined         
end  StatusErrorType; 

     
    class SurfaceContinuity;
    ---Purpose:
    -- This  class  computes  and gives  tools to check  the  local
    -- continuity  between two points situated  on 2  surfaces
    
    
    class CurveContinuity; 
    ---Purpose:
    -- This  class  compute
    -- s  and gives  tools to check  the  local
    -- continuity  between two points situated  on 2  curves) 
    
    
    
   
    Dump( surfconti : SurfaceContinuity from LocalAnalysis;
          o: in out OStream);	
    ---Purpose:
    -- This fonction gives informations  about a  variable CurveContinuity
	  
    Dump( curvconti : CurveContinuity from LocalAnalysis;
          o: in out OStream);	
    ---Purpose:
    -- This fonction gives informations  about a variable SurfaceContinuity 
	  
    	  	  
end LocalAnalysis; 




















