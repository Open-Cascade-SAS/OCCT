-- Created on: 1996-12-05
-- Created by: Flore Lantheaume/Odile Olivier
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Chamf2dDimension from AIS inherits Relation from AIS

	---Purpose: A framework to define display of 2D chamfers.
    	-- A chamfer is displayed with arrows and text. The text
    	-- gives the length of the chamfer if it is a symmetrical
    	-- chamfer, or the angle if it is not.


uses

    PresentationManager3d from PrsMgr,
    Presentation          from Prs3d,
    Selection             from SelectMgr,
    Shape                 from TopoDS,
    Pnt                   from gp,
    Plane                 from Geom,
    Dir                   from gp,
    Projector             from Prs3d,
    Transformation        from Geom,
    ExtendedString        from TCollection,
    ArrowSide             from DsgPrs,
    KindOfDimension       from AIS 
    
is
    Create (aFShape     : Shape          from TopoDS;
            aPlane        : Plane        from Geom;
	    aVal        : Real           from Standard;
	    aText       : ExtendedString from TCollection)	    
	---Purpose: Constructs the display object for 2D chamfers.
    	-- This object is defined by the face aFShape, the
    	-- dimension aVal, the plane aPlane and the text aText.
        
    returns Chamf2dDimension from AIS;

    Create (aFShape     : Shape          from TopoDS;
            aPlane        : Plane        from Geom;
	    aVal        : Real           from Standard;
	    aText       : ExtendedString from TCollection;	    
	    aPosition   : Pnt            from gp;
	    aSymbolPrs  : ArrowSide      from DsgPrs;    
    	    anArrowSize : Real           from Standard = 0.0)
	---Purpose:  Constructs the display object for 2D chamfers.
    	-- This object is defined by the face aFShape, the plane
    	-- aPlane, the dimension aVal, the position aPosition,
    	-- the type of arrow aSymbolPrs with the size
    	-- anArrowSize, and the text aText.
    returns Chamf2dDimension from AIS;

    KindOfDimension(me) 
	---Purpose: Indicates that we are concerned with a 2d length.
	---C++: inline
    returns KindOfDimension from AIS 
    is redefined;
    
    IsMovable(me) returns Boolean from Standard 
	---Purpose: Returns true if the 2d chamfer dimension is movable.
	---C++: inline    
    is redefined;
    
    -- Methods from PresentableObject
    
    Compute(me            : mutable;
  	    aPresentationManager: PresentationManager3d from PrsMgr;
    	    aPresentation : Presentation from Prs3d;
    	    aMode         : Integer from Standard= 0) 
    is redefined static private;
    
    Compute(me:mutable;
    	        aProjector: Projector from Prs3d;
                aPresentation: Presentation from Prs3d)
    is redefined static private;     

    Compute(me            : mutable;
    	    aProjector    : Projector from Prs3d;
    	    aTrsf         : Transformation from Geom;
	    aPresentation : Presentation from Prs3d)
    is redefined;
	 ---Purpose: computes the presentation according to a point of view
	 --          given by <aProjector>. 
	 --          To be Used when the associated degenerated Presentations 
	 --          have been transformed by <aTrsf> which is not a Pure
	 --          Translation. The HLR Prs can't be deducted automatically
	 --          WARNING :<aTrsf> must be applied
	 --          to the object to display before computation  !!!

    ComputeSelection(me         : mutable;
    	    	     aSelection : Selection from SelectMgr;
    	    	     aMode      : Integer from Standard)
    is redefined private;
    
    
    
fields

    myPntAttach : Pnt     from gp;
    myDir       : Dir     from gp;

end Chamf2dDimension;
