-- Created on: 1998-07-30
-- Created by: Christian CAILLET
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ParamEditor  from IFSelect    inherits Editor  from IFSelect

    ---Purpose : A ParamEditor gives access for edition to a list of TypedValue
    --           (i.e. of Static too)
    --           Its definition is made of the TypedValue to edit themselves,
    --           and can add some constants, which can then be displayed but
    --           not changed (for instance, system name, processor version ...)
    --           
    --           I.E. it gives a way of editing or at least displaying
    --           parameters as global

uses CString, Transient, AsciiString, HAsciiString, HSequenceOfHAsciiString,
     InterfaceModel, EditForm, TypedValue

is

    Create (nbmax : Integer = 100; label : CString = "") returns ParamEditor;
    ---Purpose : Creates a ParamEditor, empty, with a maximum count of params
    --           (default is 100)
    --           And a label, by default it will be "Param Editor"

    AddValue (me : mutable; val : TypedValue; shortname : CString = "");
    ---Purpose : Adds a TypedValue
    --           By default, its short name equates its complete name, it can
    --           be explicited

    AddConstantText (me : mutable; val : CString;
    	    	     shortname : CString; completename : CString = "");
    ---Purpose : Adds a Constant Text, it will be Read Only
    --           By default, its long name equates its shortname


    Label (me) returns AsciiString;

    Recognize (me; form : EditForm) returns Boolean;

    StringValue (me; form : EditForm;  num : Integer)
    	returns HAsciiString from TCollection;

    Load (me; form : EditForm; ent : Transient; model : InterfaceModel)
    	returns Boolean;

    Apply (me; form : EditForm; ent : Transient; model : InterfaceModel)
    	returns Boolean;



    StaticEditor (myclass; list : HSequenceOfHAsciiString;
    	    	  label : CString = "") returns ParamEditor;
    ---Purpose : Returns a ParamEditor to work on the Static Parameters of
    --           which names are listed in <list>
    --           Null Handle if <list> is null or empty

fields

    thelabel : AsciiString;

end ParamEditor;
