-- Created on: 2001-09-10
-- Created by: Sergey KUUL
-- Copyright (c) 2001-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class MapContainer from Transfer inherits TShared from MMgt

	---Purpose: 

uses

    DataMapOfTransientTransient from TColStd

is

    Create returns mutable MapContainer from Transfer;
     
    SetMapObjects(me : mutable; theMapObjects : in out DataMapOfTransientTransient from TColStd);
    	---Purposes:Set map already translated geometry objects.
	
    GetMapObjects(me: mutable) returns DataMapOfTransientTransient from TColStd;
    	---Purposes:Get map already translated geometry objects.
    	---C++:return &
fields

  myMapObj           : DataMapOfTransientTransient from TColStd;
  
end MapContainer;
