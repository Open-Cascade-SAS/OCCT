-- Created on: 1995-05-23
-- Created by: Robert COUBLANC
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class SensitiveArc from Select2D 
inherits SensitiveEntity from Select2D

	---Purpose: sensitive Areas for an Arc Of Circle
	--          One gives Radius and center,and limits.
	--          or a geometric circle.

uses
    Ax2d from gp,
    EntityOwner from SelectBasics,
    ListOfBox2d from SelectBasics

is
    Create (OwnerId      : EntityOwner from SelectBasics;
    	    OriginAxis   : Ax2d from gp;
	    Angle        : Real from Standard;
	    Radius       : Real from Standard;
    	    MaxPoints    : Integer=9)
    returns mutable SensitiveArc ;
    	---Level: Public 
    	---Purpose: Constructs a 2D sensitive arc object defined by the
    	-- owner OwnerId, the axis of origin OriginAxis, the
    	-- angle Angle, the radius Radius, and the maximum
    	-- number of points MaxPoints.
    	--          
    	--               _.
    	--       \ angle /|
    	--        \_____/
    	--         \   /  direction
    	--          \ /
    	--	         *

    Areas (me:mutable ; aresul : in out ListOfBox2d from SelectBasics) is static;
    	---Level: Public 
    	---Purpose: returns the sensitive areas for a circle...    
    
    Matches (me  : mutable ;
             X,Y : Real from Standard;
             aTol: Real from Standard;
             DMin: out Real from Standard) 
    returns Boolean is static;     
    	---Purpose: returns true if the minimum distance DMin
    	--          between the postion x,y and the circle is less than aTol..

	     
    Matches (me  :mutable; 
             XMin,YMin,XMax,YMax : Real from Standard;
             aTol: Real from Standard) 
    returns Boolean
    is static;

fields

    myradius : Real;
    myax2d   : Ax2d from gp;
    myangle  : Real;
    mynbpt   : Integer;
end SensitiveArc;

