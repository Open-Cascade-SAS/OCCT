-- Created on: 2000-06-07
-- Created by: Galina KULIKOVA
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class FixSmallBezierCurves from ShapeUpgrade inherits FixSmallCurves from ShapeUpgrade

	---Purpose: 

uses

    --HArray1OfCurve from TColGeom,
    --HArray1OfCurve from TColGeom2d,
    --HSequenceOfReal from TColStd,
    Edge from TopoDS,
    Face from TopoDS,
    Curve from Geom,
    Curve from Geom2d,
    Status from ShapeExtend
is

    Create returns FixSmallBezierCurves from ShapeUpgrade;
    ---Purpose :
    
    Approx(me : mutable; Curve3d :  out Curve from Geom;
    	   	    	 Curve2d :  out Curve from Geom2d;
    	    	    	 Curve2dR : out Curve from Geom2d;
    	    	    	 First, Last : in out Real) returns Boolean is redefined;
    --Perform(me : mutable; theSegments3d :in out HArray1OfCurve from TColGeom;
    --	    	    	 theKnots3d : in out HSequenceOfReal from TColStd;
    --	    	    	 theSegments2d :in out HArray1OfCurve from TColGeom2d;
    --	    	    	 theKnots2d : in out HSequenceOfReal from TColStd) returns Boolean is redefined;
    ---Purpose :
    


end FixSmallBezierCurves;
