-- File:	StdSelect_BRepSelectionTool.cdl
-- Created:	Wed Mar  8 16:20:52 1995
-- Author:	Mister rmi
--		<rmi@photon>
--           	 
--           	 Fri Apr 10 98 : rob : Add Boolean for automatic
--           	                       Triangulation on faces...
--           	 
---Copyright:	 Matra Datavision 1995



class BRepSelectionTool from StdSelect 

	---Purpose: Tool to create specific selections (sets of primitives)
	--          for Shapes from Topology.
	--          These Selections may be used  in dynamic selection 
	--          Mechanism 
	--          Given a Shape and a mode of selection 
	--          (selection of vertices,
	--          edges,faces ...) , This Tool Computes corresponding sensitive primitives,
	--          puts them in an entity called Selection (see package SelectMgr) and returns it. 
	--          
	--          
	--          A Priority for the decomposed pickable objects can be given ;
    	--         by default There is A Preset Hierachy:
    	--             Vertex             priority : 5
    	--             Edge               priority : 4
    	--             Wire               priority : 3
    	--             Face               priority : 2
    	--             Shell,solid,shape  priority : 1
	--         the default priority in the following methods has no sense - it's only taken in account
    	--         when the user gives a value between 0 and 10. 
	--          IMPORTANT : This decomposition creates BRepEntityOwner instances (from StdSelect).
	--                      which are stored in the Sensitive Entities coming from The Decomposition.
	--                      
	--                      the result of picking in a ViewerSelector return EntityOwner from SelectMgr;
	--                      to know what kind of object was picked :
	--                      
	--   ENTITY_OWNER -> Selectable() gives the selectableobject which
        --                          was decomposed into pickable elements.
	--  Handle(StdSelect_BRepOwner)::DownCast(ENTITY_OWNER) -> Shape() 
	--                            gives the real picked shape (edge,vertex,shape...)
	--                     

uses
    Selection         from SelectMgr,
    Shape             from TopoDS,
    Face              from TopoDS,
    ShapeEnum         from TopAbs,
    SelectableObject  from SelectMgr,
    BRepOwner         from StdSelect,
    SensitiveEntity   from Select3D,
    ListOfSensitive   from Select3D
is
    
    Load(myclass;
    	 aSelection        : mutable Selection from SelectMgr;
    	 aShape            : Shape             from TopoDS;
	 aType             : ShapeEnum         from TopAbs;
     theDeflection : Real from Standard;
     theDeviationAngle : Real from Standard;
	 AutoTriangulation : Boolean from Standard = Standard_True;
    	 aPriority         : Integer =-1;
    	 NbPOnEdge         : Integer = 9;
    	 MaximalParameter  : Real from Standard = 500);
    	---Level: Public 
    	---Purpose: Decomposition of <aShape> into sensitive entities following
    	--         a mode of decomposition <aType>. These entities are stored in <aSelection>.
    	--         BrepOwners are created to store the identity of the picked shapes
    	--         during the selection process.
    	--         In those BRepOwners is also stored the original shape.
    	--         But One can't get the selectable object which was decomposed to give
    	--         the sensitive entities.
    	--        maximal parameter is used for infinite objects, to limit the sensitive Domain....
    	--         If AutoTriangulation = True, a Triangulation will be 
    	--         computed for faces which have no existing one.
    	--         if AutoTriangulation = False the old algorithm will be 
    	--         called to compute sensitive entities on faces.



    Load(myclass;
    	 aSelection : mutable Selection from SelectMgr;
    	 Origin     : SelectableObject  from SelectMgr;
    	 aShape     : Shape             from TopoDS;
	 aType      : ShapeEnum         from TopAbs;
	     theDeflection : Real from Standard;
	     theDeviationAngle : Real from Standard;
       	 AutoTriangulation : Boolean from Standard = Standard_True;
    	 aPriority  : Integer =-1;
    	 NbPOnEdge  : Integer = 9;
    	 MaximalParameter : Real from Standard = 500);
    	---Purpose:  Same  functionnalities  ; the  only
    	--        difference is that  the selectable object from which the
    	--        selection comes is stored in each Sensitive EntityOwner;


   -- Load(myclass;
    --	 aSelection : mutable Selection from SelectMgr;
    --	 Users      : SequenceOfAddress from SelectBasics;
    --	 aShape     : Shape             from TopoDS;
    -- aType      : ShapeEnum         from TopAbs;
    --   	 AutoTriangulation : Boolean from Standard = Standard_True;
    --	 aPriority  : Integer =-1;
    --	 NbPOnEdge  : Integer = 9;
    --	 MaximalParameter : Real from Standard = 500);
    	---Level: Public 
    	---Purpose:decomposition of <aShape> into sensitive entities following
    	--         a mode of decomposition <aType>. These entities are stored in <aSelection> 
    	--         The Major difference is that the known users are first inserted in the
    	--         BRepOwners. the original shape is the last user...
    	--         (see EntityOwner from SelectBasics and BrepOwner)...


    GetStandardPriority(myclass; 
    	    	    	aShap: Shape     from TopoDS;
    	    	    	aType: ShapeEnum from TopAbs)
    returns Integer from Standard;
    	---Purpose: Returns the standard priority of the shape aShap having the type aType.
    	-- This priority is passed to a StdSelect_BRepOwner object.
    	-- You can use the function Load to modify the
    	-- selection priority of an owner to make one entity
    	-- more selectable than another one.

    ComputeSensitive(myclass;
    	    	     aShape     : Shape     from TopoDS;
		     anOwner    : BRepOwner from StdSelect;
		     aSelection : mutable Selection from SelectMgr;
		     theDeflection : Real from Standard;
		     theDeviationAngle : Real from Standard;
    	    	     NbPOnEdge  : Integer;
    	    	     MaximalParameter : Real from Standard;
    		     AutoTriangulation : Boolean from Standard = Standard_True) ;
    	---Purpose: Computes the sensitive primitives corresponding to
    	-- the subshape aShape with the owner anOwner.
    	-- Stores them in the SelectMgr_Selection object, and returns this object.
    	-- The number NbPOnEdge is used to define edges and wires.
    	-- In the case of infinite objects, the value
    	-- MaximalParameter serves to limit computation time
    	-- by limiting the sensitive area. The default value is 500.
    	-- If AutoTriangulation is true, triangulation will be
    	-- computed for the faces which have none. If it is false,
    	-- sensitive entities on these faces will be calculated.

    GetEdgeSensitive(myclass;
    	    	     aShape     : Shape     from TopoDS;
		     anOwner    : BRepOwner from StdSelect;
		     aSelection : mutable Selection from SelectMgr;
		     theDeflection : Real from Standard;
		     theDeflectionAngle : Real from Standard;
    	    	     NbPOnEdge  : Integer;
    	    	     MaximalParameter : Real from Standard;
    	    	     aSensitive : in out SensitiveEntity from Select3D) 
    is private;
    	---Level: Internal
    	---Purpose:	


    GetSensitiveForFace(myclass;
    	    	        aFace             : Face from TopoDS;
			anOwner           : BRepOwner from StdSelect;
			OutList           : in out ListOfSensitive from Select3D;
			AutoTriangulation : Boolean from Standard = Standard_True;
			NbPOnEdge         : Integer = 9;
    	    	        MaxiParam         : Real from Standard =500;
    	    	        InteriorFlag      : Boolean from Standard = Standard_True)
    returns Boolean from Standard;
    	---Purpose:   appends   to <OutList>   the  3D
	--          sensitive entities  created  for  selection of <aFace>
	--         if<InteriorFlag> =  False  the face  will  be sensitive only on its boundary
    	    	    	    	


end BRepSelectionTool;




