-- File:	BRepFill_MultiLineTool.cdl
-- Created:	Mon Nov 14 15:01:41 1994
-- Author:	Bruno DUMORTIER
--		<dub@fuegox>
---Copyright:	 Matra Datavision 1994

private class MultiLineTool from BRepFill

    ---Purpose: private  class   used  to  instantiate the  continuous
    --          approximations routines.

uses
     Pnt           from gp,
     Pnt2d         from gp,
     Vec           from gp,
     Vec2d         from gp,
     Array1OfPnt   from TColgp,
     Array1OfPnt2d from TColgp,
     Array1OfVec   from TColgp,
     Array1OfVec2d from TColgp,
     MultiLine     from BRepFill

is
    
    FirstParameter(myclass; ML: MultiLine from BRepFill) 
    	---Purpose: returns the first parameter of the Line.
    returns Real from  Standard;


    LastParameter(myclass; ML: MultiLine from BRepFill) 
    	---Purpose: returns the last parameter of the Line.
    returns Real from Standard;


    NbP2d(myclass; ML: MultiLine from BRepFill) 
    	---Purpose: Returns the number of 2d points of a MLine
    returns Integer from Standard;


    NbP3d(myclass; ML: MultiLine from BRepFill) 
    	---Purpose: Returns the number of 3d points of a MLine.
    returns Integer from Standard;


    Value(myclass; ML   :     MultiLine   from BRepFill; 
    	    	   U    :     Real        from Standard; 
    	    	   tabPt: out Array1OfPnt from TColgp);
    	---Purpose: returns the 3d points of the multipoint <MPointIndex>
    	--          when only 3d points exist.


    Value(myclass; ML     :     MultiLine     from BRepFill; 
    	    	   U      :     Real          from Standard; 
                   tabPt2d: out Array1OfPnt2d from TColgp);
    	---Purpose: returns the 2d points of the multipoint <MPointIndex>
    	--          when only 2d points exist.


    Value(myclass; ML     :     MultiLine     from BRepFill;
    	    	   U      :     Real          from Standard; 
            	   tabPt  : out Array1OfPnt   from TColgp;
    	    	   tabPt2d: out Array1OfPnt2d from TColgp);
    	---Purpose: returns the 3d and 2d points of the multipoint 
    	--          <MPointIndex>.


    D1(myclass; ML  :     MultiLine   from BRepFill;
    	    	U   :     Real        from Standard; 
    	    	tabV: out Array1OfVec from TColgp)
    returns Boolean from Standard;
    	---Purpose: returns the 3d derivative values of the multipoint 
    	--          <MPointIndex> when only 3d points exist.
    	--          returns False if the derivative cannot be computed.


    D1(myclass; ML    :     MultiLine     from BRepFill; 
    	        U     :     Real          from Standard; 
    	        tabV2d: out Array1OfVec2d from TColgp)
    returns Boolean from Standard;
    	---Purpose: returns the 2d derivative values of the multipoint 
    	--          <MPointIndex> only when 2d points exist.
    	--          returns False if the derivative cannot be computed.


    D1(myclass; ML    :     MultiLine     from BRepFill; 
    	    	U     :     Real          from Standard; 
             	tabV  : out Array1OfVec   from TColgp; 
    	    	tabV2d: out Array1OfVec2d from TColgp)
    returns Boolean from Standard;
    	---Purpose: returns the 3d and 2d derivative values of the 
    	--          multipoint <MPointIndex>.
    	--          returns False if the derivative cannot be computed.

end MultiLineTool;    
    
