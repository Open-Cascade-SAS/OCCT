-- Created on: 1996-09-23
-- Created by: Philippe MANGIN
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Modified:	Fri Jul 10 11:23:35 1998
--              JCT : Add WithRatio,MinM


class CompCurveToBSplineCurve from GeomConvert 

	---Purpose: Concat several curve in an BSplineCurve

uses
 ParameterisationType from Convert,
 BoundedCurve from Geom,
 BSplineCurve from Geom

--raises

is

    Create (BasisCurve : BoundedCurve from Geom; 
     	    Parameterisation : ParameterisationType from Convert 
    	    	       =  Convert_TgtThetaOver2)
	 ---Purpose: Initialize the algorithme with one curve
	 --        - Parameterisation is used to convert 
    returns CompCurveToBSplineCurve;
    
    Add (me : in out; 
         NewCurve   :  BoundedCurve from Geom;
         Tolerance  :  Real from Standard;
         After      :  Boolean from Standard = Standard_False; 
         WithRatio  :  Boolean from Standard = Standard_True; 
         MinM       :  Integer  from  Standard  =  0)
	---Purpose: Append a curve in  the BSpline Return False if the
	--          curve is not G0  with the BSplineCurve.  Tolerance
	--             is   used to   check   continuity  and decrease
	--          Multiplicity at the common Knot until MinM
	--          if MinM = 0, the common Knot can be removed
    returns Boolean;
       
    
    Add (me : in out; 
         FirstCurve : in out BSplineCurve from Geom;
    	 SecondCurve: in out BSplineCurve from Geom;
         After      : Boolean from Standard; 
         WithRatio  : Boolean from Standard; 
         MinM       : Integer from Standard)
	---Purpose: Concat two BSplineCurves.
    	is private;    
    
    BSplineCurve(me) returns BSplineCurve from Geom;

fields
 myCurve :  BSplineCurve from Geom;
 myTol   :  Real;
 myType  :  ParameterisationType from Convert;

end CompCurveToBSplineCurve;
