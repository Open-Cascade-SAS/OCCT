-- Created on: 1994-03-03
-- Created by: Joelle CHAUVET
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Modified:	Mon Nov  3 10:24:07 1997
--		new class CurveConstraint
-- Modified:	Mon Jan 12 10:46:37 1998
--		new method Organize
-- Modified:	Mon Feb 23 09:28:33 1998
--		new methods SameNumber, ComputeACR, InsertACR
--		for sections with different number of elements
-- Modified:	Thu Apr 30 15:27:04 1998
--		methods Organize and SameNumber are dispatched in
--		new methods SearchOrigin and SameNumberByACR for open wires
--		and SameNumberByPolarMethod and ComputeOrigin for closed wires
-- Modified:	Tue Nov  3 10:41:06 1998
--		add classe CompatibleWires


package BRepFill


uses
    MMgt,
    TCollection,
    TColStd,
    GeomAbs,
    gp, 
    Bnd,
    TopLoc,
    TColgp,
    MAT,
    Geom2d,
    TColGeom2d,
    TopAbs,
    TopoDS,
    TopTools,
    Geom,
    TColGeom,
    Geom2dAdaptor,
    Approx,
    Bisector,
    BRep,
    BRepTools,
    BRepAlgo,
    BRepSweep,
    GeomFill,
    BRepMAT2d,
    StdFail, 
    GeomPlate, 
    Adaptor3d, 
    Law, 
    GeomLProp

is
    enumeration TransitionStyle 
    is Modified, Right, Round end; 
    
    enumeration TypeOfContact
    is NoContact, Contact, ContactOnBorder end;
    
--    private class FilledPair;
    	---Purpose: A pair of bound shapes with the result.

    
    class Generator;

    deferred class SectionLaw; 
    	class ShapeLaw; 
    	class NSections; 
          
    class  Draft;
     
    deferred  class LocationLaw;  
    	class DraftLaw;
   	class Edge3DLaw; 
	class EdgeOnSurfLaw;
   	class ACRLaw; 

    class Pipe;

    class PipeShell; 

    class Evolved;

    class Sweep; 

    class CompatibleWires;

    class OffsetWire;

    class OffsetAncestors;


    class ListOfOffsetWire instantiates 
    	List from TCollection (OffsetWire from BRepFill);
    private class ApproxSeewing;

    imported MultiLine;
    
    private class ComputeCLine instantiates 
    	ComputeCLine from Approx (MultiLine);
	

    private class TrimSurfaceTool;

    private class TrimEdgeTool;

    private class  SectionPlacement;  
     
    private class  Section;  

    --class  TrimCorner;

--modified by NIZHNY-MKK  Tue Oct 21 17:43:15 2003
    class TrimShellCorner;
			     
    private  class  SequenceOfSection  instantiates   
    	Sequence  from TCollection (Section); 
	
    class DataMapOfNodeDataMapOfShapeShape instantiates 
    	DataMap from TCollection (Node                from MAT,
    	    	    	    	  DataMapOfShapeShape from TopTools,
    	    	    	    	  MapTransientHasher  from TColStd );
   
    class DataMapOfNodeShape instantiates 
    	DataMap from TCollection (Node                from MAT,
    	    	    	    	  Shape               from TopoDS,
   	    	    	    	  MapTransientHasher  from TColStd );
				  
    class DataMapOfShapeDataMapOfShapeListOfShape instantiates
    	DataMap from TCollection (Shape                      from TopoDS,
    	    	    	    	  DataMapOfShapeListOfShape  from TopTools,
    	    	    	    	  ShapeMapHasher             from TopTools ); 
				  
    class DataMapOfShapeSequenceOfReal	instantiates
        	DataMap from TCollection (Shape          from TopoDS,
    	    	    	    	          SequenceOfReal from TColStd,
    	    	    	    	          ShapeMapHasher from TopTools );

    class DataMapOfShapeSequenceOfPnt	instantiates
        	DataMap from TCollection (Shape          from TopoDS,
    	    	    	    	          SequenceOfPnt  from TColgp,
    	    	    	    	          ShapeMapHasher from TopTools ); 

    class DataMapOfOrientedShapeListOfShape instantiates
	    DataMap from TCollection (Shape                  from TopoDS,
		    	    	      ListOfShape            from TopTools,  
    	    	    	    	      OrientedShapeMapHasher from TopTools); 

    class IndexedDataMapOfOrientedShapeListOfShape instantiates
	    IndexedDataMap from TCollection (Shape                  from TopoDS,
		    	    	      	     ListOfShape            from TopTools,  
    	    	    	    	      	     OrientedShapeMapHasher from TopTools); 

    class DataMapOfShapeHArray2OfShape	instantiates
        	DataMap from TCollection (Shape          from TopoDS,
    	    	    	    	          HArray2OfShape from TopTools,
    	    	    	    	          ShapeMapHasher from TopTools); 


    class CurveConstraint ;

    class Filling; 

    private class FaceAndOrder;
    
    private class EdgeFaceAndOrder;
    
    private class SequenceOfFaceAndOrder instantiates
    	Sequence from TCollection (FaceAndOrder from BRepFill);
    
    private class SequenceOfEdgeFaceAndOrder instantiates
    	Sequence from TCollection (EdgeFaceAndOrder from BRepFill);
				      
    Face( Edge1 : Edge from TopoDS;
    	  Edge2 : Edge from TopoDS )
	  ---Purpose: Computes a ruled surface between two edges.
    returns Face from TopoDS;

    Shell( Wire1 : Wire from TopoDS;
    	   Wire2 : Wire from TopoDS )
	   ---Purpose: Computes a ruled surface between two wires.
	   --          The wires must have the same number of edges.
    returns Shell from TopoDS;    
    
    Axe (Spine       :        Shape   from TopoDS; 
    	 Profile     :        Wire    from TopoDS; 
    	 AxeProf     : in out Ax3     from  gp;
    	 ProfOnSpine : in out Boolean from Standard;
    	 Tol         :        Real    from Standard);
	   ---Purpose: Computes  <AxeProf>  as Follow. <Location> is 
	   --          the Position of the nearest vertex V  of <Profile>
	   --          to <Spine>.<XDirection> is confused with the tangent
	   --          to <Spine> at the projected point of V on the Spine.
	   --          <Direction> is normal to <Spine>.
	   --          <Spine> is a plane wire or a plane face.

	   --          <ProfOnSpine> is <False> if the distance
	   --          between <Profile> and <Spine> is high to <Tol>.
    	   
      
    SearchOrigin( W : in out Wire from TopoDS; 
                  P : Pnt  from  gp; 
                  V : Vec  from  gp; 
    	    	  Tol  :  Real)  is  private;
	   ---Purpose: Computes origins and orientation on a closed wire
          
    	   
    ComputeACR( wire : Wire from TopoDS; 
    	    	ACR  : out  Array1OfReal from TColStd );
	   ---Purpose:  Compute ACR on a  wire
    	   
    InsertACR( wire     : Wire from TopoDS; 
    	       ACRcuts  : Array1OfReal from TColStd; 
    	       prec     : Real  from  Standard )
	   ---Purpose:  Insert ACR on a  wire
    returns Wire from TopoDS;    	   
    	   

end BRepFill;







