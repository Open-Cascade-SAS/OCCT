-- Created on: 1991-04-03
-- Created by: Remi GILET
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Pnt2dBisec

from GccAna

	---Purpose: This class implements the algorithms used to 
	--          create the bisecting line between two 2d points 
    	-- Describes functions for building a bisecting line between two 2D points.
    	-- The bisecting line between two points is the bisector of
    	-- the segment which joins the two points, if these are not coincident.
    	-- The algorithm does not find a solution if the two points are coincident.
    	-- A Pnt2dBisec object provides a framework for:
    	-- -   defining the construction of the bisecting line,
    	-- -   implementing the construction algorithm, and consulting the result.

uses Pnt2d           from gp,
     Lin2d           from gp

raises NotDone       from StdFail

is

Create(Point1    : Pnt2d from gp ;
       Point2    : Pnt2d from gp ) returns Pnt2dBisec;

    	---Purpose: Constructs a bisecting line between the points Point1 and Point2.

IsDone(me) returns Boolean from Standard
is static;
    	---Purpose: Returns true (this construction algorithm never fails).
        
HasSolution(me) returns Boolean from Standard
is static;
    	---Purpose: Returns true if this algorithm has a solution, i.e. if the
    	-- two points are not coincident.
        
ThisSolution(me) returns Lin2d from gp
raises NotDone
is static;
    	---Purpose : Returns a line, representing the solution computed by this algorithm.

fields

    WellDone : Boolean from Standard;
    -- True if the algorithm succeeded.

    HasSol : Boolean from Standard;
    -- True if there is a solution.

    linsol   : Lin2d from gp;
    ---Purpose : The solutions.

end Pnt2dBisec;


