-- Created on: 1997-01-03
-- Created by: Christian CAILLET
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class FreeFormEntity  from StepData    inherits TShared

    ---Purpose : A Free Form Entity allows to record any kind of STEP
    --           parameters, in any way of typing
    --           It is implemented with an array of fields
    --           A Complex entity can be defined, as a chain of FreeFormEntity
    --           (see Next and As)

uses CString, AsciiString from TCollection,
     HSequenceOfAsciiString from TColStd,
     Field from StepData, HArray1OfField from StepData

is

    Create returns FreeFormEntity;
    ---Purpose : Creates a FreeFormEntity, with no field, no type

    SetStepType (me : mutable; typenam : CString);
    ---Purpose : Sets the type of an entity
    --           For a complex one, the type of this member

    StepType (me) returns CString;
    ---Purpose : Returns the recorded StepType
    --           For a complex one, the type of this member

    SetNext (me : mutable; next : FreeFormEntity; last : Boolean = Standard_True);
    ---Purpose : Sets a next member, in order to define or complete a Complex
    --           entity
    --           If <last> is True (D), this next will be set as last of list
    --           Else, it is inserted just as next of <me>
    --           If <next> is Null, Next is cleared

    Next (me) returns FreeFormEntity;
    ---Purpose : Returns the next member of a Complex entity
    --           (remark : the last member has none)

    IsComplex (me) returns Boolean;
    ---Purpose : Returns True if a FreeFormEntity is Complex (i.e. has Next)

    Typed (me; typenam : CString) returns FreeFormEntity;
    ---Purpose : Returns the member of a FreeFormEntity of which the type name
    --           is given (exact match, no sub-type)

    TypeList (me) returns HSequenceOfAsciiString;
    ---Purpose : Returns the list of types (one type for a simple entity),
    --           as is (non reordered)

    Reorder (myclass; ent : in out FreeFormEntity) returns Boolean;
    ---Purpose : Reorders a Complex entity if required, i.e. if member types
    --           are not in alphabetic order
    --           Returns False if nothing done (order was OK or simple entity),
    --           True plus modified <ent> if <ent> has been reordered


    SetNbFields (me : mutable; nb : Integer);
    ---Purpose : Sets a count of Fields, from scratch

    NbFields (me) returns Integer;
    ---Purpose : Returns the count of fields

    Field (me; num : Integer) returns Field;
    ---Purpose : Returns a field from its rank, for read-only use
    ---C++ : return const &

    CField (me : mutable; num : Integer) returns Field;
    ---Purpose : Returns a field from its rank, in order to modify it
    ---C++ : return &

fields

    thetype   : AsciiString from TCollection;
    thefields : HArray1OfField;
    thenext   : FreeFormEntity;

end FreeFormEntity;
