-- Created on: 1995-12-08
-- Created by: Laurent BOURESCHE
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class CornerState from GeomFill 

	---Purpose: Class  (should    be  a  structure)   storing  the
	--          informations         about     continuity, normals
	--          parallelism,  coons conditions and bounds tangents
	--          angle on the corner of contour to be filled.

is

    Create returns CornerState from GeomFill;
    Gap(me) returns Real from Standard;
    Gap(me : in out; G : Real from Standard);
    TgtAng(me) returns Real from Standard;
    TgtAng(me : in out; Ang : Real from Standard);
    HasConstraint(me) returns Boolean from Standard;
    Constraint(me : in out);
    NorAng(me) returns Real from Standard;
    NorAng(me : in out; Ang : Real from Standard);
    IsToKill(me; Scal : out Real from Standard) 
    returns Boolean from Standard;
    DoKill(me : in out; Scal : Real from Standard);
    
fields

    gap           : Real from Standard;
    tgtang        : Real from Standard;
    isconstrained : Boolean from Standard;
    norang        : Real from Standard;
    scal          : Real from Standard;
    coonscnd      : Boolean from Standard;

end CornerState;
