-- Created on: 1993-01-11
-- Created by: CKY / Contract Toubro-Larsen ( TCD )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class NetworkSubfigure from IGESDraw  inherits IGESEntity

        ---Purpose : defines IGES Network Subfigure Instance Entity,
        --           Type <420> Form Number <0> in package IGESDraw
        --
        --           Used to specify each instance of Network Subfigure
        --           Definition Entity (Type 320, Form 0).

uses

        XYZ                   from gp,
        HAsciiString          from TCollection,
        NetworkSubfigureDef   from IGESDraw,
        TextDisplayTemplate   from IGESGraph,
        ConnectPoint          from IGESDraw,
        HArray1OfConnectPoint from IGESDraw

raises OutOfRange

is

        Create returns mutable NetworkSubfigure;

        -- specific for the entity

        Init (me               : mutable;
              aDefinition      : NetworkSubfigureDef;
              aTranslation     : XYZ;
              aScaleFactor     : XYZ;
              aTypeFlag        : Integer;
              aDesignator      : HAsciiString;
              aTemplate        : TextDisplayTemplate;
              allConnectPoints : HArray1OfConnectPoint);
        ---Purpose : This method is used to set the fields of the class
        --           NetworkSubfigure
        --       - aDefinition      : Network Subfigure Definition Entity
        --       - aTranslation     : Translation data relative to the model
        --                            space or the definition space
        --       - aScaleFactor     : Scale factors in the definition space
        --       - aTypeFlag        : Type flag
        --       - aDesignator      : Primary reference designator
        --       - aTemplate        : Primary reference designator Text
        --                            display Template Entity
        --       - allConnectPoints : Associated Connect Point Entities

        SubfigureDefinition (me) returns NetworkSubfigureDef;
        ---Purpose : returns Network Subfigure Definition Entity specified by this entity

        Translation (me) returns XYZ from gp;
        ---Purpose : returns Translation Data relative to either model space or to
        -- the definition space of a referring entity

        TransformedTranslation (me) returns XYZ from gp;
        ---Purpose : returns the Transformed Translation Data relative to either model
        -- space or to the definition space of a referring entity

        ScaleFactors (me) returns XYZ from gp;
        ---Purpose : returns Scale factor in definition space(x, y, z axes)

        TypeFlag (me) returns Integer;
        ---Purpose : returns Type Flag which implements the distinction between Logical
        -- design and Physical design data,and is required if both are present.
        --         Type Flag = 0 : Not specified (default)
        --                   = 1 : Logical
        --                   = 2 : Physical

        ReferenceDesignator (me) returns HAsciiString from TCollection;
        ---Purpose : returns the primary reference designator

        HasDesignatorTemplate (me) returns Boolean;
        ---Purpose : returns True if Text Display Template Entity is specified,
        -- else False

        DesignatorTemplate (me) returns TextDisplayTemplate;
        ---Purpose : returns primary reference designator Text Display Template Entity,
        -- or null. If null, no Text Display Template Entity specified

        NbConnectPoints (me) returns Integer;
        ---Purpose : returns the number of associated Connect Point Entities

        ConnectPoint (me; Index : Integer) returns ConnectPoint
        raises OutOfRange;
        ---Purpose : returns the Index'th  associated Connect point Entity
        -- raises exception if Index <= 0 or Index > NbConnectPoints()

fields

--
-- Class    : IGESDraw_NetworkSubfigure
--
-- Purpose  : Declaration of the variables specific to a NetworkSubfigure.
--
-- Reminder : A  Network Subfigure Instance Entity is defined by :
--                  - a Network Subfigure Definition
--                  - translation data relative to referring entity's
--                     model or definition space
--                  - the scale factors in x,y and z directions
--                  - a type flag to distinguish logical design data
--                     from physical data
--                     Type flag : 0 = not specified (default)
--                                 1 = logical
--                                 2 = physical
--                  - the pointers to associated Connect Point Entities
--

        theSubfigureDefinition   : NetworkSubfigureDef;

        theTranslation           : XYZ;

        theScaleFactor           : XYZ;

        theTypeFlag              : Integer;

        theDesignator            : HAsciiString;

        theDesignatorTemplate    : TextDisplayTemplate;

        theConnectPoints         : HArray1OfConnectPoint;

end NetworkSubfigure;
