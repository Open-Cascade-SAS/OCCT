-- Created on: 2002-11-13
-- Created by: Galina KULIKOVA
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class RemoveLocations from ShapeUpgrade inherits TShared from MMgt

	---Purpose: Removes all locations sub-shapes of specified shape

uses
    ShapeEnum from TopAbs,
    Shape from TopoDS,
    MapOfShape from TopTools,
    DataMapOfShapeShape from TopTools
is
    Create returns RemoveLocations from ShapeUpgrade;
    	---Purpose:Empy constructor
    
    Remove(me : mutable;theShape : Shape from TopoDS) returns Boolean;
    	---Purpose:Removes all location correspodingly to RemoveLevel.
    
    MakeNewShape(me : mutable;theShape , theAncShape: Shape from TopoDS; 
    	    	 theNewShape:in out Shape from TopoDS;theRemoveLoc : Boolean) 
    	    	     returns Boolean is private;
    
    GetResult(me) returns Shape from TopoDS;
    	---Purpose:Returns shape with removed locatins.
    	---C++: inline
	
    SetRemoveLevel(me: mutable; theLevel : ShapeEnum from TopAbs);
    	---Purpose:sets level starting with that location will be removed, 
    	--         by default TopAbs_SHAPE. In this case locations will be kept for specified shape
    	--         and if specified shape is TopAbs_COMPOUND for sub-shapes of first level.
    	---C++: inline
	
    RemoveLevel(me) returns ShapeEnum from TopAbs;
    	---Purpose:sets level starting with that location will be removed.Value of level can be set to
    	--         TopAbs_SHAPE,TopAbs_COMPOUND,TopAbs_SOLID,TopAbs_SHELL,TopAbs_FACE.By default TopAbs_SHAPE.
	--         In this case location will be removed for all shape types for exception of compound.
    	---C++: inline
    
	
    ModifiedShape (me; theInitShape : Shape from TopoDS) returns Shape from TopoDS;
    	---Purpose: Returns modified shape obtained from initial shape. 
	---C++: inline
    
fields
    myLevelRemoving : ShapeEnum from TopAbs;
    myShape : Shape from TopoDS;
    myMapNewShapes : DataMapOfShapeShape from TopTools;
    
end RemoveLocations;
