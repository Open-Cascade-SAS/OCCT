-- Created on: 1993-12-03
-- Created by: Christophe MARION
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


package BRepExtrema

    ---Purpose: This package gives   tools to compute  extrema between
    --          Shapes from BRep.

uses 
    Standard,
    StdFail,
    TopoDS,
    GeomAdaptor,
    BRepAdaptor,
    gp,
    Extrema,
    TColStd,
    TopTools,
    TCollection,
    Bnd
    
is

    ----------------------------------------------------------
    --  Extrema between two Shapes with triangulation.
    ----------------------------------------------------------
    imported Poly;


    ----------------------------------------------------------
    --  Extrema between a Point and an Edge.
    ----------------------------------------------------------
    imported ExtPC;


    ----------------------------------------------------------
    --  Extrema between two Edges.
    ----------------------------------------------------------
    imported ExtCC;


    ----------------------------------------------------------
    --  Extrema between a Point and a Face.
    ----------------------------------------------------------
    imported ExtPF;


    ----------------------------------------------------------
    --  Extrema between an Edge  and a Face.
    ----------------------------------------------------------
    imported ExtCF;


    ----------------------------------------------------------
    --  Extrema between two Faces.
    ----------------------------------------------------------
    imported ExtFF;


    ----------------------------------------------------------
    --  
    ----------------------------------------------------------
    exception UnCompatibleShape inherits DomainError;


    ----------------------------------------------------------
    --  enumeration used to describe the type of the support solution:                                         
    -- 	    IsVertex => The solution is a vertex.
    -- 	    IsOnEdge => The solution belongs to an Edge.
    -- 	    IsInFace => The solution is inside a Face.    
     
    ----------------------------------------------------------
    imported SupportType;


    ----------------------------------------------------------
    -- This  class gives tools  to  compute the minimum distance value
    -- between two shapes and  the corresponding couples of solution points.  
    
    ----------------------------------------------------------
    imported DistShapeShape;


    ----------------------------------------------------------
    --  This class is used to store a solution on a Shape. 
    --  (used only by class DistShapeShape)
    ----------------------------------------------------------
    imported SolutionElem;


    ----------------------------------------------------------
    -- This sequence is used to store all the solution on each Shape.
    ----------------------------------------------------------
    imported SeqOfSolution;

    imported DistanceSS;

end BRepExtrema;
