-- Created on: 1997-05-13
-- Created by: Stagiaire Francois DUMONT
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DenominatorMultiplier from GeomLib

       ---Purpose: this defines an evaluator for a function of 2 variables
       --          that will be used by CancelDenominatorDerivative in one
       --          direction.

uses

    BSplineSurface    from Geom,
    Array1OfReal      from TColStd
   
raises

    OutOfRange from Standard,
    ConstructionError from Standard
is

    Create( Surface           : BSplineSurface from Geom ;
    	    KnotVector        : Array1OfReal   from TColStd)
    returns DenominatorMultiplier from GeomLib
    raises
        ConstructionError from Standard;
       
     ---Purpose: if the surface is rational this will define the evaluator
     --          of a real function of 2 variables a(u,v) such that
     --          if we define a new surface by :
     --                       a(u,v) * N(u,v) 
     --          NewF(u,v) = ----------------
     --                       a(u,v) * D(u,v) 
    
    
    Value(me; UParameter : in Real from Standard ;
    	      VParameter : in Real from Standard) 

    returns Real from Standard
    raises
    	OutOfRange from Standard
    	---Purpose: Returns the value of 
    	--          a(UParameter,VParameter)=
    	--          
    	--            H0(UParameter)/Denominator(Umin,Vparameter)
    	--            
    	--            D Denominator(Umin,Vparameter)
        --          - ------------------------------[H1(u)]/(Denominator(Umin,Vparameter)^2)
        --            D U
        --            
        --          + H3(UParameter)/Denominator(Umax,Vparameter)
        --          
        --            D Denominator(Umax,Vparameter)
        --          - ------------------------------[H2(u)]/(Denominator(Umax,Vparameter)^2)
        --            D U
    is static;

    
fields
    
    mySurface          : BSplineSurface  from Geom  ;
    myKnotFlatVector   : Array1OfReal from TColStd  ;              
    

end MakeCurvefromApprox;



