-- File:	BRepCheck_Analyzer.cdl
-- Created:	Fri Dec  8 15:57:56 1995
-- Author:	Jacques GOUSSARD
--		<jag@bravox>
---Copyright:	 Matra Datavision 1995


class Analyzer from BRepCheck

	---Purpose: A framework to check the overall
    	-- validity of a shape. For a shape to be valid in Open
    	--  CASCADE, it - or its component subshapes - must respect certain
    	-- criteria. These criteria are checked by the function IsValid.
    	-- Once you have determined whether a shape is valid or not, you can
    	-- diagnose its specific anomalies and correct them using the services of
    	-- the ShapeAnalysis, ShapeUpgrade, and ShapeFix packages.

uses Shape                from TopoDS,
     ShapeEnum            from TopAbs,
     Result               from BRepCheck,
     DataMapOfShapeResult from BRepCheck

raises NullObject from Standard,
       NoSuchObject from Standard

is

    Create(S: Shape from TopoDS; 
           GeomControls : Boolean from Standard =  Standard_True)
    	---Purpose: Constructs a shape validation object defined by the shape S.
    	--    <S> is the  shape  to control.  <GeomControls>  If
    	--          False   only topological informaions  are checked.
    	--          The geometricals controls are
    	--          For a Vertex :
    	--          BRepCheck_InvalidToleranceValue  NYI
    	--          For an Edge :
    	--          BRepCheck_InvalidCurveOnClosedSurface,
    	--          BRepCheck_InvalidCurveOnSurface,
    	--          BRepCheck_InvalidSameParameterFlag,
   	--          BRepCheck_InvalidToleranceValue  NYI
    	--          For a face :
    	--          BRepCheck_UnorientableShape,
    	--          BRepCheck_IntersectingWires,
   	--          BRepCheck_InvalidToleranceValue  NYI
    	--          For a wire :
    	--          BRepCheck_SelfIntersectingWire

	---C++: inline
    	returns Analyzer from BRepCheck
	raises NullObject from Standard;
    	


    Init(me: in out; S: Shape from TopoDS;
                     GeomControls : Boolean from Standard =  Standard_True)
    	---Purpose: <S> is the  shape  to control.  <GeomControls>  If
    	--          False   only topological informaions  are checked.
    	--          The geometricals controls are
    	--          For a Vertex :
    	--          BRepCheck_InvalidTolerance  NYI
    	--          For an Edge :
    	--          BRepCheck_InvalidCurveOnClosedSurface,
    	--          BRepCheck_InvalidCurveOnSurface,
    	--          BRepCheck_InvalidSameParameterFlag,
   	--          BRepCheck_InvalidTolerance  NYI
    	--          For a face :
    	--          BRepCheck_UnorientableShape,
    	--          BRepCheck_IntersectingWires,
   	--          BRepCheck_InvalidTolerance  NYI
    	--          For a wire :
    	--          BRepCheck_SelfIntersectingWire

	raises NullObject from Standard
    	is static;
    
    	

    IsValid(me; S: Shape from TopoDS)
	---Purpose: <S> is a  subshape of the  original shape. Returns
	--          <STandard_True> if no default has been detected on
	--          <S> and any of its subshape.
    	returns Boolean from Standard
	raises NoSuchObject from Standard
	is static;


    IsValid(me)
    	---Purpose:  Returns true if no defect is
    	-- detected on the shape S or any of its subshapes.
    	-- Returns true if the shape S is valid.
    	-- This function checks whether a given shape is valid by checking that:
    	-- -      the topology is correct
    	-- -      parameterization of edges in particular is correct. 
    	-- For the topology to be correct, the following conditions must be satisfied:
    	-- -      edges should have at least two vertices if they are not
    	--    degenerate edges. The vertices should be within the range of
    	--  the bounding edges at the tolerance specified in the vertex,
    	-- -      edges should share at least one face. The representation of
    	--  the edges should be within the tolerance criterion assigned to them.
    	-- -      wires defining a face should not self-intersect and should be closed,
    	-- - there should be one wire which contains all other wires inside a face,
    	-- -      wires should be correctly oriented with respect to each of the edges,
    	-- -      faces should be correctly oriented, in particular with
    	--    respect to adjacent faces if these faces define a solid,
    	-- -      shells defining a solid should be closed. There should
    	--    be one enclosing shell if the shape is a solid;
    	--    To check parameterization of edge, there are 2 approaches depending on
    	--    the edge?s contextual situation.
    	-- -      if the edge is either single, or it is in the context
    	--    of a wire or a compound, its parameterization is defined by
    	--    the parameterization of its 3D curve and is considered as    valid.
    	-- -      If the edge is in the context of a face, it should
    	--    have SameParameter and SameRange flags set to Standard_True. To
    	--    check these flags, you should call the function
    	--    BRep_Tool::SameParameter and BRep_Tool::SameRange for an
    	--    edge. If at least one of these flags is set to Standard_False,
    	--    the edge is considered as invalid without any additional check.
    	--    If the edge is contained by a face, and it has SameParameter and
    	--    SameRange flags set to Standard_True, IsValid checks
    	--    whether representation of the edge on face, in context of which the
    	--    edge is considered, has the same parameterization up to the
    	--    tolerance value coded on the edge. For a given parameter t on the edge
    	--    having C as a 3D curve and one PCurve P on a surface S (base
    	--    surface of the reference face), this checks that |C(t) - S(P(t))|
    	--    is less than or equal to tolerance, where tolerance is the tolerance
    	--    value coded on the edge.
  	---C++: inline
    	returns Boolean from Standard
	is static;



    Result(me; SubS: Shape from TopoDS)
    
	---C++: return const&
	---C++: inline
    	returns any Result from BRepCheck
	raises NoSuchObject from Standard
	is static;


    --- Private implementation method

    Put(me: in out; S: Shape from TopoDS; Gctrl: Boolean from Standard)
    
    	is static private;


    Perform(me: in out; S: Shape from TopoDS)
    
	is static private;
	
    
    ValidSub(me; S: Shape from TopoDS; SubType: ShapeEnum from TopAbs)
    
    	returns Boolean from Standard
        is static private;
	
    
fields

    myShape : Shape                from TopoDS;
    myMap   : DataMapOfShapeResult from BRepCheck;
    
end Analyzer;
