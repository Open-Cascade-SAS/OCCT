-- Created on: 1994-04-01
-- Created by: Modelistation
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class HVertex from BRepTopAdaptor 

	---Purpose: 


inherits HVertex from Adaptor3d

uses Pnt2d       from gp,
     Orientation from TopAbs,
     Vertex      from TopoDS,
     HCurve2d    from Adaptor2d,
     HCurve2d    from BRepAdaptor

is

    Create(Vtx: Vertex from TopoDS; Curve: HCurve2d from BRepAdaptor)

    	returns HVertex from BRepTopAdaptor;


    Vertex(me)
    
    	returns Vertex from TopoDS
	---C++: inline
	---C++: return const&
	is static;


    ChangeVertex(me: mutable)
    
    	returns Vertex from TopoDS
	---C++: inline
	---C++: return&
	is static;


    Value(me: mutable)
    
    	returns Pnt2d from gp
	is redefined;


    Parameter(me: mutable; C: HCurve2d from Adaptor2d)
    
    	returns Real from Standard
	is redefined;


    Resolution(me: mutable; C: HCurve2d from Adaptor2d)
    
	---Purpose: Parametric resolution (2d).

    	returns Real from Standard
	is redefined;


    Orientation(me: mutable)
    
    	returns Orientation from TopAbs
	is redefined;


    IsSame(me: mutable; Other: like me)
    
    	returns Boolean from Standard
	is redefined;


fields -- redefined from HVertex from Adaptor3d

    myVtx   : Vertex   from TopoDS;
    myCurve : HCurve2d from BRepAdaptor;

end HVertex;
