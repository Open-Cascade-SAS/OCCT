-- File:	StepAP214_AppliedSecurityClassificationAssignment.cdl
-- Created:	Wed Mar 10 16:04:54 1999
-- Author:	data exchange team
--		<det@androx.nnov.matra-dtv.fr>
---Copyright:	 Matra Datavision 1999


class AppliedSecurityClassificationAssignment from StepAP214 
inherits SecurityClassificationAssignment from StepBasic
	

uses
    	HArray1OfSecurityClassificationItem from StepAP214, 
	SecurityClassificationItem from StepAP214, 
	SecurityClassification from StepBasic


is
    	Create returns mutable AppliedSecurityClassificationAssignment;
	---Purpose: Returns a AppliedSecurityClassificationAssignment


	Init (me : mutable;
	      aAssignedSecurityClassification : mutable SecurityClassification from StepBasic) is redefined;

	Init (me : mutable;
	      aAssignedSecurityClassification : mutable SecurityClassification from StepBasic;
	      aItems : mutable HArray1OfSecurityClassificationItem from StepAP214) is virtual;

	-- Specific Methods for Field Data Access --

	SetItems(me : mutable; aItems : mutable HArray1OfSecurityClassificationItem from StepAP214);
	Items (me) returns mutable HArray1OfSecurityClassificationItem from StepAP214;
	ItemsValue (me; num : Integer) returns SecurityClassificationItem;
	---C++: return const &
	NbItems (me) returns Integer;
    

fields

    items :  HArray1OfSecurityClassificationItem from StepAP214;

end AppliedSecurityClassificationAssignment;
