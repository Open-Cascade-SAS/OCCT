-- File:	StepBasic_Contract.cdl
-- Created:	Fri Nov 26 16:26:37 1999 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0
-- Copyright:	Matra Datavision 1999

class Contract from StepBasic
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity Contract

uses
    HAsciiString from TCollection,
    ContractType from StepBasic

is
    Create returns Contract from StepBasic;
	---Purpose: Empty constructor

    Init (me: mutable; aName: HAsciiString from TCollection;
                       aPurpose: HAsciiString from TCollection;
                       aKind: ContractType from StepBasic);
	---Purpose: Initialize all fields (own and inherited)

    Name (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Name
    SetName (me: mutable; Name: HAsciiString from TCollection);
	---Purpose: Set field Name

    Purpose (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Purpose
    SetPurpose (me: mutable; Purpose: HAsciiString from TCollection);
	---Purpose: Set field Purpose

    Kind (me) returns ContractType from StepBasic;
	---Purpose: Returns field Kind
    SetKind (me: mutable; Kind: ContractType from StepBasic);
	---Purpose: Set field Kind

fields
    theName: HAsciiString from TCollection;
    thePurpose: HAsciiString from TCollection;
    theKind: ContractType from StepBasic;

end Contract;
