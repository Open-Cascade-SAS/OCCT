-- Created on: 1991-07-19
-- Created by: Isabelle GRIGNON
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

private class MyRootFunction from CPnts 

inherits FunctionWithDerivative from math

---Purpose: Implements a function for the Newton algorithm to find the
--          solution of Integral(F) = L
--          (compute Length  and Derivative of the curve for Newton)

uses
    MyGaussFunction from CPnts,
    RealFunction    from CPnts

is

    Create returns MyRootFunction from CPnts;
	---C++: inline

    Init(me : in out;
           F : RealFunction from CPnts;
           D : Address from Standard;
    	   Order : Integer);
	---Purpose: F  is a pointer on a  function  D is a client data
	--          Order is the order of integration to use
	--          

    Init(me : in out; X0,L : Real);
	---Purpose: We want to solve Integral(X0,X,F(X,D)) = L

    Init(me : in out; X0,L,Tol : Real);
	---Purpose: We want to solve Integral(X0,X,F(X,D)) = L 
	--  with given tolerance
   
   Value(me:in out; X : Real; F : out Real)
    ---Purpose: This is Integral(X0,X,F(X,D)) - L
   returns Boolean
   is static;

   Derivative(me :in out; X: Real; Df : out Real)
    ---Purpose: This is F(X,D)
   returns Boolean
   is static;

   Values(me:in out; X : Real; F, Df : out Real)
   returns Boolean
   is static;

fields
   myFunction : MyGaussFunction from CPnts;
   myX0       : Real;
   myL        : Real;
   myOrder    : Integer;
   myTol      : Real;  -- rbv's modification 
end MyRootFunction;
