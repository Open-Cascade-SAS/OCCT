-- Created on: 1997-04-01
-- Created by: Christian CAILLET
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class FieldListN  from StepData    inherits FieldList  from StepData

    ---Purpose : Describes a list of fields, in a general way
    --           This basic class is for a null size list
    --           Subclasses are for 1, N (fixed) or Dynamic sizes

uses Field from StepData, Array1OfField from StepData

raises OutOfRange

is

    Create (nb : Integer) returns FieldListN;
    ---Purpose : Creates a FieldListN of <nb> Fields

    NbFields (me) returns Integer  is redefined;
    ---Purpose : Returns the count of fields. Here, returns starting <nb>

    Field  (me; num : Integer) returns Field
    ---Purpose : Returns the field n0 <num> between 1 and NbFields (read only)
	raises OutOfRange
    --           Error if <num> out of range
    	is redefined;
    ---C++ : return const &

    CField (me : in out; num : Integer) returns Field
    ---Purpose : Returns the field n0 <num> between 1 and NbFields, in order to
    --           modify its content
	raises OutOfRange
    --           Error if <num> out of range
    	is redefined;
    ---C++ : return &

    Destroy (me: in out) is virtual;
    ---C++ : alias "Standard_EXPORT virtual ~StepData_FieldListN() { Destroy(); }"


fields

    thefields : Array1OfField;

end FieldListN;
