-- Created on: 1992-11-17
-- Created by: Christian CAILLET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DispGlobal  from IFSelect  inherits Dispatch

    ---Purpose : A DispGlobal gathers all the input Entities into only one
    --           global Packet

uses AsciiString from TCollection, Graph, SubPartsIterator

is

    Create returns mutable DispGlobal;
    ---Purpose : Creates a DispGlobal

    Label (me) returns AsciiString from TCollection;
    ---Purpose : Returns as Label, "One File for all Input"

    	--  --    Evaluation    --  --

    LimitedMax (me; nbent : Integer; max : out Integer) returns Boolean
    	is redefined;
    ---Purpose : Returns True : maximum equates 1

    PacketsCount (me; G : Graph; count : out Integer) returns Boolean
    	is redefined;
    ---Purpose : Returns True (count of packets is well known) and count is 1

    Packets (me; G : Graph; packs : in out SubPartsIterator);
    ---Purpose : Computes the list of produced Packets. It is made of only ONE
    --           Packet, which gets the RootResult from the Final Selection.
    --           Remark : the inherited exception raising is never activated.

end DispGlobal;
