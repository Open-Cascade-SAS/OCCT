-- Created on: 1991-04-11
-- Created by: Michel CHAUVAT
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

--              Jean-Claude Vauthier January 1992, September 1992



generic class CGProps  from GProp (Curve     as any;
    	    	    	    	   Tool      as any -- as CurveTool(Curve)
    	    	    	    	  )

inherits GProps from GProp

	--- Purpose  : 
	--  Computes the  global properties of bounded curves 
	--  in 3D space. The curve must have at least a continuity C1. 
	--  It can be a curve as defined in the template CurveTool from 
	--  package GProp. This template gives the minimum of methods 
	--  required to evaluate the global properties of a curve 3D with  
	--  the algorithmes of GProp.

uses  Pnt   from gp
       
is

    Create returns CGProps;
  
    Create (C : Curve; CLocation : Pnt)  returns CGProps;

    SetLocation(me : in out;CLocation : Pnt) ;

    Perform(me : in out; C : Curve);

end CGProps;


