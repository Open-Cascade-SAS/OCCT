-- Created on: 2001-12-28
-- Created by: Andrey BETENEV
-- Copyright (c) 2001-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1

class EdgeBasedWireframeModel from StepShape
inherits GeometricRepresentationItem from StepGeom

    ---Purpose: Representation of STEP entity EdgeBasedWireframeModel

uses
    HAsciiString from TCollection,
    HArray1OfConnectedEdgeSet from StepShape

is
    Create returns EdgeBasedWireframeModel from StepShape;
	---Purpose: Empty constructor

    Init (me: mutable; aRepresentationItem_Name: HAsciiString from TCollection;
                       aEbwmBoundary: HArray1OfConnectedEdgeSet from StepShape);
	---Purpose: Initialize all fields (own and inherited)

    EbwmBoundary (me) returns HArray1OfConnectedEdgeSet from StepShape;
	---Purpose: Returns field EbwmBoundary
    SetEbwmBoundary (me: mutable; EbwmBoundary: HArray1OfConnectedEdgeSet from StepShape);
	---Purpose: Set field EbwmBoundary

fields
    theEbwmBoundary: HArray1OfConnectedEdgeSet from StepShape;

end EdgeBasedWireframeModel;
