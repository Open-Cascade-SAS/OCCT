-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ReparametrisedCompositeCurveSegment from StepGeom 

inherits CompositeCurveSegment from StepGeom 

uses

	Real from Standard, 
	TransitionCode from StepGeom, 
	Boolean from Standard, 
	Curve from StepGeom
is

	Create returns ReparametrisedCompositeCurveSegment;
	---Purpose: Returns a ReparametrisedCompositeCurveSegment


	Init (me : mutable;
	      aTransition : TransitionCode from StepGeom;
	      aSameSense : Boolean from Standard;
	      aParentCurve : Curve from StepGeom) is redefined;

	Init (me : mutable;
	      aTransition : TransitionCode from StepGeom;
	      aSameSense : Boolean from Standard;
	      aParentCurve : Curve from StepGeom;
	      aParamLength : Real from Standard) is virtual;

	-- Specific Methods for Field Data Access --

	SetParamLength(me : mutable; aParamLength : Real);
	ParamLength (me) returns Real;

fields

	paramLength : Real from Standard;

end ReparametrisedCompositeCurveSegment;
