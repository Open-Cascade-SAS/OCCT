-- File:	RWStepBasic_RWContractType.cdl
-- Created:	Fri Nov 26 16:26:38 1999 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0
-- Copyright:	Matra Datavision 1999

class RWContractType from RWStepBasic

    ---Purpose: Read & Write tool for ContractType

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    ContractType from StepBasic

is
    Create returns RWContractType from RWStepBasic;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : ContractType from StepBasic);
	---Purpose: Reads ContractType

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: ContractType from StepBasic);
	---Purpose: Writes ContractType

    Share (me; ent : ContractType from StepBasic;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWContractType;
