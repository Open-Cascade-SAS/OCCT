-- Created on: 1993-04-30
-- Created by: Yves FRICAUD
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class BasicElt from MAT 

	---Purpose: A    BasicELt  is  associated   to  each  elemtary
	--          constituant of  the figure.

inherits 

    TShared from MMgt

uses
    Arc            from MAT,
    Side           from MAT,
    Address        from Standard
is
    
    Create (anInteger : Integer) 
    	--- Purpose : Constructor, <anInteger> is the <index> of <me>.
    returns mutable BasicElt from MAT;

    StartArc(me)  
    	--- Purpose : Return <startArcLeft> or <startArcRight> corresponding
    	--            to <aSide>.
    returns Arc is static;

    EndArc(me)  
    	--- Purpose : Return <endArcLeft> or <endArcRight> corresponding
    	--            to <aSide>.
    returns Arc is static;
     
    Index (me) 
    	--- Purpose : Return the <index> of <me> in Graph.TheBasicElts.
    returns Integer is static;

    GeomIndex(me) 
    	--- Purpose : Return the <GeomIndex> of <me>.
    returns Integer is static;
    
    SetStartArc (me : mutable ; anArc : Arc)
    is static;
    
    SetEndArc (me : mutable ; anArc : Arc)
    is static;
    
    SetIndex (me : mutable ; anInteger : Integer)
    is static;

    SetGeomIndex(me : mutable ; anInteger : Integer)
    is static;
    
fields
    startLeftArc  : Address from Standard;
    endLeftArc    : Address from Standard;
    index         : Integer;
    geomIndex     : Integer;
    
end BasicElt;






