-- Created on: 2002-12-15
-- Created by: data exchange team
-- Copyright (c) 2002-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class ProductDefinitionFormationRelationship from StepBasic
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity ProductDefinitionFormationRelationship

uses
    HAsciiString from TCollection,
    ProductDefinitionFormation from StepBasic

is
    Create returns ProductDefinitionFormationRelationship from StepBasic;
	---Purpose: Empty constructor

    Init (me: mutable; aId: HAsciiString from TCollection;
                       aName: HAsciiString from TCollection;
                       aDescription: HAsciiString from TCollection;
                       aRelatingProductDefinitionFormation: ProductDefinitionFormation from StepBasic;
                       aRelatedProductDefinitionFormation: ProductDefinitionFormation from StepBasic);
	---Purpose: Initialize all fields (own and inherited)

    Id (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Id
    SetId (me: mutable; Id: HAsciiString from TCollection);
	---Purpose: Set field Id

    Name (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Name
    SetName (me: mutable; Name: HAsciiString from TCollection);
	---Purpose: Set field Name

    Description (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Description
    SetDescription (me: mutable; Description: HAsciiString from TCollection);
	---Purpose: Set field Description

    RelatingProductDefinitionFormation (me) returns ProductDefinitionFormation from StepBasic;
	---Purpose: Returns field RelatingProductDefinitionFormation
    SetRelatingProductDefinitionFormation (me: mutable; RelatingProductDefinitionFormation: ProductDefinitionFormation from StepBasic);
	---Purpose: Set field RelatingProductDefinitionFormation

    RelatedProductDefinitionFormation (me) returns ProductDefinitionFormation from StepBasic;
	---Purpose: Returns field RelatedProductDefinitionFormation
    SetRelatedProductDefinitionFormation (me: mutable; RelatedProductDefinitionFormation: ProductDefinitionFormation from StepBasic);
	---Purpose: Set field RelatedProductDefinitionFormation

fields
    theId: HAsciiString from TCollection;
    theName: HAsciiString from TCollection;
    theDescription: HAsciiString from TCollection;
    theRelatingProductDefinitionFormation: ProductDefinitionFormation from StepBasic;
    theRelatedProductDefinitionFormation: ProductDefinitionFormation from StepBasic;

end ProductDefinitionFormationRelationship;
