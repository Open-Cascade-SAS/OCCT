-- Created on: 1991-06-24
-- Created by: Christophe MARION
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- modified by jct (15/04/97)  add of  ModificationCommands




package GeomliteTest 

	---Purpose: this  package  provides  elementary commands for  curves  and
	--          surface.
uses
    Draw,
    Standard

is

    AllCommands(I : in out Interpretor from Draw);
	---Purpose: defines all geometric commands.
    
    CurveCommands(I : in out Interpretor from Draw);
	---Purpose: defines curve commands.
    
    SurfaceCommands(I : in out Interpretor from Draw);
	---Purpose: defines surface commands.
    
    API2dCommands(I : in out Interpretor from Draw);
	---Purpose: defines commands to test the Geom2dAPI
	--          - Intersection
	--          - Extrema
	--          - Projection
	--          - Approximation, interpolation 
    ApproxCommands(I : in out Interpretor from Draw);
	---Purpose: defines constrained curves commands.

    ModificationCommands(I : in out Interpretor from Draw);
	---Purpose: defines curves and surfaces modification commands.
	--          - Curve extension to point
	--          - Surface extension by length
    
    
end GeomliteTest;
