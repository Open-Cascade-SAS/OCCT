-- Created on: 1993-07-23
-- Created by: Jean Louis FRENKEL
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ColorPixel from Aspect inherits Pixel from Aspect

uses
    Color   from Quantity
is

    Create returns ColorPixel from Aspect;
	---Level: Public

    Create(aColor: Color from Quantity) returns ColorPixel from Aspect;
	---Level: Public

    Value (me) returns Color from Quantity is static ;
	---Level: Public
	   ---C++: return const &

    SetValue(me: in out; aColor: Color from Quantity) is static ;
	---Level: Public

    Print( me ; s : in out OStream from Standard ) is redefined static ;
	---Level: Public
	---Purpose : Prints the contents of <me> on the stream <s>

    HashCode (me; Upper : Integer ) returns Integer is redefined static ;
	---Level: Public
	---Purpose: Returns a hashed value denoting <me>. This value is in
	--         the range 1..<Upper>.
	---C++:  function call

    	IsEqual(me; Other : ColorPixel from Aspect) returns Boolean;
	    ---C++: alias operator==

    	IsNotEqual(me; Other : ColorPixel from Aspect) returns Boolean;
           ---C++: alias operator!=



fields
    myColor: Color from Quantity;

end ColorPixel from Aspect;
