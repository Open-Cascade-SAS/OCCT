-- Created on: 1991-02-22
-- Created by: Jean Claude Vauthier
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package GCPnts
        --- Purpose :
        --  This package  contains the geometric  algorithmes  used to
        --  compute characteristic points on parametrized curves.
        --  
        --  They are  high  level  algorithms based  on  the low level
        --  algorithms in CPnts.
    	---Level : Public. 
    	--  All methods of all  classes will be public.

uses Standard, TCollection, CPnts, Adaptor3d, Adaptor2d  , gp, GeomAbs,
     TColgp, StdFail, TColStd

is

   enumeration AbscissaType 
         is LengthParametrized, Parametrized, AbsComposite end;
	 
   enumeration DeflectionType 
         is Linear, Circular, Curved, DefComposite end;

   class AbscissaPoint;
   
   class UniformAbscissa;
   
   class UniformDeflection;

   class QuasiUniformDeflection;

   class QuasiUniformAbscissa;

   class TangentialDeflection;
   
end GCPnts;





