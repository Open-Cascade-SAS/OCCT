-- Created on: 1992-04-06
-- Created by: Christian CAILLET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class IGESType  from IGESData

    ---Purpose : taken from directory part of an entity (from file or model),
    --           gives "type" and "form" data, used to recognize entity's type

uses Integer

is

    Create returns IGESType;  -- default constructor (gives type = form = 0)

    Create (atype, aform : Integer) returns IGESType;

    Type (me) returns Integer  is static;
    ---Purpose : returns "type" data

    Form (me) returns Integer  is static;
    ---Purpose : returns "form" data

    IsEqual (me; another : IGESType) returns Boolean  is static;
    ---Purpose : compares two IGESTypes, avoiding comparing their fields
    ---C++ : alias operator ==

    Nullify (me : in out)  is static;
    ---Purpose : resets fields (usefull when an IGESType is stored as mask)

fields

    thetype : Integer;
    theform : Integer;

end IGESType;
