-- Created on: 1992-11-18
-- Created by: Remi LEQUETTE
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



package BRepClass 

	---Purpose: The  BRepClass packages provides    classification
	--          algorithms for the BRep topology.  It instantiates
	--          the algorithms from the package TopClass.

uses
    gp,
    TopAbs,
    TopoDS,
    TopExp,
    BRepTools,
    Geom2dInt,
    TopClass,
---    IntCurveSurface,
    Bnd




is
    class Edge;
	---Purpose: Stores the Edge and the Face.

    class Intersector;
	---Purpose: Intersect an Edge  with a segment.   This class is
	--          inherited   from   IntConicCurveOfGInter      from
	--          Geom2dInt.

    class FacePassiveClassifier instantiates Classifier2d from TopClass
    	(Edge         from BRepClass,
	 Intersector  from BRepClass);

    class FaceExplorer;
	---Purpose: Exploration of a Face to return UV edges.

    class FClassifier instantiates FaceClassifier from TopClass
    	(FaceExplorer from BRepClass,
	 Edge         from BRepClass,
	 Intersector  from BRepClass);
	 
    class FaceClassifier;
	---Purpose: Inherited    from   FClassifier   to   provide   a
	--          Constructor with a Face.

       
end BRepClass;
