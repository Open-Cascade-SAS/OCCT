-- Created on: 2002-12-12
-- Created by: data exchange team
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class FeaAxis2Placement3d from StepFEA
inherits Axis2Placement3d from StepGeom

    ---Purpose: Representation of STEP entity FeaAxis2Placement3d

uses
    HAsciiString from TCollection,
    CartesianPoint from StepGeom,
    Direction from StepGeom,
    CoordinateSystemType from StepFEA

is
    Create returns FeaAxis2Placement3d from StepFEA;
	---Purpose: Empty constructor

    Init (me: mutable; aRepresentationItem_Name: HAsciiString from TCollection;
                       aPlacement_Location: CartesianPoint from StepGeom;
                       hasAxis2Placement3d_Axis: Boolean;
                       aAxis2Placement3d_Axis: Direction from StepGeom;
                       hasAxis2Placement3d_RefDirection: Boolean;
                       aAxis2Placement3d_RefDirection: Direction from StepGeom;
                       aSystemType: CoordinateSystemType from StepFEA;
                       aDescription: HAsciiString from TCollection);
	---Purpose: Initialize all fields (own and inherited)

    SystemType (me) returns CoordinateSystemType from StepFEA;
	---Purpose: Returns field SystemType
    SetSystemType (me: mutable; SystemType: CoordinateSystemType from StepFEA);
	---Purpose: Set field SystemType

    Description (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Description
    SetDescription (me: mutable; Description: HAsciiString from TCollection);
	---Purpose: Set field Description

fields
    theSystemType: CoordinateSystemType from StepFEA;
    theDescription: HAsciiString from TCollection;

end FeaAxis2Placement3d;
