-- Created on: 1993-03-24
-- Created by: JCV
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Line from Geom2d inherits Curve from Geom2d

        --- Purpose : Describes an infinite line in the plane (2D space).
    	-- A line is defined and positioned in the plane with an
    	-- axis (gp_Ax2d object) which gives it an origin and a unit vector.
    	-- The Geom2d_Line line is parameterized as follows:
    	-- P (U) = O + U*Dir
    	-- where:
    	-- - P is the point of parameter U,
    	-- - O is the origin and Dir the unit vector of its positioning axis.
    	--   The parameter range is ] -infinite, +infinite [.
    	-- The orientation of the line is given by the unit vector
    	-- of its positioning axis.
    	-- See Also
    	-- GCE2d_MakeLine which provides functions for more
    	-- complex line constructions
    	-- gp_Ax2d
    	-- gp_Lin2d for an equivalent, non-parameterized data structure.
       

uses Ax2d     from gp,
     Dir2d    from gp, 
     Lin2d    from gp, 
     Pnt2d    from gp, 
     Vec2d    from gp,
     Trsf2d   from gp,
     Geometry from Geom2d,
     Shape    from GeomAbs


raises RangeError  from Standard

is

  Create (A : Ax2d)   returns mutable Line;
        --- Purpose :
        --  Creates a line located in 2D space with the axis placement A.
        --  The Location of A is the origin of the line. 


  Create (L : Lin2d)  returns mutable Line;
        --- Purpose :
        --  Creates a line by conversion of the gp_Lin2d line L.


  Create (P : Pnt2d; V : Dir2d)    returns mutable Line;
        --- Purpose : Constructs a line passing through point P and parallel to
    	--   vector V (P and V are, respectively, the origin
    	--   and the unit vector of the positioning axis of the line).


  SetLin2d (me : mutable; L : Lin2d);
        --- Purpose :
        --  Set <me> so that <me> has the same geometric properties as L.


  SetDirection (me : mutable; V : Dir2d);
        --- Purpose : changes the direction of the line.


  Direction (me) returns Dir2d from gp;
        --- Purpose : changes the direction of the line.
	---C++: return const &

  SetLocation (me : mutable; P : Pnt2d);
        --- Purpose : 
        --  Changes the "Location" point (origin) of the line.

  Location (me) returns Pnt2d from gp;
        --- Purpose : 
        --  Changes the "Location" point (origin) of the line.
	---C++: return const &

  SetPosition (me : mutable; A : Ax2d);
        --- Purpose :
        --  Changes the "Location" and a the "Direction" of <me>.

  Position(me) returns Ax2d from gp
	---C++: return const &
  is static;

  Lin2d (me)  returns Lin2d;
        --- Purpose : 
        --  Returns non persistent line from gp with the same geometric
        --  properties as <me>


  Reverse (me : mutable);
        --- Purpose : Changes the orientation of this line. As a result, the
    	-- unit vector of the positioning axis of this line is reversed.
      

  ReversedParameter(me; U : Real) returns Real;
	---Purpose: Computes the parameter on the reversed line for the
    	-- point of parameter U on this line.
    	-- For a line, the returned value is -U.


  FirstParameter (me)  returns Real;
        --- Purpose : Returns RealFirst  from  Standard.


  LastParameter (me)   returns Real;
        --- Purpose : Returns RealLast  from Standard


  IsClosed (me)  returns Boolean;
        --- Purpose : Returns False


  IsPeriodic (me)   returns Boolean;
        --- Purpose : Returns False


  Continuity (me)   returns Shape from GeomAbs;
        --- Purpose : Returns GeomAbs_CN, which is the global continuity of any line.

        
  Distance (me; P : Pnt2d)   returns Real;
        --- Purpose : Computes the distance between <me> and the point P.


  IsCN (me; N : Integer)   returns Boolean;
        --- Purpose : Returns True.

  D0(me; U : Real; P : out Pnt2d);
	---Purpose: Returns in P the point of parameter U.
       	--  P (U) = O + U * Dir where O is the "Location" point of the 
       	--  line and Dir the direction of the line.

  D1 (me; U : Real; P : out Pnt2d; V1 : out Vec2d);
        --- Purpose :
        --  Returns the point P of parameter u and the first derivative V1.


  D2 (me; U : Real; P : out Pnt2d; V1, V2 : out Vec2d);
        --- Purpose :
        --  Returns the point P of parameter U, the first and second 
        --  derivatives V1 and V2. V2 is a vector with null magnitude
        --  for a line.


  D3 (me; U : Real; P : out Pnt2d; V1, V2, V3 : out Vec2d);
        --- Purpose :
        --  V2 and V3 are vectors with null magnitude for a line.

        
  DN (me; U : Real; N : Integer)   returns Vec2d
        --- Purpose : For the point of parameter U of this line, computes
    	-- the vector corresponding to the Nth derivative.
    	-- Note: if N is greater than or equal to 2, the result is a
    	-- vector with null magnitude.
    	-- Exceptions Standard_RangeError if N is less than 1.
          raises RangeError;
    


  Transform (me : mutable; T : Trsf2d);
    	---Purpose: Applies the transformation T to this line.
    
    
  TransformedParameter(me; U : Real; T : Trsf2d from gp) returns Real
	---Purpose: Computes the parameter on the line transformed by
    	-- T for the point of parameter U on this line.
    	-- For a line, the returned value is equal to U multiplied
    	-- by the scale factor of transformation T.
     is redefined;  

  ParametricTransformation(me; T : Trsf2d from gp) returns Real
	---Purpose: Returns the coefficient required to compute the
    	-- parametric transformation of this line when
    	-- transformation T is applied. This coefficient is the
    	-- ratio between the parameter of a point on this line
    	-- and the parameter of the transformed point on the
    	-- new line transformed by T.
    	-- For a line, the returned value is the scale factor of the transformation T.
     is redefined;  




  Copy (me)  returns mutable like me;
    	---Purpose: Creates a new object, which is a copy of this line. 
    
fields

  pos : Ax2d;

end;
