-- Created on: 1994-12-16
-- Created by: Frederic MAUPAS
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Builder from StepToTopoDS
    inherits Root from StepToTopoDS
    
    ---Purpose:
    --         


uses

    ManifoldSolidBrep           from StepShape,
    BrepWithVoids               from StepShape,
    FacetedBrep                 from StepShape,
    FacetedBrepAndBrepWithVoids from StepShape,
    ShellBasedSurfaceModel      from StepShape,
    EdgeBasedWireframeModel     from StepShape,
    FaceBasedSurfaceModel       from StepShape,
    GeometricSet                from StepShape,
    Shape                       from TopoDS,
    BuilderError                from StepToTopoDS,
    TransientProcess            from Transfer,
    NMTool                      from StepToTopoDS
    
    raises NotDone from StdFail
     
is 

    Create returns Builder from StepToTopoDS;
    
    Create (S  : ManifoldSolidBrep from StepShape;
       	    TP : TransientProcess  from Transfer )
	returns Builder from StepToTopoDS;
     
    Create (S  : BrepWithVoids from StepShape;
            TP : TransientProcess  from Transfer )
    	returns Builder from StepToTopoDS;

    Create ( S : FacetedBrep from StepShape;
            TP : TransientProcess  from Transfer )
    	returns Builder from StepToTopoDS;

    Create (S  : FacetedBrepAndBrepWithVoids from StepShape;
            TP : TransientProcess  from Transfer )
    	returns Builder from StepToTopoDS;

    Create (S      : ShellBasedSurfaceModel from StepShape;
            TP     : TransientProcess  from Transfer;
            NMTool : in out NMTool from StepToTopoDS )
    	returns Builder from StepToTopoDS;

    Create ( S : GeometricSet from StepShape;
            TP : TransientProcess  from Transfer )
    	returns Builder from StepToTopoDS;

    Init (me : in out;
    	  S  : ManifoldSolidBrep from StepShape;
          TP : TransientProcess  from Transfer );

    Init (me : in out;
    	  S  : BrepWithVoids from StepShape;
          TP : TransientProcess  from Transfer );

    Init (me : in out;
    	  S  : FacetedBrep from StepShape;
          TP : TransientProcess  from Transfer );

    Init (me : in out;
    	  S  : FacetedBrepAndBrepWithVoids from StepShape;
          TP : TransientProcess  from Transfer );
	  
    Init (me     : in out;
    	   S     : ShellBasedSurfaceModel from StepShape;
          TP     : TransientProcess  from Transfer;
	  NMTool : in out NMTool from StepToTopoDS );
	  
    Init (me : in out;
    	  S  : EdgeBasedWireframeModel from StepShape;
          TP : TransientProcess  from Transfer );
	  
    Init (me : in out;
    	  S  : FaceBasedSurfaceModel from StepShape;
          TP : TransientProcess  from Transfer );
	  
    Init (me : in out;
    	  S  : GeometricSet from StepShape;
          TP : TransientProcess  from Transfer );
	  
    Value (me) returns Shape from TopoDS
    	raises NotDone
    	is static;
    	---C++: return const&
    
    Error (me) returns BuilderError from StepToTopoDS
    	is static;

fields

    myError  : BuilderError from StepToTopoDS;    
    
    myResult : Shape from TopoDS;
    
end Builder;
