-- Created on: 1993-06-11
-- Created by: Martine LANGLOIS
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MakeCartesianPoint from GeomToStep inherits Root from GeomToStep

    ---Purpose: This class implements the mapping between classes 
    --          CartesianPoint from Geom and Pnt from gp, and the class
    --          CartesianPoint from StepGeom which describes a point from
    --          Prostep. 
  
uses Pnt from gp,
     Pnt2d from gp,
     CartesianPoint from Geom,
     CartesianPoint from Geom2d,
     CartesianPoint from StepGeom
     
raises NotDone from StdFail
     
is 

Create ( P : Pnt from gp ) returns MakeCartesianPoint;

Create ( P : Pnt2d from gp ) returns MakeCartesianPoint;

Create ( P : CartesianPoint from Geom ) returns MakeCartesianPoint;

Create ( P : CartesianPoint from Geom2d ) returns MakeCartesianPoint;

Value (me) returns CartesianPoint from StepGeom
    raises NotDone
    is static;
    ---C++: return const&
    
fields

    theCartesianPoint : CartesianPoint from StepGeom;
    	-- The solution from StepGeom
    	
end MakeCartesianPoint;


