-- Created on: 1992-06-22
-- Created by: Gilles DEBARBOUILLE
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



deferred class FuzzyDefinitionsDictionary from Dynamic

inherits

    TShared from MMgt

	---Purpose: This  class groups   in  a dictionary  all  of the
	--          various definitions of  an object. It  also allows
	--          the  sharing of the   same definition by more than
	--          one  FuzzyInstance to  preserve a global coherence
	--          and also to manage  the memory.  To use this class
	--          an  inheritance  is  necessary with  perhaps   the
	--          overload  of  the  Switch  method if the parameter
	--          types   are   not  of  the  type BooleanParameter,
	--          IntegerParameter,        RealParameter         and
	--          StringParameter.
  
uses

    OStream from Standard,
    Integer from Standard,
    Boolean from Standard,
    CString from Standard,
    HAsciiString               from TCollection,
    Parameter                  from Dynamic,
    SequenceOfFuzzyDefinitions from Dynamic,
    FuzzyClass                 from Dynamic

is

    Initialize;
    
    ---Level: Internal 
    
    ---Purpose: Deferred constructor of the class.
    
    Creates(me : mutable ; afilename : CString from Standard)
    
    ---Level: Internal 
    
    ---Purpose: Starting with   a file named  <afilename>,  fills  the
    --          dictionary with all the wishes definitions.
    
    is static;
    
    Switch(me ; aname , atype , avalue : CString from Standard)
    
    ---Level: Internal 
    
    ---Purpose: This virtual method allows the user to add recognition
    --          of its  own  parameters when reading  the file to fill
    --          the dictionary.
    
    returns Parameter from Dynamic

    is virtual;
    
    Definition(me ; atype       : CString from Standard
                  ; adefinition : out FuzzyClass from Dynamic) returns Boolean from Standard
		  
    ---Level: Public 
    
    ---Purpose: Returns from     the dictionary in  the   out variable
    --          <adefinition> a reference to the right instance of the
    --          definition identified  by its type <atype>. The method
    --          returns true if the definition exist, false otherwise.
    
    is static;
    
    UpToDate(me) returns Boolean from Standard
    
    ---Level: Advanced 
    
    ---Purpose: Returns true if there has been  no modification of the
    --          file  fuzzyclasses.dat  since  the   creation  of  the
    --          dictionary object, false otherwise.
    
    is static;
    
    NumberOfDefinitions(me) returns Integer from Standard
    
    ---Level: Public 
    
    ---Purpose: Returns    the number  of  definitions  stored  in the
    --          dictionary.
    
    is static;
    
    Definition(me ; anindex : Integer from Standard) returns any FuzzyClass from Dynamic
    
    ---Level: Public 
    
    ---Purpose: Returns a  reference on the  definition identified  by
    --          the index <anidex>.
    
    is static;
    
    Dump(me ; astream : in out OStream from Standard)
    
    ---Level: Internal 
    
    ---Purpose: Useful for debugging.
    
    is static;

fields

    thefilename                   : HAsciiString               from TCollection;
    thetime                       : Integer from Standard                                ;
    thesequenceoffuzzydefinitions : SequenceOfFuzzyDefinitions from Dynamic    ;

end FuzzyDefinitionsDictionary;
