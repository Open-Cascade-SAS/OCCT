-- File:        FaceOuterBound.cdl
-- Created:     Mon Dec  4 12:02:26 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWFaceOuterBound from RWStepShape

	---Purpose : Read & Write Module for FaceOuterBound

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     FaceOuterBound from StepShape,
     EntityIterator from Interface

is

	Create returns RWFaceOuterBound;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable FaceOuterBound from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : FaceOuterBound from StepShape);

	Share(me; ent : FaceOuterBound from StepShape; iter : in out EntityIterator);

end RWFaceOuterBound;
