-- Created on: 1996-12-23
-- Created by: Alexander BRIVIN
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class SFRotation from Vrml 

	---Purpose: defines SFRotation type of VRML field types.
    	--          The  4  values  represent  an  axis  of  rotation  followed  by  amount  of 
	--          right-handed  rotation  about  the  that  axis, in  radians. 
is
 
    Create returns SFRotation from Vrml;

    Create ( aRotationX, aRotationY, aRotationZ : Real from Standard;
             anAngle : Real from Standard )   
    returns SFRotation from Vrml;

    SetRotationX ( me : in out; aRotationX : Real from Standard );
    RotationX ( me )  returns Real from Standard;

    SetRotationY ( me : in out; aRotationY : Real from Standard );
    RotationY ( me )  returns Real from Standard;

    SetRotationZ ( me : in out; aRotationZ : Real from Standard );
    RotationZ ( me )  returns Real from Standard;

    SetAngle ( me : in out; anAngle : Real from Standard );
    Angle ( me )  returns  Real from Standard;

fields

    myRotationX : Real from Standard;
    myRotationY : Real from Standard;
    myRotationZ : Real from Standard;
    myAngle     : Real from Standard;

end SFRotation;

