-- Created on: 1995-10-19
-- Created by: Andre LIEUTIER
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class D2 from Plate
---Purpose : define an order 2 derivatives of a 3d valued
--          function of a 2d variable
--         

uses XYZ from gp

is
    Create(duu,duv,dvv : XYZ from gp) returns D2;
    Create(ref  :  D2  from  Plate) returns D2;

fields
    
    Duu, Duv,Dvv : XYZ from gp;

friends
    class GtoCConstraint from Plate,
    class FreeGtoCConstraint from Plate    
end;
