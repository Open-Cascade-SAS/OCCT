-- Created on: 1993-01-22
-- Created by: Gilles DEBARBOUILLE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DynamicClass from Dynamic

inherits

    TShared from MMgt 
	---Purpose: A  dynamic class  is  defined   as a  sequence  of
	--          parameters and   as a   sequence of   methods. The
	--          specifications  are similar   to C++  classes. The
	--          class  has  to  be   defined  in terms  of  fields
	--          (Parameters) and methods. An instance of the class
	--          must be   made to set  the  fields and to  use the
	--          functionalities.

    
uses

    OStream from Standard,
    CString from Standard,
    HAsciiString      from TCollection,
    DynamicInstance   from Dynamic,
    Parameter         from Dynamic,
    ParameterNode     from Dynamic,
    Method            from Dynamic,
    SequenceOfMethods from Dynamic

    
is

    Create(aname : CString from Standard) returns mutable DynamicClass from Dynamic;
    
    ---Level: Public 
    
    ---Purpose: Creates a new empty instance of DynamicClass.
    
    Parameter(me : mutable ; aparameter : Parameter from Dynamic)
    
    ---Level: Public 
    
    ---Purpose: Adds another parameter <aparameter> to the sequence of
    --          parameter definitions.
    
    is static;
    
    CompiledMethod(me : mutable ; amethod , anaddress : CString from Standard)
    
    ---Level: Public 
    
    ---Purpose: Adds another method to the sequence of methods. It has
    --          <amethod> as name  and <anaddress> as mangled  name of
    --          the corresponding C++ function which must be called.
    
    is static;
    
    InterpretedMethod(me : mutable ; amethod , afile : CString from Standard)
    
    ---Level: Public 
    
    ---Purpose: Adds  another method to the  sequence of methods.   It
    --          has <amethod> as name and <afile> as interpreted file.
    
    is static;
    
    Method(me ; amethod : CString from Standard) returns any Method from Dynamic
    
    ---Level: Public 
    
    ---Purpose: Returns a reference to the method object identified by
    --          the string <amethod>.
    
    is virtual;
    
    Instance(me) returns mutable DynamicInstance from Dynamic
    
    ---Level: Public 
    
    ---Purpose: Returns an instance object of this class.

    is virtual;

    Dump(me ; astream : in out OStream from Standard)
    
    ---Level: Internal 
    
    ---Purpose: useful for debugging.

    is virtual;
    
fields

    thename               : HAsciiString      from TCollection;
    thefirstparameternode : ParameterNode     from Dynamic;
    thesequenceofmethods  : SequenceOfMethods from Dynamic;

end ;
