-- Created on: 1995-10-17
-- Created by: Andre LIEUTIER
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package Plate

uses
     TCollection,  TColStd,
     math, gp, TColgp
is

    class Plate; 
    
-- Basic  Constraints Class
    class PinpointConstraint;
    class LinearScalarConstraint;
    class LinearXYZConstraint;
--
-- geometric Constraints Class
--
    class GlobalTranslationConstraint;  
--    
    class PlaneConstraint; 
    class LineConstraint;  
--  
    class SampledCurveConstraint;
--   
--  class LinearizedHighlightConstraint;
--  
--  class DirectionalPressureConstraint;
--  
--  
--  Geometric contact of order k Constraint 
    class GtoCConstraint;
    class FreeGtoCConstraint;


-- utilities and internal Classes
    class D1;
    class D2;
    class D3;
    imported SequenceOfPinpointConstraint;
    imported SequenceOfLinearXYZConstraint;
    imported SequenceOfLinearScalarConstraint;
    imported Array1OfPinpointConstraint;    
    imported transient class HArray1OfPinpointConstraint;    
end Plate;
