-- Created on: 1992-11-17
-- Created by: Remi LEQUETTE
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package TopClass 

	---Purpose: The  package TopClass   provides    Classification
	--          algorithms.  A Classification algorithm is used to
	--          compute if  a  point is inside,  outside or on the
	--          boundary of a Shape.

uses
    gp,
    TopTrans, -- complex transitions
    TopAbs,   -- enumerations Orientation and State
    TopoDS,   
    IntRes2d,  -- to describe the result of intersections
    IntCurveSurface
---    TopExp   ------------- Pas Utilise mais sinon ca plante !!! 

is

    deferred generic class Intersection2d; 
	---Purpose: Describes   the  intersection algorithm     for 2d
	--          classifications. 
	
    generic class Classifier2d;
	---Purpose: Basic algorithm for 2d classifications.

    deferred generic class FaceExplorer;
	---Purpose: Defines  the   description  of   a  face  for  the
	--          FaceClassifier.

    generic class  FaceClassifier, FClass2d;
	---Purpose: Algorithm for classification in a Face.

	


    deferred class Intersection3d;
	---Purpose: Describes the intersection algorithm for 3d 
	--          classifications.    	    
		
    generic class Classifier3d;
    	---Purpose: Basic algorithm for 3d classification.
    	          
    deferred class SolidExplorer;
    	---Purpose: Defines the description of a solid for the 
    	--          SolidClassifier.
       
    generic class SolidClassifier;
    	---Purpose: Algorithm for classification in a Solid.
    
    
    
end TopClass;
