-- File:        Conic.cdl
-- Created:     Fri Dec  1 11:11:17 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class Conic from StepGeom 

inherits Curve from StepGeom 

uses

	Axis2Placement from StepGeom, 
	HAsciiString from TCollection
is

	Create returns mutable Conic;
	---Purpose: Returns a Conic


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aPosition : Axis2Placement from StepGeom) is virtual;

	-- Specific Methods for Field Data Access --

	SetPosition(me : mutable; aPosition : Axis2Placement);
	Position (me) returns Axis2Placement;

fields

	position : Axis2Placement from StepGeom; -- a SelectType

end Conic;
