-- File:	RWStepFEA_RWFeaShellMembraneBendingCouplingStiffness.cdl
-- Created:	Thu Dec 12 17:51:06 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWFeaShellMembraneBendingCouplingStiffness from RWStepFEA

    ---Purpose: Read & Write tool for FeaShellMembraneBendingCouplingStiffness

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    FeaShellMembraneBendingCouplingStiffness from StepFEA

is
    Create returns RWFeaShellMembraneBendingCouplingStiffness from RWStepFEA;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : FeaShellMembraneBendingCouplingStiffness from StepFEA);
	---Purpose: Reads FeaShellMembraneBendingCouplingStiffness

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: FeaShellMembraneBendingCouplingStiffness from StepFEA);
	---Purpose: Writes FeaShellMembraneBendingCouplingStiffness

    Share (me; ent : FeaShellMembraneBendingCouplingStiffness from StepFEA;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWFeaShellMembraneBendingCouplingStiffness;
