-- Created on: 2000-05-11
-- Created by: data exchange team
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1

class CharacterizedDefinition from StepRepr
inherits SelectType from StepData

    ---Purpose: Representation of STEP SELECT type CharacterizedDefinition

uses
    CharacterizedObject from StepBasic,
    ProductDefinition from StepBasic,
    ProductDefinitionRelationship from StepBasic,
    ProductDefinitionShape from StepRepr,
    ShapeAspect from StepRepr,
    ShapeAspectRelationship from StepRepr,
    DocumentFile from StepBasic

is
    Create returns CharacterizedDefinition from StepRepr;
	---Purpose: Empty constructor

    CaseNum (me; ent: Transient) returns Integer;
	---Purpose: Recognizes a kind of CharacterizedDefinition select type
	--          1 -> CharacterizedObject from StepBasic
	--          2 -> ProductDefinition from StepBasic
	--          3 -> ProductDefinitionRelationship from StepBasic
	--          4 -> ProductDefinitionShape from StepRepr
	--          5 -> ShapeAspect from StepRepr
	--          6 -> ShapeAspectRelationship from StepRepr
	--          7 -> DocumentFile from StepBasic
	--          0 else

    CharacterizedObject (me) returns CharacterizedObject from StepBasic;
	---Purpose: Returns Value as CharacterizedObject (or Null if another type)

    ProductDefinition (me) returns ProductDefinition from StepBasic;
	---Purpose: Returns Value as ProductDefinition (or Null if another type)

    ProductDefinitionRelationship (me) returns ProductDefinitionRelationship from StepBasic;
	---Purpose: Returns Value as ProductDefinitionRelationship (or Null if another type)

    ProductDefinitionShape (me) returns ProductDefinitionShape from StepRepr;
	---Purpose: Returns Value as ProductDefinitionShape (or Null if another type)
 
    ShapeAspect (me) returns ShapeAspect from StepRepr;
	---Purpose: Returns Value as ShapeAspect (or Null if another type)

    ShapeAspectRelationship (me) returns ShapeAspectRelationship from StepRepr;
	---Purpose: Returns Value as ShapeAspectRelationship (or Null if another type)

    DocumentFile (me) returns DocumentFile from StepBasic;
	---Purpose: Returns Value as DocumentFile (or Null if another type)

end CharacterizedDefinition;
