-- Created on: 2000-04-09
-- Created by: Sergey MOZOKHIN
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package STEPCAFControl

    ---Purpose : This package provides external access and control for STEP,
    --           on the level of CAF (shapes with attributes, external 
    --           references etc.)

uses 
    Dico,
    TCollection,
    TColStd,
    TopTools,
    TopoDS,
    IFSelect,
    Transfer,
    XSControl,
    STEPControl,
    STEPConstruct,
    StepShape,
    StepRepr,
    StepBasic,
    ShapeBuild,
    TDF,
    TDocStd,
    XCAFDoc,
    MoniTool

is

    class Reader;

    class Writer;

    class ExternFile;

    class ActorWrite;
    class Controller;

    class DictionaryOfExternFile instantiates 
    	  Dictionary from Dico (ExternFile from STEPCAFControl);

    imported DataMapOfShapeSDR;

    imported DataMapIteratorOfDataMapOfShapeSDR;

    --- skl
    imported DataMapOfShapePD;
    imported DataMapIteratorOfDataMapOfShapePD;

    imported DataMapOfSDRExternFile;

    imported DataMapIteratorOfDataMapOfSDRExternFile;

    --- skl
    imported DataMapOfPDExternFile;
    imported DataMapIteratorOfDataMapOfPDExternFile;

    imported DataMapOfLabelShape;

    imported DataMapIteratorOfDataMapOfLabelShape;

    imported DataMapOfLabelExternFile;

    imported DataMapIteratorOfDataMapOfLabelExternFile;

end STEPCAFControl;
