-- Created by: Peter KURNEV
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Tools from BOPDS 

	---Purpose: 
    	-- The class BOPDS_Tools contains  
    	-- a set auxiliary static functions  
	-- of the package BOPDS 

uses
    ShapeEnum from TopAbs 
  
--raises

is 
    TypeToInteger(myclass; 
    	    theT1: ShapeEnum from TopAbs; 
    	    theT2: ShapeEnum from TopAbs) 
    	returns Integer from Standard; 
    ---C++: inline  
     	---Purpose:  
     	--- Converts the conmbination of two types  
    	--  of shape <theT1>,<theT2>  
	--- to the one integer value, that is returned       
  
    TypeToInteger(myclass; 
    	    theT: ShapeEnum from TopAbs) 
    	returns Integer from Standard; 
    ---C++: inline  
     	---Purpose:  
     	--- Converts the type of shape <theT>,  
	--- to integer value, that is returned      	 
	
    HasBRep(myclass; 
    	    theT: ShapeEnum from TopAbs) 
    	returns Boolean from Standard;  
    ---C++: inline  
    	---Purpose:   
	--- Returns true if the type  <theT> correspond 
	--- to a shape having boundary representation 
  
    IsInterfering(myclass; 
    	    theT: ShapeEnum from TopAbs) 
	returns Boolean from Standard;   
    ---C++: inline 
    	---Purpose: 
        --- Returns true if the type <theT> can be participant of  
        --- an interference 	  

end Tools;
