-- Created on: 1994-06-10
-- Created by: Laurent PAINNOT
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



generic class WFRestrictedFace from Prs3d 
         (DrawFaceIso     as any;
    	  RestrictionTool as any)
	  
inherits Root from Prs3d
	 

	---Purpose: 

uses
    HSurface             from BRepAdaptor,
    Presentation         from Prs3d,
    Drawer               from Prs3d, 
    NListOfSequenceOfPnt from Prs3d,
    Length               from Quantity

--  Description of the isoparametric curves:
--  

is
    Add(myclass; aPresentation: Presentation from Prs3d; 
        	 aFace: HSurface from BRepAdaptor;
    	    	 aDrawer: Drawer from Prs3d);
		 
    AddUIso(myclass; aPresentation: Presentation from Prs3d; 
        	     aFace: HSurface from BRepAdaptor;
    	    	     aDrawer: Drawer from Prs3d);
		 
    AddVIso(myclass; aPresentation: Presentation from Prs3d; 
        	     aFace: HSurface from BRepAdaptor;
    	    	     aDrawer: Drawer from Prs3d);

    Add(myclass;  aPresentation: Presentation from Prs3d; 
    	          aFace: HSurface from BRepAdaptor;
		  DrawUIso, DrawVIso: Boolean from Standard;
		  Deflection: Length from Quantity;
		  NBUiso,NBViso: Integer from Standard;
		  aDrawer: Drawer from Prs3d; 
    	    	  Curves: out NListOfSequenceOfPnt from Prs3d);
		   
    Match(myclass; X,Y,Z: Length from Quantity;
                   aDistance: Length from Quantity;
        	   aFace: HSurface from BRepAdaptor;
    	    	   aDrawer: Drawer from Prs3d)
    returns Boolean from Standard;
		 
    MatchUIso(myclass; X,Y,Z: Length from Quantity;
                       aDistance: Length from Quantity;
        	       aFace: HSurface from BRepAdaptor;
    	    	       aDrawer: Drawer from Prs3d)
    returns Boolean from Standard;
		 
    MatchVIso(myclass; X,Y,Z: Length from Quantity;
                       aDistance: Length from Quantity;
         	       aFace: HSurface from BRepAdaptor;
    	    	       aDrawer: Drawer from Prs3d)
    returns Boolean from Standard;
		 
    Match(myclass;  X,Y,Z: Length from Quantity;
                  aDistance: Length from Quantity;
    	          aFace: HSurface from BRepAdaptor;
		  DrawUIso, DrawVIso: Boolean from Standard;
		  Deflection: Length from Quantity;
		  NBUiso,NBViso: Integer from Standard;
		  aDrawer: Drawer from Prs3d)

    returns Boolean from Standard;	  
		   
end WFRestrictedFace;

