-- File:        PlanarExtent.cdl
-- Created:     Mon Dec  4 12:02:28 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWPlanarExtent from RWStepVisual

	---Purpose : Read & Write Module for PlanarExtent

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     PlanarExtent from StepVisual

is

	Create returns RWPlanarExtent;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable PlanarExtent from StepVisual);

	WriteStep (me; SW : in out StepWriter; ent : PlanarExtent from StepVisual);

end RWPlanarExtent;
