-- Created on: 2007-05-29
-- Created by: Vlad Romashko
-- Copyright (c) 2007-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Tick from TDataStd inherits Attribute from TDF

    ---Purpose: Defines a boolean attribute.
    --          If it exists at a label - true,
    --          Otherwise - false.

uses 

    Attribute         from TDF,
    Label             from TDF,
    GUID              from Standard,
    Integer           from Standard,
    DataSet           from TDF,
    RelocationTable   from TDF

is

    ---Purpose: Static methods
    --          ==============

    GetID (myclass)   
    ---C++: return const &  
    returns GUID from Standard;


    Set (myclass; label : Label from TDF)  
    ---Purpose: Find, or create, a Tick attribute.
    returns Tick from TDataStd;  


    ---Purpose: Tick methods
    --          ============

    Create
    returns mutable Tick from TDataStd;


    ---Category: Inherited methods
    --           =================

    ID (me)
    ---C++: return const & 
    returns GUID from Standard;

    Restore (me: mutable; With : Attribute from TDF);

    NewEmpty (me)
    returns mutable Attribute from TDF;

    Paste (me; Into : mutable Attribute from TDF;
	       RT   : mutable RelocationTable from TDF);    

    Dump (me; anOS : in out OStream from Standard)
    returns OStream from Standard
    is redefined;
    ---C++: return &


end Tick;
