-- Created on: 1993-12-02
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

generic class Iterator from Blend (Item as any)

	---Purpose: Template class for an iterator.
	--          A Sequence from TCollection can implement this iterator.

is

    Create

	---Purpose: Creates an empty iterator.

    	returns Iterator;


    Clear(me: in out);

	---Purpose: Clears the content of the iterator.



    Append(me: in out; I: Item);

	---Purpose: Adds an element in the iterator.


    Length(me: in out)
    
	---Purpose: Returns the number of elements in the iterator.

    	returns Integer;


    Value(me: in out; Index: Integer from Standard)
    
	---Purpose: Returns the element of range Index.
    
    	returns any Item;
	---C++: return const&
	---C++: alias operator()


end Iterator;
