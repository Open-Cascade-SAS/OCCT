-- Created on: 1997-03-28
-- Created by: Philippe MANGIN
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

private class SearchSing from ChFi3d inherits FunctionWithDerivative from math

	---Purpose: F(t) = (C1(t) - C2(t)).(C1'(t) - C2'(t));

uses Curve from Geom

is
    Create(C1, C2 : Curve from Geom)
    returns SearchSing from ChFi3d;

    Value(me: in out; X: Real; F: out Real)
    	---Purpose: computes the value of the function <F> for the 
    	--          variable <X>. 
    	--          returns True if the computation was done successfully,
    	--          False otherwise.
    returns Boolean;
    
    Derivative(me: in out; X: Real; D: out Real)
         ---Purpose: computes the derivative <D> of the function 
         --          for the variable <X>.
    	--           Returns True if the calculation were successfully done, 
    	--           False otherwise.

    returns Boolean;    

    Values(me: in out; X: Real; F, D: out Real)
    	---Purpose: computes the value <F> and the derivative <D> of the 
    	--          function for the variable <X>.
    	--          Returns True if the calculation were successfully done,
    	--          False otherwise.

    returns Boolean;

fields
myC1 : Curve from Geom;
myC2 : Curve from Geom;
end SearchSing;
