-- Created on: 1994-02-14
-- Created by: model
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



generic class GenHSurface from Adaptor3d
    (TheSurface as Surface from Adaptor3d)
 
inherits HSurface from Adaptor3d 
    
	---Purpose: Generic class used to create a surface manipulated
      	--          with Handle from a surface described by the class Surface. 
	
uses

     Surface      from Adaptor3d


raises

    OutOfRange          from Standard,
    NoSuchObject        from Standard,
    DomainError         from Standard


is

    Create
    
	---Purpose: Creates an empty GenHSurface.
    	returns mutable GenHSurface from Adaptor3d; 
    

    Create(S: TheSurface)
    
	---Purpose: Creates a GenHSurface from a Surface.
    	returns mutable GenHSurface from Adaptor3d; 


    Set(me: mutable; S: TheSurface)
    
	---Purpose: Sets the field of the GenHSurface.
    	is static;

    --
    --  Access to the surface
    --  
    
    Surface(me) returns Surface from Adaptor3d;
	---Purpose: Returns a reference to the Surface inside the HSurface.
	--          This is redefined from HSurface, cannot be inline.
	--          
	---C++: return const &

    ChangeSurface(me : mutable)
    
	---Purpose: Returns the surface used to create the GenHSurface.
	--          
	---C++: return &
	---C++: inline

    	returns TheSurface;


fields

    mySurf: TheSurface is protected;

end GenHSurface;
