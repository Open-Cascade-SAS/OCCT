-- Created on: 1995-03-17
-- Created by: Dieter THIEMANN
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MakeGeometricCurveSet from TopoDSToStep inherits
    Root from TopoDSToStep

    ---Purpose: This class implements the mapping between a Shape 
    --          from TopoDS and a GeometricCurveSet from StepShape in order
    --          to create a GeometricallyBoundedWireframeRepresentation.
  
uses Shape from TopoDS,
     GeometricCurveSet from StepShape,
     FinderProcess from Transfer
          
raises NotDone from StdFail
     
is 

Create ( SH : Shape from TopoDS;
         FP : mutable FinderProcess from Transfer)
        returns MakeGeometricCurveSet;

Value (me) returns GeometricCurveSet from StepShape
    raises NotDone
    is static;
    ---C++: return const&

fields

    theGeometricCurveSet : GeometricCurveSet from StepShape;
    
    
end MakeGeometricCurveSet;    
