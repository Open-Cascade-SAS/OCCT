-- Created on: 1996-09-25
-- Created by: Christian CAILLET
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class SelectExplore  from IFSelect  inherits SelectDeduct

    ---Purpose : A SelectExplore determines from an input list of Entities,
    --           a list obtained by a way of exploration. This implies the
    --           possibility of recursive exploration : the output list is
    --           itself reused as input, etc...
    --           Examples : Shared Entities, can be considered at one level
    --           (immediate shared) or more, or max level
    --           
    --           Then, for each input entity, if it is not rejected, it can be
    --           either taken itself, or explored : it then produces a list.
    --           According to a level, either the produced lists or taken
    --           entities give the result (level one), or lists are themselves
    --           considered and for each item, is it taken or explored.
    --           
    --           Remark that rejection is just a safety : normally, an input
    --             entity is, either taken itself, or explored
    --           A maximum level can be specified. Else, the process continues
    --           until all entities have been either taken or rejected

uses AsciiString from TCollection, InterfaceModel, EntityIterator,  Graph

is

    Initialize (level : Integer);
    ---Purpose : Initializes a SelectExplore : the level must be specified on
    --           starting. 0 means all levels, 1 means level one only, etc...

    Level (me) returns Integer;
    ---Purpose : Returns the required exploring level

    RootResult (me; G : Graph) returns EntityIterator;
    ---Purpose : Returns the list of selected entities. Works by calling the
    --           method Explore on each input entity : it can be rejected,
    --           taken for output, or to explore. If the maximum level has not
    --           yet been attained, or if no max level is specified, entities
    --           to be explored are themselves used as if they were input

    Explore (me; level : Integer; ent : Transient; G : Graph;
    	     explored : in out EntityIterator)
    	returns Boolean  is deferred;
    ---Purpose : Analyses and, if required, Explores an entity, as follows :
    --           The explored list starts as empty, it has to be filled by this
    --           method.
    --           If it returns False, <ent> is rejected for result (this is to
    --               be used only as safety)
    --           If it returns True and <explored> remains empty, <ent> is
    --             taken itself for result, not explored
    --           If it returns True and <explored> is not empty, the content
    --             of this list is considered :
    --             If maximum level is attained, it is taken for result
    --             Else (or no max), each of its entity will be itself explored

    Label (me) returns AsciiString from TCollection;
    ---Purpose : Returns a text saying "(Recursive)" or "(Level nn)" plus
    --           specific criterium returned by ExploreLabel (see below)

    ExploreLabel (me) returns AsciiString from TCollection  is deferred;
    ---Purpose : Returns a text defining the way of exploration

fields

    thelevel : Integer;

end SelectExplore;
