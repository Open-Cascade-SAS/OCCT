-- File:	StepFEA_Curve3dElementRepresentation.cdl
-- Created:	Thu Dec 12 17:51:03 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class Curve3dElementRepresentation from StepFEA
inherits ElementRepresentation from StepFEA

    ---Purpose: Representation of STEP entity Curve3dElementRepresentation

uses
    HAsciiString from TCollection,
    HArray1OfRepresentationItem from StepRepr,
    RepresentationContext from StepRepr,
    HArray1OfNodeRepresentation from StepFEA,
    FeaModel3d from StepFEA,
    Curve3dElementDescriptor from StepElement,
    Curve3dElementProperty from StepFEA,
    ElementMaterial from StepElement

is
    Create returns Curve3dElementRepresentation from StepFEA;
	---Purpose: Empty constructor

    Init (me: mutable; aRepresentation_Name: HAsciiString from TCollection;
                       aRepresentation_Items: HArray1OfRepresentationItem from StepRepr;
                       aRepresentation_ContextOfItems: RepresentationContext from StepRepr;
                       aElementRepresentation_NodeList: HArray1OfNodeRepresentation from StepFEA;
                       aModelRef: FeaModel3d from StepFEA;
                       aElementDescriptor: Curve3dElementDescriptor from StepElement;
                       aProperty: Curve3dElementProperty from StepFEA;
                       aMaterial: ElementMaterial from StepElement);
	---Purpose: Initialize all fields (own and inherited)

    ModelRef (me) returns FeaModel3d from StepFEA;
	---Purpose: Returns field ModelRef
    SetModelRef (me: mutable; ModelRef: FeaModel3d from StepFEA);
	---Purpose: Set field ModelRef

    ElementDescriptor (me) returns Curve3dElementDescriptor from StepElement;
	---Purpose: Returns field ElementDescriptor
    SetElementDescriptor (me: mutable; ElementDescriptor: Curve3dElementDescriptor from StepElement);
	---Purpose: Set field ElementDescriptor

    Property (me) returns Curve3dElementProperty from StepFEA;
	---Purpose: Returns field Property
    SetProperty (me: mutable; Property: Curve3dElementProperty from StepFEA);
	---Purpose: Set field Property

    Material (me) returns ElementMaterial from StepElement;
	---Purpose: Returns field Material
    SetMaterial (me: mutable; Material: ElementMaterial from StepElement);
	---Purpose: Set field Material

fields
    theModelRef: FeaModel3d from StepFEA;
    theElementDescriptor: Curve3dElementDescriptor from StepElement;
    theProperty: Curve3dElementProperty from StepFEA;
    theMaterial: ElementMaterial from StepElement;

end Curve3dElementRepresentation;
