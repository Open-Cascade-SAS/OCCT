-- Created on: 1994-06-01
-- Created by: Christian CAILLET
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SetVersion5  from IGESSelect  inherits ModelModifier from IGESSelect

    ---Purpose : Sets IGES Version (coded in global parameter 23) to be at least
    --           IGES 5.1 . If it is older, it is set to IGES 5.1, and
    --           LastChangeDate (new Global n0 25) is added (current time)
    --           Else, it does nothing (i.e. changes neither IGES Version nor
    --           LastChangeDate)

uses AsciiString from TCollection,
     IGESModel, CopyTool, ContextModif

is

    Create returns mutable SetVersion5;
    ---Purpose : Creates an SetVersion5, which uses the system Date for Last
    --           Change Date

    Performing (me; ctx : in out ContextModif;
    	        target  : mutable IGESModel;
                TC      : in out CopyTool);
    ---Purpose : Specific action : only <target> is used : IGES Version (coded)
    --           is upgraded to 5.1 if it is older, and it this case the new
    --           global parameter 25 (LastChangeDate) is set to current time

    Label (me) returns AsciiString from TCollection;
    ---Purpose : Returns a text which is
    --           "Update IGES Version to 5.1"

end SetVersion5;
