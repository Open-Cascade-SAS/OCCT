-- Created on: 1991-04-03
-- Created by: Remi GILET
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class CircLin2dBisec

from GccAna

	---Purpose: Describes functions for building bisecting curves between a 2D line and a 2D circle.
    	-- A bisecting curve between a circle and a line is a curve
    	-- such that each of its points is at the same distance from
    	-- the circle and the line. It can be a parabola or a line,
    	-- depending of the relative position of the line and the
    	-- circle. The algorithm computes all the elementary curves which are solutions.
    	-- A CircLin2dBisec object provides a framework for:
    	-- -   defining the construction of the bisecting curves,
    	-- -   implementing the construction algorithm, and
    	-- -   consulting the result.


uses Lin2d  from gp,
     Circ2d from gp,
     Bisec  from GccInt
     
raises OutOfRange        from Standard,
       NotDone           from StdFail
       
is

Create(Circle  : Circ2d from gp;
       Line    : Lin2d  from gp) returns CircLin2dBisec;

    	---Purpose: Constructs bisecting curves between the circle Circle and the line Line. 

IsDone(me) returns Boolean from Standard
is static;

    	--- Purpose: Returns true (this construction algorithm never fails).
        
NbSolutions(me) returns Integer from Standard
raises NotDone
is static;
    	---Purpose:
    	-- Returns the number of curves, representing solutions computed by this algorithm.
    
ThisSolution(me                           ; 
    	     Index : Integer from Standard) returns Bisec from GccInt
raises OutOfRange, NotDone
is static;
    	---Purpose : Returns the solution number Index and raises OutOfRange 
    	--         exception if Index is greater than the number of solutions 
    	--    Exceptions
    	-- Standard_OutOfRange if Index is less than zero or
    	-- greater than the number of solutions computed by this algorithm.

fields

    WellDone : Boolean from Standard;
    	---Purpose: True if the algorithm succeeded.

    NbrSol   : Integer from Standard;
    	---Purpose: The number of possible solutions. We have to decide about the
    	--          status of the multiple solutions...

    circle   : Circ2d from gp;
    	---Purpose: The first argument used for ThisSolution.

    line   : Lin2d from gp;
    	---Purpose: The second argument used for ThisSolution.

end CircLin2dBisec;
