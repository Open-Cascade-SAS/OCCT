-- Created on: 1997-03-26
-- Created by: Christian CAILLET
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PresentationLayerUsage  from StepVisual    inherits TShared

    ---Purpose : Added from StepVisual Rev2 to Rev4

uses
     PresentationLayerAssignment from StepVisual,
     PresentationRepresentation from StepVisual

is

    Create returns PresentationLayerUsage;

    Init (me : mutable;
    	  aAssignment : PresentationLayerAssignment from StepVisual;
	  aPresentation : PresentationRepresentation from StepVisual);

    SetAssignment (me : mutable; aAssignment : PresentationLayerAssignment from StepVisual);
    Assignment (me) returns PresentationLayerAssignment from StepVisual;

    SetPresentation (me : mutable; aPresentation : PresentationRepresentation from StepVisual);
    Presentation (me) returns PresentationRepresentation from StepVisual;

fields

    theAssignment : PresentationLayerAssignment from StepVisual;
    thePresentation : PresentationRepresentation from StepVisual;

end PresentationLayerUsage;
