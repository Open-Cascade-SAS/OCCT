-- Created on: 2005-12-15
-- Created by: Julia GERASIMOVA
-- Copyright (c) 2005-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class EigenValuesSearcher from math
        ---Purpose: This class finds eigen values and vectors of
        --          real symmetric tridiagonal matrix

uses 
     
    Array1OfReal  from TColStd, 
    HArray1OfReal from TColStd, 
    HArray2OfReal from TColStd, 
    Vector        from math
    
raises 
 
    NotDone from StdFail

is 
    Create(Diagonal    : Array1OfReal from TColStd; 
    	   Subdiagonal : Array1OfReal from TColStd)
    returns EigenValuesSearcher
    raises NotDone;  -- if length(Subdiagonal) != length(Diagonal)-1 
    
    IsDone(me)
     	---Purpose: Returns Standard_True if computation is performed 
        --          successfully.
    returns Boolean from Standard;

    Dimension(me)
     	---Purpose: Returns the dimension of matrix
    returns Integer from Standard;

    EigenValue(me; Index : Integer from Standard)
     	---Purpose: Returns the Index_th eigen value of matrix
        --          Index must be in [1, Dimension()]
    returns Real from Standard;

    EigenVector(me; Index : Integer from Standard)
     	---Purpose: Returns the Index_th eigen vector of matrix
        --          Index must be in [1, Dimension()]
    returns Vector from math;
     
fields 

    myDiagonal    : HArray1OfReal from TColStd;
    mySubdiagonal : HArray1OfReal from TColStd;  
    
    myIsDone       : Boolean from Standard; 
    myN            : Integer from Standard;
    myEigenValues  : HArray1OfReal from TColStd; 
    myEigenVectors : HArray2OfReal from TColStd;

end EigenValuesSearcher;
