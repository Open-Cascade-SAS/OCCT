-- Created on: 1994-11-25
-- Created by: Frederic MAUPAS
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package TopoDSToStep

    ---Purpose: This package implements the mapping between CAS.CAD
    --  Shape representation and AP214 Shape Representation.
    --  The target schema is pms_c4 (a subset of AP214)
    --  
    --  How to use this Package :
    --  
    --  Entry point are context dependent. It can be :
    --     MakeManifoldSolidBrep
    --     MakeBrepWithVoids
    --     MakeFacetedBrep
    --     MakeFacetedBrepAndBrepWithVoids
    --     MakeShellBasedSurfaceModel
    --  Each of these classes call the Builder
    --  The class tool centralizes some common informations.   

uses TopoDS, StdFail, TCollection, TColStd, TopTools, Transfer, MoniTool,
     BRepTools, TopLoc, GeomAbs, Geom2d, Geom, gp,
     StepGeom, StepShape

is

--  ------------------------------------------------------
--  Enumeration
--  ------------------------------------------------------

    enumeration BuilderError is
    	BuilderDone,
	NoFaceMapped,
	BuilderOther
    end BuilderError;
    
    enumeration MakeFaceError is
    	FaceDone,
	InfiniteFace,
	NonManifoldFace,
	NoWireMapped,
    	FaceOther
    end MakeFaceError;
    
    enumeration MakeWireError is
    	WireDone,
	NonManifoldWire,
    	WireOther
    end MakeWireError;
    
    enumeration MakeEdgeError is
    	EdgeDone,
	NonManifoldEdge,
    	EdgeOther
    end MakeEdgeError;
    
    enumeration MakeVertexError is
    	VertexDone,
    	VertexOther
    end MakeVertexError;
    
    enumeration FacetedError is
	FacetedDone,    
    	SurfaceNotPlane,
	PCurveNotLinear
    end FacetedError;

--  ------------------------------------------------------
--  Package Classes
--  ------------------------------------------------------

    private deferred class Root;

    class MakeManifoldSolidBrep;

    class MakeBrepWithVoids;

    class MakeFacetedBrep;

    class MakeFacetedBrepAndBrepWithVoids;

    class MakeShellBasedSurfaceModel;

    class MakeGeometricCurveSet;
    
    class Builder;
    
    class WireframeBuilder;
    
    class Tool;
    
    class FacetedTool;
    
    class MakeStepFace;
    
    class MakeStepWire;
    
    class MakeStepEdge;
    
    class MakeStepVertex;
    
--    private class DirectModification;
--    private class ConicalSurfModif;
    
--  ------------------------------------------------------
--  Instanciated Class
--  ------------------------------------------------------

--    class DataMapOfShape instantiates
--    	  DataMap from TCollection 
--    	    (Shape                         from TopoDS,
--    	     TopologicalRepresentationItem from StepShape,
--	     ShapeMapHasher                from TopTools);

--  ------------------------------------------------------
--  Package Method
--  ------------------------------------------------------

    DecodeBuilderError(E : BuilderError from TopoDSToStep)
    	returns HAsciiString from TCollection;   
   
    DecodeFaceError(E : MakeFaceError from TopoDSToStep)
    	returns HAsciiString from TCollection;
	
    DecodeWireError(E : MakeWireError from TopoDSToStep)
    	returns HAsciiString from TCollection;   
   
    DecodeEdgeError(E : MakeEdgeError from TopoDSToStep)
    	returns HAsciiString from TCollection;
	
    DecodeVertexError(E : MakeVertexError from TopoDSToStep)
    	returns HAsciiString from TCollection;
	
--    DirectFaces(S : Shape from TopoDS)
--    	returns Shape from TopoDS;
	---Purpose: Returns a new shape without undirect surfaces.
	
    AddResult (FP: FinderProcess from Transfer;
     	       Shape: Shape from TopoDS;
	       entity: Transient from Standard);
	---Purpose: Adds an entity into the list of results (binders) for
	--          shape stored in FinderProcess

    AddResult (FP: FinderProcess from Transfer;
     	       Tool: Tool from TopoDSToStep);
	---Purpose: Adds all entities recorded in Tool into the map of results
	--          (binders) stored in FinderProcess

end TopoDSToStep;
