-- Created on: 1993-07-15
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Face from DBRep inherits TShared from MMgt
	---Purpose: Display of a face. Face + Array of iso + color.
uses
    Face            from TopoDS,
    IsoType         from GeomAbs,
    Array1OfInteger from TColStd,
    Array1OfReal    from TColStd,
    Color           from Draw

is
    Create (F : Face from TopoDS; 
    	    N : Integer;
    	    C : Color from Draw)
    returns Face from DBRep;
	---Purpose: N is the number of iso intervals.
    
    Face(me) returns Face from TopoDS
	---C++: return const &
	---C++: inline
    is static;

    Face(me : mutable; F : Face from TopoDS)
	---C++: inline
    is static;
    
    NbIsos(me) returns Integer
	---C++: inline
    is static;

    Iso(me : mutable; 
    	I           : Integer; 
    	T           : IsoType from GeomAbs; 
    	Par, T1, T2 : Real)
	---C++: inline
    is static;

    GetIso(me;
    	   I           : Integer; 
    	   T           : out IsoType from GeomAbs; 
    	   Par, T1, T2 : out Real)
	---C++: inline
    is static;

    Color(me) returns Color from Draw
	---C++: return const &
	---C++: inline
    is static;

    Color(me : mutable; C : Color from Draw)
	---C++: inline
    is static;
    
fields
    myFace   : Face            from TopoDS;
    myColor  : Color           from Draw;
    myTypes  : Array1OfInteger from TColStd;
    myParams : Array1OfReal    from TColStd;

end Face;
