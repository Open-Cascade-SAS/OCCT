-- Created on: 1993-03-10
-- Created by: JCV
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class SurfaceOfRevolution from Geom inherits SweptSurface from Geom

        ---Purpose : Describes a surface of revolution (revolved surface).
    	-- Such a surface is obtained by rotating a curve (called
    	-- the "meridian") through a complete revolution about
    	-- an axis (referred to as the "axis of revolution"). The
    	-- curve and the axis must be in the same plane (the
    	-- "reference plane" of the surface).
    	-- Rotation around the axis of revolution in the
    	-- trigonometric sense defines the u parametric
    	-- direction. So the u parameter is an angle, and its
    	-- origin is given by the position of the meridian on the surface.
    	-- The parametric range for the u parameter is: [ 0, 2.*Pi ]
    	-- The v parameter is that of the meridian.
    	-- Note: A surface of revolution is built from a copy of the
    	-- original meridian. As a result the original meridian is
    	-- not modified when the surface is modified.
    	-- The form of a surface of revolution is typically a
    	-- general revolution surface
    	-- (GeomAbs_RevolutionForm). It can be:
    	-- - a conical surface, if the meridian is a line or a
    	--   trimmed line (GeomAbs_ConicalForm),
    	-- - a cylindrical surface, if the meridian is a line or a
    	--   trimmed line parallel to the axis of revolution
    	--   (GeomAbs_CylindricalForm),
    	-- - a planar surface if the meridian is a line or a
    	--   trimmed line perpendicular to the axis of revolution
    	--   of the surface (GeomAbs_PlanarForm),
    	-- - a toroidal surface, if the meridian is a circle or a
    	--   trimmed circle (GeomAbs_ToroidalForm), or
    	-- - a spherical surface, if the meridian is a circle, the
    	--   center of which is located on the axis of the
    	--   revolved surface (GeomAbs_SphericalForm).
    	--   Warning
    	-- Be careful not to construct a surface of revolution
    	-- where the curve and the axis or revolution are not
    	-- defined in the same plane. If you do not have a
    	-- correct configuration, you can correct your initial
    	-- curve, using a cylindrical projection in the reference plane.
        
        
        
uses Ax1         from gp, 
     Ax2         from gp,
     Dir         from gp,
     Pnt         from gp,
     Trsf        from gp,
     GTrsf2d     from gp,
     Vec         from gp,
     Curve       from Geom,
     Geometry    from Geom,
     Shape       from GeomAbs,
    BSplineCurve from Geom  

raises ConstructionError   from Standard,
       RangeError          from Standard, 
       UndefinedDerivative from Geom
 

is


  Create (C : Curve; A1 : Ax1)   returns mutable SurfaceOfRevolution;
        ---Purpose :
        --  C : is the meridian  or the referenced curve.
        --  A1 is the axis of revolution. 
        --  The form of a SurfaceOfRevolution can be :
        --  . a general revolution surface (RevolutionForm),
        --  . a conical surface if the meridian is a line or a trimmed line
        --    (ConicalForm),
        --  . a cylindrical surface if the meridian is a line or a trimmed
        --    line parallel to the revolution axis (CylindricalForm),
        --  . a planar surface if the meridian is a line perpendicular to
        --    the revolution axis of the surface (PlanarForm).  
        --  . a spherical surface,
        --  . a toroidal surface,
        --  . a quadric surface.
        -- Warnings :
        --  It is not checked that the curve C is planar and that the
        --  surface axis is in the plane of the curve.
        --  It is not checked that the revolved curve C doesn't 
        --  self-intersects.


  SetAxis (me : mutable; A1 : Ax1);
        ---Purpose : Changes the axis of revolution.
        -- Warnings :
        --  It is not checked that the axis is in the plane of the 
        --  revolved curve.


  SetDirection (me : mutable; V : Dir);
        ---Purpose : Changes the direction of the revolution axis.
        -- Warnings :
        --  It is not checked that the axis is in the plane of the 
        --  revolved curve.



  SetBasisCurve (me : mutable; C : Curve);
        ---Purpose : Changes the revolved curve of the surface.
        -- Warnings :
        --  It is not checked that the curve C is planar and that the
        --  surface axis is in the plane of the curve.
        --  It is not checked that the revolved curve C doesn't 
        --  self-intersects.


  SetLocation (me : mutable; P : Pnt);
        ---Purpose : Changes the location point of the revolution axis.
        -- Warnings :
        --  It is not checked that the axis is in the plane of the 
        --  revolved curve.


  Axis (me)  returns Ax1;
        ---Purpose : Returns the revolution axis of the surface.


  Location (me)  returns Pnt;
        ---Purpose :
        --  Returns the location point of the axis of revolution.
    	---C++: return const&


  ReferencePlane (me)   returns Ax2
        ---Purpose :
        --  Computes the position of the reference plane of the surface
        --  defined by the basis curve and the symmetry axis.
        --  The location point is the location point of the revolution's
        --  axis, the XDirection of the plane is given by the revolution's
        --  axis and the orientation of the normal to the plane is given
        --  by the sense of revolution.
     raises ConstructionError;
        ---Purpose :
        --  Raised if the revolved curve is not planar or if the revolved 
        --  curve and the symmetry axis are not in the same plane or if 
        --  the maximum of distance between the axis and the revolved
        --  curve is lower or equal to Resolution from gp.


  UReverse (me : mutable);
    	---Purpose : Changes the orientation of this surface of revolution
    	-- in the u  parametric direction. The bounds of the
    	-- surface are not changed but the given parametric
    	-- direction is reversed. Hence the orientation of the
    	-- surface is reversed.
    	-- As a consequence:
    	-- - UReverse reverses the direction of the axis of
    	--   revolution of this surface,


  UReversedParameter ( me; U : Real) returns Real;
    	---Purpose: Computes the u  parameter on the modified
    	-- surface, when reversing its u  parametric
    	-- direction, for any point of u parameter U  on this surface of revolution.
    	-- In the case of a revolved surface:
    	-- - UReversedParameter returns 2.*Pi - U

  
  VReverse (me : mutable);
       	---Purpose : Changes the orientation of this surface of revolution
    	-- in the v parametric direction. The bounds of the
    	-- surface are not changed but the given parametric
    	-- direction is reversed. Hence the orientation of the
    	-- surface is reversed.
    	-- As a consequence:
    	-- - VReverse reverses the meridian of this surface of revolution. 

  VReversedParameter (me; V : Real) returns Real;
	---Purpose: Computes the  v parameter on the modified
    	-- surface, when reversing its  v parametric
    	-- direction, for any point of v parameter V on this surface of revolution.
    	-- In the case of a revolved surface:
    	-- - VReversedParameter returns the reversed
    	--   parameter given by the function
    	--   ReversedParameter called with V on the meridian.

  TransformParameters(me; U,V : in out Real; T : Trsf from gp)
	---Purpose: Computes the  parameters on the  transformed  surface for
	--          the transform of the point of parameters U,V on <me>.
	--          
	--          me->Transformed(T)->Value(U',V')
	--          
	--          is the same point as
	--          
	--          me->Value(U,V).Transformed(T)
	--          
	--          Where U',V' are the new values of U,V after calling
	--          
	--          me->TranformParameters(U,V,T)
	--          
	--          This methods multiplies V by 
	--          BasisCurve()->ParametricTransformation(T)
     is redefined;  

  ParametricTransformation(me; T : Trsf from gp) returns GTrsf2d from gp
	---Purpose: Returns a 2d transformation  used to find the  new
	--          parameters of a point on the transformed surface.
	--          
	--          me->Transformed(T)->Value(U',V')
	--          
	--          is the same point as
	--          
	--          me->Value(U,V).Transformed(T)
	--          
	--          Where U',V' are  obtained by transforming U,V with
	--          th 2d transformation returned by
	--          
	--          me->ParametricTransformation(T)
	--          
	--          This  methods  returns  a scale  centered  on  the
	--          U axis with BasisCurve()->ParametricTransformation(T)
     is redefined;  
  
  Bounds (me; U1, U2, V1, V2 : out Real);
        ---Purpose : Returns the parametric bounds U1, U2 , V1 and V2 of this surface.
    	-- A surface of revolution is always complete, so U1 = 0, U2 = 2*PI.


  IsUClosed (me) returns Boolean;
        ---Purpose : IsUClosed always returns true.


  IsVClosed (me)  returns Boolean;
        ---Purpose : IsVClosed returns true if the meridian of this
    	--   surface of revolution is closed.


  IsCNu (me; N : Integer)  returns Boolean;
        ---Purpose : IsCNu always returns true.


  IsCNv (me; N : Integer)  returns Boolean
        ---Purpose : IsCNv returns true if the degree of continuity of the
    	--   meridian of this surface of revolution is at least N.
     raises RangeError;
        ---Purpose : Raised if N < 0.


  IsUPeriodic (me)   returns Boolean;
        ---Purpose : Returns True.


  IsVPeriodic (me)  returns Boolean;
        ---Purpose :  IsVPeriodic returns true if the meridian of this
    	--   surface of revolution is periodic.


  UIso (me; U : Real)   returns mutable Curve;
    	---Purpose :  Computes the U isoparametric curve of this surface
    	-- of revolution. It is the curve obtained by rotating the
    	-- meridian through an angle U about the axis of revolution.


  VIso (me; V : Real)  returns mutable Curve;
    	---Purpose :  Computes the U isoparametric curve of this surface
    	-- of revolution. It is the curve obtained by rotating the
    	-- meridian through an angle U about the axis of revolution.


  D0 (me; U, V : Real; P : out Pnt);
        ---Purpose :  Computes the  point P (U, V) on the surface.
        --  U is the angle of the rotation around the revolution axis.
        --  The direction of this axis gives the sense of rotation.
        --  V is the parameter of the revolved curve.

  
  D1 (me; U, V : Real; P : out Pnt; D1U, D1V : out Vec)
        ---Purpose :
        --  Computes the current point and the first derivatives 
        --  in the directions U and V.
     raises UndefinedDerivative;
        ---Purpose : Raised if the continuity of the surface is not C1.


  D2 (me; U, V : Real; P : out Pnt; D1U, D1V, D2U, D2V, D2UV : out Vec)
        ---Purpose :
        --  Computes the current point, the first and the second derivatives
        --  in the directions U and V.
     raises UndefinedDerivative;
        ---Purpose : Raised if the continuity of the surface is not C2.


  D3 (me; U, V : Real; P : out Pnt; 
      D1U, D1V, D2U, D2V, D2UV, D3U, D3V, D3UUV, D3UVV : out Vec)
        ---Purpose :
        --  Computes the current point, the first,the second and the third 
        --  derivatives in the directions U and V.
     raises UndefinedDerivative;
        ---Purpose : Raised if the continuity of the surface is not C3.


  DN (me; U, V : Real; Nu, Nv : Integer)
        ---Purpose :
        --  Computes the derivative of order Nu in the direction u and 
        --  Nv in the direction v.
     returns Vec
     raises UndefinedDerivative,
        ---Purpose : 
        --  Raised if the continuity of the surface is not CNu in the u
        --  direction and CNv in the v direction.
            RangeError;
        ---Purpose : Raised if Nu + Nv < 1 or Nu < 0 or Nv < 0.



    	---Purpose : The following  functions  evaluates the  local 
    	-- derivatives on surface. Useful to manage discontinuities 
	-- on the surface. 
	--           if    Side  =  1  ->  P  =  S( U+,V ) 
        --           if    Side  = -1  ->  P  =  S( U-,V ) 
    	--           else  P  is betveen discontinuities   
	--           can be evaluated using methods  of  
    	--           global evaluations    P  =  S( U ,V )      
   
  LocalD0 (me; U, V : Real; USide : Integer;
    	       P : out Pnt);
 
  LocalD1 (me; U, V : Real;  USide : Integer;
          P : out Pnt; D1U, D1V : out Vec);
 
  LocalD2 (me; U, V : Real; USide : Integer;
           P : out Pnt; D1U, D1V, D2U, D2V, D2UV : out Vec);
 
  LocalD3 (me; U, V : Real; USide : Integer;
           P : out Pnt; D1U, D1V, D2U, D2V, D2UV, D3U, D3V, D3UUV, D3UVV :
           out Vec);
  
  LocalDN (me; U, V : Real; USide : Integer; 
           Nu, Nv : Integer)
     returns Vec;

  Transform (me : mutable; T : Trsf);
    	---Purpose: Applies the transformation T to this surface of revolution.
   Copy (me)  returns mutable like me;
    	---Purpose: Creates a new object which is a copy of this surface of revolution.
fields

  loc  : Pnt;

end;
