-- Created on: 1994-09-29
-- Created by: Dieter THIEMANN
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package UnitsMethods

uses

    Standard, Geom, Geom2d
    
is

    InitializeFactors(LengthFactor :     Real from Standard;
                      PlaneAngleFactor : Real from Standard;
                      SolidAngleFactor : Real from Standard);

       ---Purpose: Initializes the 3 factors for the conversion of
       --          units

    LengthFactor       
    	returns   Real from Standard;

    PlaneAngleFactor   
    	returns   Real from Standard;

    SolidAngleFactor   
    	returns   Real from Standard;

    Set3dConversion(B : Boolean from Standard);
    
    Convert3d          
    	returns   Boolean from Standard;
    
    RadianToDegree(C : Curve from Geom2d; 
    	    	   S : Surface from Geom)
    	returns Curve from Geom2d;
		   
    DegreeToRadian(C : Curve from Geom2d; 
    	    	   S : Surface from Geom)
    	returns Curve from Geom2d;

    MirrorPCurve(C : Curve from Geom2d)
	returns Curve from Geom2d;

    GetLengthFactorValue (param: Integer) returns Real;
    	---Purpose: Returns value of unit encoded by parameter param
        --          (integer value denoting unit, as described in IGES
        --          standard) in millimeters
	
    GetCasCadeLengthUnit returns Real;
    	---Purpose: Returns value of current internal unit for CASCADE
	--          in millemeters
	
    SetCasCadeLengthUnit (param: Integer);
    	---Purpose: Sets value of current internal unit for CASCADE
	--          by parameter param (integer value denoting unit, 
        --          as described in IGES standard) 
	--          GetCasCadeLengthUnit() will then return value 
	--          equal to GetLengthFactorValue(param)
	
end UnitsMethods;
