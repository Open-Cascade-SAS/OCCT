-- Created on: 2001-04-24
-- Created by: Christian CAILLET
-- Copyright (c) 2001-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class ValueQualifier  from StepShape    inherits SelectType  from StepData

    ---Purpose : Added for Dimensional Tolerances

uses
    PrecisionQualifier from StepShape,
    TypeQualifier from StepShape

is

    Create returns ValueQualifier from StepShape;

    CaseNum (me; ent : Transient) returns Integer;
    ---Purpose : Recognizes a kind of ValueQualifier Select Type :
    --           1 -> PrecisionQualifier from StepShape
    --           2 -> TypeQualifier from StepShape
    --           3 -> UnceraintyQualifier .. not yet implemented

    PrecisionQualifier (me) returns PrecisionQualifier from StepShape;
    ---Purpose : Returns Value as PrecisionQualifier

    TypeQualifier (me) returns TypeQualifier from StepShape;
    ---Purpose : Returns Value as TypeQualifier

end ValueQualifier;
