-- File:	IGESGeom_ToolTabulatedCylinder.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolTabulatedCylinder  from IGESGeom

    ---Purpose : Tool to work on a TabulatedCylinder. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses TabulatedCylinder from IGESGeom,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolTabulatedCylinder;
    ---Purpose : Returns a ToolTabulatedCylinder, ready to work


    ReadOwnParams (me; ent : mutable TabulatedCylinder;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : TabulatedCylinder;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : TabulatedCylinder;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a TabulatedCylinder <ent>, from
    --           its specific (own) parameters

    DirChecker (me; ent : TabulatedCylinder) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : TabulatedCylinder;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : TabulatedCylinder; entto : mutable TabulatedCylinder;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : TabulatedCylinder;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolTabulatedCylinder;
