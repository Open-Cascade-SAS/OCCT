-- Created on: 1991-01-21
-- Created by: Christophe MARION
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

private class ItemLocation from TopLoc

	---Purpose: An ItemLocation is an elementary coordinate system
	--          in a Location.
	--          
	--          The  ItemLocation     contains :
	--          
	--          * The elementary Datum.
	--          
	--          * The exponent of the elementary Datum.
	--          
	--          * The transformation associated to the composition.
	--          

uses
    Datum3D   from TopLoc,
    Trsf      from gp,
    TrsfPtr from TopLoc
    
is
    Create(D : Datum3D      from TopLoc; 
    	   P : Integer      from Standard;
           fromTrsf : Boolean from Standard = Standard_False) returns ItemLocation from TopLoc;
	---Purpose: Sets the elementary Datum to <D>
	--          Sets the exponent to <P>

    Create(anOther : ItemLocation from TopLoc) returns ItemLocation from TopLoc;
    
    Assign(me : in out; anOther : ItemLocation from TopLoc) returns ItemLocation from TopLoc;
    ---C++: alias operator=
    ---C++: return &

    Destroy(me : in out);
    ---C++: alias ~

fields
    myDatum  : Datum3D   from TopLoc;
    myPower  : Integer   from Standard;
    myTrsf   : TrsfPtr   from TopLoc;

friends
    class Location from TopLoc
    
end ItemLocation;
