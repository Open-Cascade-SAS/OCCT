-- Created by: Tanya COOL
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class AspectHidingPoly from Prs2d inherits AspectRoot from Prs2d

 ---Purpose: defines the attributes when drawing a hiding 
 --          polyhedral simplification Presentation.
uses

  NameOfColor from Quantity,
  TypeOfLine from Aspect,
  WidthOfLine from Aspect 

is
 
    Create ( HidingColorInd: NameOfColor from Quantity;
             FrameColorInd:  NameOfColor from Quantity;
             FrameTypeInd:   TypeOfLine from Aspect;
             FrameWidthInd:  WidthOfLine from Aspect)
	   returns mutable AspectHidingPoly from Prs2d;
	    
    SetHidingColor (me: mutable; aColorInd:      NameOfColor from Quantity ) is static;
    SetFrameColor  (me: mutable; aFrameColorInd: NameOfColor from Quantity ) is static;
    SetFrameType   (me: mutable; aFrameTypeInd:  TypeOfLine from Aspect) is static;
    SetFrameWidth  (me: mutable; aFrameWidthInd: WidthOfLine from Aspect ) is static;

    Values( me;
	      HidingColorInd: out NameOfColor from Quantity;
            FrameColorInd:  out NameOfColor from Quantity;
            FrameTypeInd:   out TypeOfLine from Aspect;
            FrameWidthInd:  out WidthOfLine from Aspect );

 fields
    
    myHidingColorInd: NameOfColor from Quantity;
    myFrameColorInd:  NameOfColor from Quantity;
    myFrameTypeInd:   TypeOfLine  from Aspect;
    myFrameWidthInd:  WidthOfLine from Aspect; 

end AspectHidingPoly from Prs2d;
