-- Created on: 1993-05-07
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class WPointInterIterator from TopOpeBRep

uses

    LineInter from TopOpeBRep,
    PLineInter from TopOpeBRep,
    WPointInter from TopOpeBRep
    
is

    -- ==========================
    -- Restriction Point iterator
    -- ==========================

    Create returns WPointInterIterator from TopOpeBRep;
    Create (LI : LineInter from TopOpeBRep) 
    returns WPointInterIterator from TopOpeBRep; 

    Init(me:in out; LI : LineInter from TopOpeBRep) is static;
    Init(me:in out) is static;
    More(me) returns Boolean from Standard is static;
    Next(me:in out) is static;
 
    CurrentWP(me:in out) returns WPointInter from TopOpeBRep 
    ---C++: return const &
    is static;

    PLineInterDummy(me) returns PLineInter from TopOpeBRep;

fields

    myLineInter : PLineInter from TopOpeBRep;
    myWPointIndex : Integer from Standard;
    myWPointNb : Integer from Standard;
    
end WPointInterIterator from TopOpeBRep;
