-- Created on: 2000-08-11
-- Created by: Andrey BETENEV
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package XCAFPrs 

    ---Purpose: Presentation (visualiation, selection etc.) tools for
    --          DECAF documents

uses
    Quantity,
    TCollection,
    TopAbs,
    TopLoc,
    TopoDS,
    TopTools,
    Graphic3d,
    Prs3d,
    PrsMgr,
    TPrsStd,
    AIS,
    TDF,
    XCAFDoc

is

    class Driver;
    	---Purpose: Implements a presentation driver for DECAF

    class AISObject;
    	---Purpose: Implements an interactive object for DECAF

    class Style;
        ---Purpose: Object representing a set of style settings
	
    class DataMapOfShapeStyle instantiates
    	DataMap from TCollection(Shape from TopoDS,
	    	    	    	 Style from XCAFPrs,
                                 ShapeMapHasher from TopTools);

    class DataMapOfStyleShape instantiates
    	DataMap from TCollection(Style from XCAFPrs,
                                 Shape from TopoDS,
	    	    	    	 Style from XCAFPrs);

    class DataMapOfStyleTransient instantiates
    	DataMap from TCollection(Style from XCAFPrs,
                                 Transient from Standard,
	    	    	    	 Style from XCAFPrs);

    ---Methods: Work with styles of the document
    
    CollectStyleSettings (L: Label from TDF;
			  loc: Location from TopLoc;
			  settings: in out DataMapOfShapeStyle from XCAFPrs);
    	---Purpose: Collect styles defined for shape on label L
    	--          and its components and subshapes and fills a map of 
	--          shape - style correspondence
	--          The location <loc> is for internal use, it 
	--          should be Null location for external call
	
    DispatchStyles (shape: Shape from TopoDS; 
    	    	    settings: DataMapOfShapeStyle from XCAFPrs; 
		    items: in out DataMapOfStyleShape from XCAFPrs;
		    DefStyle: Style from XCAFPrs;
		    force: Boolean = Standard_True;
    	    	    context: ShapeEnum from TopAbs = TopAbs_SHAPE)
    returns Boolean;
    	---Purpose: Iterates on shape (recursively) and splits it
	--          on parts each of which has its own style
	--          (basing on settings collected by CollectStyleSettings())
	--          The DefStyle is default style applied to a shape if
	--          no specific style assignment is applied to it
	--          If force is True, the <shape> is added to a map
	--          even if no styles are redefined for it or its
	--          subshapes
	--          The context is for internal use, it indicates
	--          the type of the shape to which <shape> belongs

    SetViewNameMode ( viewNameMode: Boolean from Standard);

    	---Purpose: Set ViewNameMode for indicate display names or not.
	
    GetViewNameMode returns Boolean;

        	   	    	
end XCAFPrs;
