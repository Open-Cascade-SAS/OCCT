-- Created on: 1991-01-10
-- Created by: Arnaud BOUZY
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class NamedExpression from Expr
    
inherits GeneralExpression from Expr  

    ---Purpose: Describe an expression used  by its name (as constants 
    --          or variables). A single reference is made to a 
    --          NamedExpression in every Expression (i.e. a 
    --          NamedExpression is shared).

uses AsciiString from TCollection


is

    GetName(me)
    returns AsciiString
    ---C++: return const &
    ---Level: Advanced
    is static;

    SetName(me : mutable; name : AsciiString)
    ---Level: Internal
    is static;

    IsShareable(me)
    ---Purpose: Tests if <me> can be shared by one or more expressions 
    --          or must be copied. This method redefines to a True 
    --          value the GeneralExpression method.
    returns Boolean
    is redefined;
    
    IsIdentical(me; Other : GeneralExpression)
    ---Purpose: Tests if <me> and <Other> define the same expression.
    --          This method does not include any simplification before
    --          testing.
    returns Boolean;

    String(me)
    ---Purpose: returns a string representing <me> in a readable way.
    returns AsciiString from TCollection;

fields

    myName : AsciiString;

end NamedExpression;
