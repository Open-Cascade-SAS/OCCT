-- Created on: 1993-06-22
-- Created by: Jean Louis FRENKEL, Gerard GRAS
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


-- Modified: TCL G002A, 28-11-00, new section "inquire methods"


class InfiniteLine from Graphic2d inherits Line from Graphic2d

	---Version:

	---Purpose: The primitive InfiniteLine

	---Keywords: Primitive, InfiniteLine
	---Warning:
	---References:

uses
	Drawer          from Graphic2d,
	GraphicObject	from Graphic2d,
	Length          from Quantity, 
	FStream         from Aspect,
	IFStream	from Aspect


raises
	InfiniteLineDefinitionError	from Graphic2d

is
	-------------------------
	-- Category: Constructors
	-------------------------

	Create (aGraphicObject: GraphicObject from Graphic2d;
		X, Y, DX, DY: Length from Quantity)
	returns mutable InfiniteLine from Graphic2d
	---Level: Public
	---Purpose: Creates an infinite line.
	--	    The reference point is <X>, <Y>.
	--	    The slope is <DX>, <DY>.
	--  Warning: Raises InfiniteLineDefinitionError if the
	--          <DX> and <DY> are null.
	raises InfiniteLineDefinitionError from Graphic2d;

	--------------------------
	-- Category: Draw and Pick
	--------------------------

	Draw (me : mutable; aDrawer: Drawer from Graphic2d)
	is static protected;
	---Level: Internal
	---Purpose: Draws the infinite line <me>.

	Pick (me : mutable; X, Y: ShortReal from Standard;
		aPrecision: ShortReal from Standard;
		aDrawer: Drawer from Graphic2d)
	returns Boolean from Standard is static protected;
	---Level: Internal
	---Purpose: Returns Standard_True if the infinite line <me> is picked,
	--	    Standard_False if not.

	--------------------------------------
	-- Category: Inquire methods
	--------------------------------------

    Reference( me; X, Y: out Length from Quantity );  
	---Level: Public
	---Purpose: returns the coordinates of the reference point
	
	Slope( me; dX, dY: out Length from Quantity );
	---Level: Public
	---Purpose: returns the slope <dX>, <dY>

	----------------------------------------------------------------------

	Save( me; aFStream: in out FStream from Aspect ) is virtual;
	Retrieve(myclass; anIFStream: in out IFStream from Aspect;
		aGraphicObject: GraphicObject from Graphic2d);
fields

	myX:	ShortReal from Standard;
	myY:	ShortReal from Standard;
	myDX:	ShortReal from Standard;
	myDY:	ShortReal from Standard;

end InfiniteLine from Graphic2d;
