-- Created on: 1998-07-22
-- Created by: Philippe MANGIN
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

private  class Section from BRepFill 

	---Purpose: To store section definition
uses 
    Shape  from TopoDS, 
    Wire   from TopoDS,
    Vertex from TopoDS  

is 
  Create returns Section from BRepFill;  
   
  Create (Profile : Shape  from TopoDS;   
          V       : Vertex from TopoDS; 
    	  WithContact    :  Boolean ; 
          WithCorrection :  Boolean) 
  returns Section from BRepFill;  
   
  Set(me  :  in  out;  IsLaw  :  Boolean); 
   
  Wire(me)   
  ---C++: return const & 
  ---C++: inline    
  returns  Wire  from  TopoDS; 
   
  Vertex(me)   
  ---C++: return const & 
  ---C++: inline    
  returns  Vertex  from  TopoDS;   

  IsLaw(me)   
   ---C++: inline
  returns  Boolean; 
   
  WithContact(me)  
   ---C++: inline
  returns  Boolean; 
   
  WithCorrection(me)  
   ---C++: inline
  returns  Boolean;  
   
     

fields
    wire    :  Wire  from  TopoDS; 
    vertex  :  Vertex from TopoDS;       
    islaw   :  Boolean;
    contact :  Boolean; 
    correction:Boolean; 
end Section;
