-- Created on: 1992-05-27
-- Created by: Remi LEQUETTE
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class TEdge from PBRep inherits TEdge from PTopoDS

	---Purpose: The TEdge from PBRep is  inherited from  the  TEdge
	--          from TopoDS. It contains the geometric data.
	--          
	--          The TEdge contains :
	--           
	--           * Flags : SameParameter, SameRange, Degenerated
	--          
	--           * A tolerance.
	--           
	--           * A list of representations.
	--           

uses
    CurveRepresentation       from PBRep

is
    Create returns TEdge from PBRep;
	---Purpose: Creates an empty TEdge.
    	---Level: Internal 

    Tolerance(me) returns Real
    is static;
    	---Level: Internal 
    	
    Tolerance(me : mutable; T : Real)
    is static;
    	---Level: Internal 
    
    SameParameter(me) returns Boolean
    is static;
    	---Level: Internal 
    
    SameParameter(me : mutable; S : Boolean)
    is static;
    	---Level: Internal 
    
    SameRange(me) returns Boolean
    is static;
    	---Level: Internal 
    
    SameRange(me : mutable; S : Boolean)
    is static;
    	---Level: Internal 
    
    Degenerated(me) returns Boolean
    is static;
    	---Level: Internal 
    
    Degenerated(me : mutable; S : Boolean)
    is static;
    	---Level: Internal 
    
    Curves(me) returns CurveRepresentation from PBRep
    is static;
    	---Level: Internal 
    
    Curves(me : mutable; C : CurveRepresentation from PBRep)
    is static;
    	---Level: Internal 
    

fields

    myTolerance     : Real;
    myFlags         : Integer;
    myCurves        : CurveRepresentation from PBRep;

end TEdge;
