-- Created on: 1991-11-18
-- Created by: Remi GILET
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


generic class ParGenCurve from GccGeo (TheCurve as any)

    ---Purpose: Definition of a virtual curve.

uses Pnt2d  from gp,
     Vec2d  from gp
     
is

Create returns ParGenCurve;

Create(C : TheCurve) returns ParGenCurve;

Create(C : TheCurve               ;
       D : Real     from Standard ) returns ParGenCurve;

Value(me; U : Real)returns Pnt2d;
    --- Purpose : Computes the point of parameter U on the curve 

D1 (me; U : Real; P : out Pnt2d from gp ; V : out Vec2d from gp);
    --- Purpose : Computes the point of parameter U on the curve with its
    --  first derivative.

D2 (me; U : Real; P : out Pnt2d from gp ; V1,V2 : out Vec2d from gp);
    --- Purpose : Computes the point of parameter U on the curve with its
    --  first derivative and second derivative.


FirstParameter(me)  returns Real;
    	
LastParameter(me) returns Real;

GetResolution(me) returns Real;

GetIntervals(me) returns Integer;

fields

Cu  : TheCurve              ;
Dep : Real     from Standard;

end ParGenCurve;
