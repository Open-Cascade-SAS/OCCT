-- Created on: 2000-07-03
-- Created by: Andrey BETENEV
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1

class QuantifiedAssemblyComponentUsage from StepRepr
inherits AssemblyComponentUsage from StepRepr

    ---Purpose: Representation of STEP entity QuantifiedAssemblyComponentUsage

uses
    HAsciiString from TCollection,
    ProductDefinition from StepBasic,
    MeasureWithUnit from StepBasic

is
    Create returns QuantifiedAssemblyComponentUsage from StepRepr;
	---Purpose: Empty constructor

    Init (me: mutable; aProductDefinitionRelationship_Id: HAsciiString from TCollection;
                       aProductDefinitionRelationship_Name: HAsciiString from TCollection;
                       hasProductDefinitionRelationship_Description: Boolean;
                       aProductDefinitionRelationship_Description: HAsciiString from TCollection;
                       aProductDefinitionRelationship_RelatingProductDefinition: ProductDefinition from StepBasic;
                       aProductDefinitionRelationship_RelatedProductDefinition: ProductDefinition from StepBasic;
                       hasAssemblyComponentUsage_ReferenceDesignator: Boolean;
                       aAssemblyComponentUsage_ReferenceDesignator: HAsciiString from TCollection;
                       aQuantity: MeasureWithUnit from StepBasic);
	---Purpose: Initialize all fields (own and inherited)

    Quantity (me) returns MeasureWithUnit from StepBasic;
	---Purpose: Returns field Quantity
    SetQuantity (me: mutable; Quantity: MeasureWithUnit from StepBasic);
	---Purpose: Set field Quantity

fields
    theQuantity: MeasureWithUnit from StepBasic;

end QuantifiedAssemblyComponentUsage;
