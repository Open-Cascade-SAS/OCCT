-- Created by: Peter KURNEV
-- Copyright (c) 2010-2014 OPEN CASCADE SAS
-- Copyright (c) 2007-2010 CEA/DEN, EDF R&D, OPEN CASCADE
-- Copyright (c) 2003-2007 OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN, CEDRAT,
--                         EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class BuilderArea from BOPAlgo 
    	inherits Algo from BOPAlgo 
	 
	---Purpose: The root class for algorithms to build  
    	--          faces/solids from set of edges/faces  

uses 
    Shape from TopoDS, 
    BaseAllocator from BOPCol, 
    ListOfShape from BOPCol,
    MapOfOrientedShape from BOPCol, 
    Context  from BOPInt 
    
--raises

is 
    Initialize  
    	returns BuilderArea from BOPAlgo; 
    ---C++: alias "Standard_EXPORT virtual ~BOPAlgo_BuilderArea();"  
     
    Initialize(theAllocator: BaseAllocator from BOPCol)   
    	returns BuilderArea from BOPAlgo; 
     
    SetContext(me:out; 
    	    theContext:Context from BOPInt);  
    	
    Shapes(me) 
    	returns ListOfShape from BOPCol;   
    ---C++:  return const &   
    ---C++: alias "Standard_EXPORT void SetShapes(const BOPCol_ListOfShape& theLS);"  
    
    Loops(me)  
    	returns ListOfShape from BOPCol; 
    ---C++:  return const &   
     
    Areas(me) 
    	returns ListOfShape from BOPCol; 
    ---C++:  return const &     
     
    PerformShapesToAvoid(me:out) 
    	is deferred protected; 
	 
    PerformLoops(me:out) 
    	is deferred protected;  
	 
    PerformAreas(me:out)   
    	is deferred protected;  

    PerformInternalShapes(me:out)   
    	is deferred protected;  

fields  
    myContext        :  Context from BOPInt is protected; 
    myShapes         :  ListOfShape from BOPCol is protected;  
    myLoops          :  ListOfShape from BOPCol is protected;  
    myLoopsInternal  :  ListOfShape from BOPCol is protected;
    
    myAreas          :  ListOfShape from BOPCol is protected;  
    myShapesToAvoid  :  MapOfOrientedShape from BOPCol is protected;  
    --
       	 

end BuilderArea; 

