-- Created on: 2018-03-15
-- Created by: Stephan GARNAUD (ARM)
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Host from OSD

 ---Purpose: Carries information about a Host


uses SysType, OEMType, Error, AsciiString from TCollection
raises ConstructionError, NullObject, OSDError

 is

  Create returns Host;
    ---Purpose: Initializes current host by default.
    ---Level: Advanced

  SystemVersion (me : in out) returns AsciiString is static;
    ---Purpose: Returns system name and version
    ---Level: Advanced

  SystemId (me) returns SysType is static;
    ---Purpose: Returns the system type (UNIX System V, UNIX BSD, MS-DOS...)
    ---Level: Advanced

  HostName (me : in out) returns AsciiString is static;
    ---Purpose: Returns host name.
    ---Level: Advanced

  AvailableMemory (me : in out)  returns Integer is static;
    ---Purpose: Returns available memory in Kilobytes.
    ---Level: Obsolete syntax. Will be removed in next version

  InternetAddress (me : in out) returns AsciiString is static;
    ---Purpose: Returns Internet address of current host.
    ---Level: Advanced

  MachineType (me : in out) returns OEMType is static;
    ---Purpose: Returns type of current machine.
    ---Level: Advanced

 Failed (me) returns Boolean is static;
   ---Purpose: Returns TRUE if an error occurs
   ---Level: Advanced

 Reset (me : in out) is static;
   ---Purpose: Resets error counter to zero
   ---Level: Advanced
      
 Perror (me : in out)
   ---Purpose: Raises OSD_Error
   ---Level: Advanced
   raises OSDError is static;

 Error (me) returns Integer is static;
   ---Purpose: Returns error number if 'Failed' is TRUE.
   ---Level: Advanced

fields
  myName   : AsciiString;
  myError  : Error;
end Host from OSD;


