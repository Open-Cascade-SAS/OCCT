-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Axis2Placement from StepGeom inherits SelectType from StepData

	-- <Axis2Placement> is an EXPRESS Select Type construct translation.
	-- it gathers : Axis2Placement2d, Axis2Placement3d

uses

	Axis2Placement2d,
	Axis2Placement3d
is

	Create returns Axis2Placement;
	---Purpose : Returns a Axis2Placement SelectType

	CaseNum (me; ent : Transient) returns Integer;
	---Purpose: Recognizes a Axis2Placement Kind Entity that is :
	--        1 -> Axis2Placement2d
	--        2 -> Axis2Placement3d
	--        0 else

	Axis2Placement2d (me) returns any Axis2Placement2d;
	---Purpose : returns Value as a Axis2Placement2d (Null if another type)

	Axis2Placement3d (me) returns any Axis2Placement3d;
	---Purpose : returns Value as a Axis2Placement3d (Null if another type)


end Axis2Placement;

