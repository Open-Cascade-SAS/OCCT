-- Created on: 1997-03-26
-- Created by: Christian CAILLET
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ApprovalDateTime  from StepBasic    inherits TShared

    ---Purpose : Added from StepBasic Rev2 to Rev4

uses
    DateTimeSelect from StepBasic,
    Approval from StepBasic

is

    Create returns ApprovalDateTime;

    Init (me : mutable;
    	  aDateTime : DateTimeSelect;
	  aDatedApproval : Approval);

    SetDateTime (me : mutable; aDateTime : DateTimeSelect);
    DateTime    (me) returns DateTimeSelect;

    SetDatedApproval (me : mutable; aDatedApproval : Approval);
    DatedApproval    (me) returns Approval;

fields

    theDateTime : DateTimeSelect;
    theDatedApproval : Approval;

end ApprovalDateTime;
