-- File:        TypeQualifier.cdl
-- Created:     Mon Dec  4 12:02:23 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWTypeQualifier from RWStepShape

	---Purpose : Read & Write Module for TypeQualifier

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     TypeQualifier from StepShape

is

	Create returns RWTypeQualifier;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable TypeQualifier from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : TypeQualifier from StepShape);

end RWTypeQualifier;
