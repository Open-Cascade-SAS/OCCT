-- Created on: 1997-05-09
-- Created by: Christian CAILLET
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ECDescr  from StepData    inherits EDescr  from StepData

    ---Purpose : Describes a Complex Entity (Plex) as a list of Simple ones

uses HSequenceOfAsciiString from TColStd, SequenceOfTransient from TColStd,
     ESDescr from StepData, Described from StepData

is

    Create returns ECDescr;
    ---Purpose : Creates an ECDescr, empty

    Add (me : mutable; member : ESDescr);
    ---Purpose : Adds a member
    --  Warning : members are added in alphabetic order

    NbMembers (me) returns Integer;
    ---Purpose : Returns the count of members

    Member (me; num : Integer) returns ESDescr;
    ---Purpose : Returns a Member from its rank

    TypeList (me) returns HSequenceOfAsciiString;
    ---Purpose : Returns the ordered list of types


    	--  inherited

    Matches    (me; steptype : CString) returns Boolean;
    ---Purpose : Tells if a ESDescr matches a step type : exact or super type

    IsComplex  (me) returns Boolean;
    ---Purpose : Returns True

    NewEntity  (me) returns Described;
    ---Purpose : Creates a described entity (i.e. a complex one, made of one
    --           simple entity per member)

fields

    thelist : SequenceOfTransient;

end ECDescr;
