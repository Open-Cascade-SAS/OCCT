-- Created on: 2008-04-17
-- Created by: Customer Support
-- Copyright (c) 2008-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class LayerMgr from V3d inherits TShared from MMgt

    ---Purpose: Class to manage layers

uses

    ExtendedString from TCollection,
    Color from Quantity,
    Layer from Visual3d,
    ColorScale from Aspect,
    ColorScale from V3d,
    ColorScaleLayerItem from V3d,
    View from V3d,
    ViewPointer from V3d
    

is

    ---Category: Public

    Create (aView : View from V3d)
    returns mutable LayerMgr from V3d;
    
    Overlay (me)
    returns mutable Layer from Visual3d;
    ---C++: return const &
    ---C++: inline

    View (me)
    returns mutable View from V3d;
    ---C++: inline

    ColorScaleDisplay (me : mutable);
    ColorScaleErase (me : mutable);
    ColorScaleIsDisplayed (me) returns Boolean from Standard;
    ColorScale (me) returns mutable ColorScale from Aspect;

    Compute (me : mutable);
    ---Purpose: Recompute layer with objects

    Resized(me : mutable);

    ---Category: Protected

    Begin (me : mutable) returns Boolean from Standard is virtual protected;
    ---Purpose: Begin layers recomputation

    Redraw (me : mutable) is virtual protected;
    ---Purpose: Perform layers recomputation

    End (me : mutable) is virtual protected;
    ---Purpose: End layers recomputation

fields

    myView       : ViewPointer from V3d is protected;
    myOverlay    : Layer from Visual3d is protected;
    myColorScale : ColorScale from V3d is protected;
    
    myColorScaleLayerItem: ColorScaleLayerItem from V3d is protected;

end LayerMgr;
