-- File:	IGESDraw_ToolSegmentedViewsVisible.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolSegmentedViewsVisible  from IGESDraw

    ---Purpose : Tool to work on a SegmentedViewsVisible. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses SegmentedViewsVisible from IGESDraw,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolSegmentedViewsVisible;
    ---Purpose : Returns a ToolSegmentedViewsVisible, ready to work


    ReadOwnParams (me; ent : mutable SegmentedViewsVisible;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : SegmentedViewsVisible;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : SegmentedViewsVisible;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a SegmentedViewsVisible <ent>, from
    --           its specific (own) parameters

    DirChecker (me; ent : SegmentedViewsVisible) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : SegmentedViewsVisible;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : SegmentedViewsVisible; entto : mutable SegmentedViewsVisible;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : SegmentedViewsVisible;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolSegmentedViewsVisible;
