-- Created on: 1993-07-23
-- Created by: Jean Louis FRENKEL
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class ColorPixel from Aspect inherits Pixel from Aspect

uses
    Color   from Quantity
is

    Create returns ColorPixel from Aspect;
	---Level: Public

    Create(aColor: Color from Quantity) returns ColorPixel from Aspect;
	---Level: Public

    Value (me) returns Color from Quantity is static ;
	---Level: Public
	   ---C++: return const &

    SetValue(me: in out; aColor: Color from Quantity) is static ;
	---Level: Public

    Print( me ; s : in out OStream from Standard ) is redefined static ;
	---Level: Public
	---Purpose : Prints the contents of <me> on the stream <s>

    HashCode (me; Upper : Integer ) returns Integer is redefined static ;
	---Level: Public
	---Purpose: Returns a hashed value denoting <me>. This value is in
	--         the range 1..<Upper>.
	---C++:  function call

    	IsEqual(me; Other : ColorPixel from Aspect) returns Boolean;
	    ---C++: alias operator==

    	IsNotEqual(me; Other : ColorPixel from Aspect) returns Boolean;
           ---C++: alias operator!=



fields
    myColor: Color from Quantity;

end ColorPixel from Aspect;
