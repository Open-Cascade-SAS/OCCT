-- Created on: 1997-05-27
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Modified by skv - Mon May 31 12:26:27 2004 OCC5865


private class BuildWires from LocOpe 

	---Purpose: 

-- Modified by skv - Mon May 31 12:53:04 2004 OCC5865 Begin
uses ListOfShape from TopTools,
     ProjectedWires from LocOpe
-- Modified by skv - Mon May 31 12:53:05 2004 OCC5865 End

raises NotDone from StdFail

is

    Create
    
    	returns BuildWires from LocOpe;


-- Modified by skv - Mon May 31 12:54:10 2004 OCC5865 Begin
    Create(Ledges: ListOfShape from TopTools;
    	   PW    : ProjectedWires  from  LocOpe)
-- Modified by skv - Mon May 31 12:54:11 2004 OCC5865 End
    
    	returns BuildWires from LocOpe;


-- Modified by skv - Mon May 31 12:54:10 2004 OCC5865 Begin
    Perform(me: in out; Ledges: ListOfShape from TopTools; 
    	    	        PW    : ProjectedWires  from  LocOpe)
-- Modified by skv - Mon May 31 12:54:11 2004 OCC5865 End
    
    	is static;


    IsDone(me)
    
    	returns Boolean from Standard
	is static;


    Result(me)
    
    	returns ListOfShape from TopTools
	---C++: return const&
    	raises NotDone from StdFail
	is static;



fields

    myDone : Boolean from Standard;
    myRes  : ListOfShape from TopTools;

end BuildWires;
