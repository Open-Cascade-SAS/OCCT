-- File:	IGESSelect_CounterOfLevelNumber.cdl
-- Created:	Tue May 31 14:32:15 1994
-- Author:	Modelistation
--		<model@bravox>
---Copyright:	 Matra Datavision 1994


class CounterOfLevelNumber  from IGESSelect  inherits SignCounter

    ---Purpose : This class gives information about Level Number. It counts
    --           entities according level number, considering also the
    --           multiple level (see the class LevelList) for which an entity
    --           is attached to each of the listed levels.
    --           
    --           Data are available, as level number, or as their alphanumeric
    --           counterparts ("LEVEL nnnnnnn", " NO LEVEL", " LEVEL LIST")

uses Integer, Transient, MapOfTransient, HAsciiString from TCollection,
     HArray1OfInteger from TColStd, HSequenceOfInteger from TColStd,
     Messenger from Message,
     HSequenceOfTransient, InterfaceModel

is

    Create (withmap  : Boolean = Standard_True;
    	    withlist : Boolean = Standard_False)
    	 returns mutable CounterOfLevelNumber;
    ---Purpose : Creates a CounterOfLevelNumber, clear, ready to work
    --           <withmap> and <withlist> are transmitted to SignCounter

    Clear (me : mutable) is redefined;
    ---Purpose : Resets already memorized informations : also numeric data

    AddSign  (me : mutable; ent : Transient; model : InterfaceModel)
    	is redefined;
    ---Purpose : Adds an entity by considering its lrvrl number(s)
    --	         A level is added both in numeric and alphanumeric form,
    --           i.e. LevelList gives "LEVEL LIST", others (no level or
    --           positive level) displays level number on 7 digits (C : %7d)
    --           Remark : an entity attached to a Level List is added for
    --           " LEVEL LIST", and for each of its constituant levels

    AddLevel (me : mutable; ent : Transient; level : Integer);
    ---Purpose : The internal action to record a new level number, positive,
    --           null (no level) or negative (level list)

    HighestLevel (me) returns Integer;
    ---Purpose : Returns the highest value found for a level number

    NbTimesLevel (me; level : Integer) returns Integer;
    ---Purpose : Returns the number of times a level is used,
    --           0 if it has not been recorded at all
    --           <level> = 0 counts entities attached to no level
    --           <level> < 0 counts entities attached to a LevelList

    Levels (me) returns HSequenceOfInteger;
    ---Purpose : Returns the ordered list of used positive Level numbers

    Sign (me; ent : Transient; model : InterfaceModel) returns HAsciiString  is redefined;
    ---Purpose : Determines and returns the value of the signature for an
    --           entity as an HAsciiString. Redefined, gives the same result
    --           as AddSign, see this method ("LEVEL LIST" or "nnnnnnn")

    PrintCount (me; S : Messenger from Message)  is redefined;
    ---Purpose : Prints the counts of items (not the list) then the Highest
    --           Level Number recorded

fields

    thehigh    : Integer;
    thenblists : Integer;
    thelevels  : HArray1OfInteger;

end CounterOfLevelNumber;
