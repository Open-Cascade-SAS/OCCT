-- Created by: Peter KURNEV
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Curve from BOPDS 

	---Purpose:  
    	-- The class BOPDS_Curve is to store  
    	-- the information about intersection curve 

uses 
    Box from Bnd,
    Curve from IntTools, 
    ListOfInteger from BOPCol, 
    BaseAllocator from BOPCol, 
    ListOfPaveBlock from BOPDS, 
    PaveBlock from BOPDS 
    
--raises

is 
    Create 
    	returns Curve from BOPDS;  
    ---C++: alias "virtual ~BOPDS_Curve();" 
    ---C++: inline  
	---Purpose:  
    	--- Empty contructor  
    	--- 
    Create (theAllocator: BaseAllocator from BOPCol) 
    	returns Curve from BOPDS;      
    ---C++: inline   
     	---Purpose:  
    	---  Contructor    
    	---  <theAllocator> - the allocator to manage the memory     
    	---  
	
    SetCurve(me:out; 
    	     theC:Curve from IntTools);  
    ---C++: inline  
    	---Purpose: 
    	--- Modifier   
	--- Sets the curve <theC> 
	 
    Curve(me)
    	returns Curve from IntTools; 
    ---C++: return const &  
    ---C++: inline 
      	---Purpose: 
    	--- Selector   
	--- Returns the curve  
	 
    SetBox(me:out; 
    	    theBox:Box from Bnd); 
    ---C++: inline 
     	---Purpose: 
    	--- Modifier   
	--- Sets the bounding box <theBox> of the curve 
	 
    Box(me) 
    	returns Box from Bnd; 
    ---C++: return const &    
    ---C++: inline 
     	---Purpose: 
    	--- Selector   
	--- Returns the bounding box of the curve 
	 
    ChangeBox(me:out) 
    	returns Box from Bnd; 
    ---C++: return  &    
    ---C++: inline  
    	---Purpose: 
    	--- Selector/Modifier  
	--- Returns the bounding box of the curve 
    SetPaveBlocks(me:out; 
    	    theLPB:ListOfPaveBlock from BOPDS); 
	     
    PaveBlocks (me) 
        returns ListOfPaveBlock from BOPDS;  
    ---C++: return const &   
    ---C++: inline       
     	---Purpose: 
    	--- Selector   
	--- Returns the list of pave blocks  
    	--- of the curve 
	 
    ChangePaveBlocks (me:out) 
        returns ListOfPaveBlock from BOPDS; 
    ---C++: return & 
    ---C++: inline      
      	---Purpose: 
    	--- Selector/Modifier   
	--- Returns the list of pave blocks   
	--- of the curve  
	
    InitPaveBlock1(me:out); 
    ---C++: inline 
    	---Purpose: 
	--- Creates  initial pave block   
	--- of the curve   
	
    ChangePaveBlock1(me:out) 
    	returns PaveBlock from BOPDS; 
    ---C++: return &  
    ---C++: inline  
    	---Purpose:  
	--- Selector/Modifier 
	--- Returns  initial pave block   
	--- of the curve   

    TechnoVertices (me) 
    	returns ListOfInteger from BOPCol; 
    ---C++: return const &  
    ---C++: inline      
     	---Purpose:  
	--- Selector
	--- Returns list of indices of technologic vertices   
	--- of the curve    
	
    ChangeTechnoVertices (me:out) 
    	returns ListOfInteger from BOPCol; 
    ---C++:  return & 
    ---C++: inline  
     	---Purpose:  
	--- Selector/Modifier 
	--- Returns list of indices of technologic vertices   
	--- of the curve   
	 
    HasEdge(me) 
    	returns Boolean from Standard;  
    ---C++: inline 
    	---Purpose:  
	--- Query 
	--- Returns true if at least one pave block of the curve  
    	--  has edge  
fields 
    myAllocator      : BaseAllocator from BOPCol is protected;
    myCurve          : Curve from IntTools is protected; 
    myPaveBlocks     : ListOfPaveBlock from BOPDS is protected; 
    myTechnoVertices : ListOfInteger from BOPCol is protected;  
    myBox            : Box from Bnd is protected; 

end Curve;
