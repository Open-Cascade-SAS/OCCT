-- File:        EdgeCurve.cdl
-- Created:     Mon Dec  4 12:02:26 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWEdgeCurve from RWStepShape

	---Purpose : Read & Write Module for EdgeCurve
	--           Check added by CKY , 7-OCT-1996

uses Check from Interface, ShareTool from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     EdgeCurve from StepShape,
     EntityIterator from Interface

is

	Create returns RWEdgeCurve;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable EdgeCurve from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : EdgeCurve from StepShape);

	Share(me; ent : EdgeCurve from StepShape; iter : in out EntityIterator);

	Check(me; ent : EdgeCurve from StepShape; shares : ShareTool; ach : in out Check);

end RWEdgeCurve;
