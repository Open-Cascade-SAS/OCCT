-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class AutoDesignDateAndTimeItem from StepAP214 inherits SelectType from StepData

	-- <AutoDesignDateAndTimeItem> is an EXPRESS Select Type construct translation.
	-- it gathers : ApprovalPersonOrganization, AutoDesignDateAndPersonAssignment

uses

	ApprovalPersonOrganization from StepBasic,
	AutoDesignDateAndPersonAssignment from StepAP214,
	ProductDefinitionEffectivity from StepBasic
is

	Create returns AutoDesignDateAndTimeItem;
	---Purpose : Returns a AutoDesignDateAndTimeItem SelectType

	CaseNum (me; ent : Transient) returns Integer;
	---Purpose: Recognizes a AutoDesignDateAndTimeItem Kind Entity that is :
	--        1 -> ApprovalPersonOrganization
	--        2 -> AutoDesignDateAndPersonAssignment
	--        0 else

	ApprovalPersonOrganization (me) returns any ApprovalPersonOrganization;
	---Purpose : returns Value as a ApprovalPersonOrganization (Null if another type)

	AutoDesignDateAndPersonAssignment (me) returns any AutoDesignDateAndPersonAssignment;
	---Purpose : returns Value as a AutoDesignDateAndPersonAssignment (Null if another type)

    	ProductDefinitionEffectivity (me) returns ProductDefinitionEffectivity;

end AutoDesignDateAndTimeItem;
