-- Created on: 1997-01-08
-- Created by: Robert COUBLANC
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ConnectedInteractive from AIS inherits InteractiveObject from AIS

	---Purpose: Creates an arbitrary located instance of another Interactive Object,
    	-- which serves as a reference.
    	-- This allows you to use the Connected Interactive
    	-- Object without having to recalculate presentation,
    	-- selection or graphic structure. These are deduced
    	-- from your reference object.
    	-- The relation between the connected interactive object
    	-- and its source is generally one of geometric transformation. 
        -- AIS_ConnectedInteractive class supports selection mode 0 for any InteractiveObject and
        -- all standard modes if its reference based on AIS_Shape.
        -- Descendants may redefine ComputeSelection() though.
    	-- Also ConnectedInteractive will handle HLR if its reference based on AIS_Shape.

uses
    Location              from TopLoc,
    Shape                 from TopoDS,
    Transformation        from Geom,
    PresentationManager3d from PrsMgr,
    Presentation          from Prs3d,
    TypeOfPresentation3d  from PrsMgr,
    Selection             from SelectMgr,
    Projector             from Prs3d,
    KindOfInteractive     from AIS,
    Trsf                  from gp
raises
    NotImplemented from Standard

is

    Create (aTypeOfPresentation3d: TypeOfPresentation3d from PrsMgr = PrsMgr_TOP_AllView) 
    returns  ConnectedInteractive  from  AIS;
    	---Purpose:
    	-- Disconnects the previous view and sets highlight
    	-- mode to 0. This highlights the wireframe presentation
    	-- aTypeOfPresentation3d.
    	-- Top_AllView deactivates hidden line removal.
    
    Type(me) returns KindOfInteractive from AIS 
    is redefined virtual;
  	---Purpose: Returns KOI_Object

    Signature(me) returns Integer from Standard
    is redefined virtual;
	---Purpose: Returns 1


    Connect(me          : mutable; 
    	    anotherIObj : InteractiveObject from AIS) is virtual;
    	---Purpose: Establishes the connection between the Connected
    	-- Interactive Object, anotherIobj, and its reference.


    Connect(me:mutable;
    	    anotherIobj: InteractiveObject from AIS;
	        aLocation : Trsf from gp) is virtual;
        ---Purpose: Establishes the connection between the Connected
        -- Interactive Object, anotherIobj, and its reference.
        -- Locates instance in aLocation.
	    

    HasConnection(me) returns Boolean from Standard;
        ---C++: inline
    	---Purpose:
    	-- Returns true if there is a connection established
    	-- between the presentation and its source reference.
	
    ConnectedTo(me) returns any InteractiveObject from AIS;
     	---C++: inline
	---C++: return const&
    	---Purpose:
    	-- Returns the connection with the reference Interactive Object.

	    
    Disconnect(me:mutable);
	---Purpose: Clears the connection with a source reference. The
    	-- presentation will no longer be displayed.
    	-- Warning Must be done before deleting the presentation.

    Compute(me                   : mutable;
            aPresentationManager : PresentationManager3d from PrsMgr;
            aPresentation        : Presentation from Prs3d;
            aMode                : Integer from Standard = 0)
	---Level: Public 
	---Purpose: Calculates the view aPresentation and its updates.
    	-- The latter are managed by aPresentationManager.
    	-- The display mode aMode is 0 by default.
    	--    this method is redefined virtual;
	--          when the instance is connected to another
    	--          InteractiveObject,this method doesn't
    	--          compute anything, but just uses the 
	--          presentation of this last object, with
	--          a transformation if there's one stored. 
    is redefined virtual private;

    Compute(me            : mutable;
    	    aProjector    : Projector from Prs3d;
    	    aTrsf         : Transformation from Geom;
	    aPresentation : Presentation from Prs3d)
    is redefined virtual private;
	---Purpose: Computes the presentation according to a point of view
	--          given by <aProjector>. 
	--          To be Used when the associated degenerated Presentations 
	--          have been transformed by <aTrsf> which is not a Pure
	--          Translation. The HLR Prs can't be deducted automatically
	--          WARNING :<aTrsf> must be applied
	--           to the object to display before computation  !!!


    Compute(me:mutable;
    	        aProjector: Projector from Prs3d;
                aPresentation: Presentation from Prs3d)
    is redefined virtual private;
    ---Purpose: Computes the presentation according to a point of view
    --          given by <aProjector>. 
    
    ComputeSelection(me:mutable; theSelection : Selection from SelectMgr;
                                 theMode      : Integer) is redefined virtual private;
	---Level: Public 
	---Purpose: Generates sensitive entities by copying 
        -- them from myReference selection, creates and sets an entity 
        -- owner for this entities and adds them to theSelection

    computeSubShapeSelection (me:mutable; theSelection : Selection from SelectMgr;
                                          theMode      : Integer) is private;
    ---Level: Public 
    ---Purpose: Generates sensitive entities by copying 
        -- them from myReference sub shapes selection, creates and sets an entity 
        -- owner for this entities and adds them to theSelection

    AcceptShapeDecomposition(me) returns Boolean from Standard is 
    redefined virtual;
        ---C++: inline
        ---Purpose:  Informs the graphic context that the interactive Object
        -- may be decomposed into sub-shapes for dynamic selection.


    updateShape(me:mutable;WithLocation:Boolean from Standard = Standard_True)
    is static private;
    
    Compute(me:mutable;
                aProjector   :         Projector    from Prs3d;
                aPresentation: Presentation from Prs3d;
                aShape       :         Shape from TopoDS)
    is  private;
    ---Purpose: Computes the presentation according to a point of view
    --          given by <aProjector>. 
    
fields

    myReference : InteractiveObject from AIS is protected; -- reference object
    myShape : Shape from TopoDS; -- used for HLR

end ConnectedInteractive;


