-- File:        UncertaintyMeasureWithUnit.cdl
-- Created:     Mon Dec  4 12:02:32 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWUncertaintyMeasureWithUnit from RWStepBasic

	---Purpose : Read & Write Module for UncertaintyMeasureWithUnit

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     UncertaintyMeasureWithUnit from StepBasic,
     EntityIterator from Interface

is

	Create returns RWUncertaintyMeasureWithUnit;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable UncertaintyMeasureWithUnit from StepBasic);

	WriteStep (me; SW : in out StepWriter; ent : UncertaintyMeasureWithUnit from StepBasic);

	Share(me; ent : UncertaintyMeasureWithUnit from StepBasic; iter : in out EntityIterator);

end RWUncertaintyMeasureWithUnit;
