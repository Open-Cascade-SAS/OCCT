-- Created on: 1999-09-21
-- Created by: Edward AGAPOV
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ExtPRevS from Extrema inherits Transient from Standard
		    
	---Purpose: It calculates all the extremum (minimum and
	--          maximum) distances between a point and a surface
	--          of revolution.
		    
uses
    POnSurf from Extrema,
    GenExtPS from Extrema,

    HSurfaceOfRevolution from Adaptor3d,

    Ax2 from gp,
    Pnt from gp

raises 
    NotDone from StdFail,
    OutOfRange


is

    Create returns ExtPRevS from Extrema;

    Create (P: Pnt; S: HSurfaceOfRevolution from Adaptor3d;
		    Umin, Usup, Vmin, Vsup: Real; 
		    TolU,TolV: Real) 
		    returns ExtPRevS from Extrema;
    ---Purpose: It calculates all the distances between a point 
    --          from gp and a SurfacePtr from Adaptor3d.
    
    Create (P: Pnt; S: HSurfaceOfRevolution from Adaptor3d; 
		    TolU,TolV: Real) 
		    returns ExtPRevS from Extrema;
    ---Purpose: It calculates all the distances between a point 
    --          from gp and a SurfacePtr from Adaptor3d.
    
    Initialize(me: mutable; S: HSurfaceOfRevolution from Adaptor3d; 
			   Umin, Usup, Vmin, Vsup: Real; 
			   TolU,TolV: Real)
		    is static;
    
    Perform (me: mutable; P: Pnt)
		    is static;
    
    IsDone (me) returns Boolean
    ---Purpose: Returns True if the distances are found.
    		    is static;
    
    NbExt (me) returns Integer
    ---Purpose: Returns the number of extremum distances.
    		    raises  NotDone from StdFail
	    	-- if IsDone(me)=False.
    		    is static;

    SquareDistance (me; N: Integer) returns Real
    ---Purpose: Returns the value of the Nth resulting square distance.
    		    raises  NotDone from StdFail,
    	    	-- if IsDone(me)=False.
    	        OutOfRange
		-- if N < 1 or N > NbPoints(me).
    		    is static;

    Point (me; N: Integer) returns POnSurf
    ---C++: return const &
    ---Purpose: Returns the point of the Nth resulting distance.
    		    raises  NotDone from StdFail,
    	    	-- if IsDone(me)=False.
    	        OutOfRange
		-- if N < 1 or N > NbPoints(me).
    		    is static;

fields
    myS      : HSurfaceOfRevolution from Adaptor3d;
    myvinf   : Real                 from Standard;
    myvsup   : Real                 from Standard;
    mytolv   : Real                 from Standard;
    
    myPosition  : Ax2      from gp;
    myExtPS     : GenExtPS from Extrema;
    
    myIsAnalyticallyComputable : Boolean  from Standard;

    myDone : Boolean;
    myNbExt: Integer;
    mySqDist: Real [8];
    myPoint: POnSurf from Extrema [8];

end ExtPRevS;
