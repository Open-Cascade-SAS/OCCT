-- File:	IGESSolid_ToolSolidOfLinearExtrusion.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolSolidOfLinearExtrusion  from IGESSolid

    ---Purpose : Tool to work on a SolidOfLinearExtrusion. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses SolidOfLinearExtrusion from IGESSolid,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolSolidOfLinearExtrusion;
    ---Purpose : Returns a ToolSolidOfLinearExtrusion, ready to work


    ReadOwnParams (me; ent : mutable SolidOfLinearExtrusion;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : SolidOfLinearExtrusion;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : SolidOfLinearExtrusion;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a SolidOfLinearExtrusion <ent>, from
    --           its specific (own) parameters

    DirChecker (me; ent : SolidOfLinearExtrusion) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : SolidOfLinearExtrusion;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : SolidOfLinearExtrusion; entto : mutable SolidOfLinearExtrusion;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : SolidOfLinearExtrusion;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolSolidOfLinearExtrusion;
