-- Created on: 1994-02-18
-- Created by: Remi LEQUETTE
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- modified by Michael KLOKOV  Wed Mar  6 15:01:25 2002

class Section from BRepAlgoAPI inherits BooleanOperation from BRepAlgoAPI

    	---Purpose: Computes the intersection of two shapes or geometries.
    	-- Geometries can be surfaces of planes.
    	-- Geometries are converted to faces
    	-- When a geometry has been converted to
    	-- topology the created shape can be found using
    	-- the methods Shape1 and Shape2 inherited from the class BooleanOperation.
    	-- The result (Shape() method) is a compound containing 
    	-- edges built on intersection curves.
    	-- By default, the section is performed immediatly in 
    	-- class constructors, with default values :
    	-- - geometries built are NOT approximated.
    	-- - PCurves are NOT computed on both parts.
    	-- Example : giving two shapes S1,S2 accessing faces,
    	-- let compute the section edges R on S1,S2, 
    	-- performing approximation on new curves,
    	-- performing PCurve on part 1 but not on part 2 :
    	-- Standard_Boolean PerformNow = Standard_False;
    	-- BRepBoolAPI_Section S(S1,S2,PerformNow);
    	-- S.ComputePCurveOn1(Standard_True);
    	-- S.Approximation(Standard_True);
    	-- S.Build();
    	-- TopoDS_Shape R = S.Shape();
    	-- On Null Shapes of geometries, NotDone() is called. 

uses
    Pln   from gp,
    Shape from TopoDS,
    Surface from Geom,
    Curve   from Geom2d,
    DSFiller from BOPTools,
    ListOfShape from TopTools
    
is
        Create (S1,S2 : Shape from TopoDS; 
    	    aDSF:DSFiller from BOPTools;
    	    PerformNow : Boolean = Standard_True)  
    	returns Section from BRepAlgoAPI;

    Create(Sh1,Sh2 : Shape from TopoDS;
    	   PerformNow : Boolean = Standard_True)
    	---Purpose: see upper
    	---Level: Public
    	returns Section from BRepAlgoAPI;

    Create(Sh : Shape from TopoDS; Pl : Pln from gp;
    	   PerformNow : Boolean = Standard_True)
    	---Purpose: see upper
    	---Level: Public
    	returns Section from BRepAlgoAPI;

    Create(Sh : Shape from TopoDS; Sf : Surface from Geom;
 	   PerformNow : Boolean = Standard_True)
    	---Purpose: see upper
    	---Level: Public
    	returns Section from BRepAlgoAPI;

    Create(Sf : Surface from Geom; Sh : Shape from TopoDS;
 	   PerformNow : Boolean = Standard_True)
    	---Purpose: see upper
    	---Level: Public
	returns Section from BRepAlgoAPI;

    Create(Sf1 : Surface from Geom; Sf2 : Surface from Geom;
    	PerformNow : Boolean = Standard_True)
    	---Purpose: This and the above classes construct a framework for
    	-- computing the section lines of:
    	-- -       two shapes Sh1 and Sh2, or
    	-- -       shape Sh and plane Pl,  or
    	-- -       shape Sh and surface Sf, or
    	-- -       surface Sf and shape Sh, or
    	-- -       two surfaces Sf1 and Sf2,
    	--   and builds a result if PerformNow equals true, its
    	-- default value. If PerformNow equals false, the intersection
    	-- will be computed later by the function Build.
    	--  The constructed shape will be returned by the function Shape.
    	-- This is a compound object composed of edges. These
    	-- intersection edges may be built:
    	-- -      on new intersection lines, or
    	-- -      on coincident portions of edges in the two intersected    shapes.
    	--   These intersection edges are independent: they are not
    	-- chained or grouped in wires. If no intersection edge exists, the
    	-- result is an empty compound object.
    	-- Note that other objects than TopoDS_Shape shapes involved in
    	-- these syntaxes are converted into faces or shells before
    	-- performing the computation of the intersection. A shape
    	-- resulting from this conversion can be retrieved with the
    	-- function Shape1 or Shape2.
    	-- Parametric 2D curves on intersection edges
    	-- No parametric 2D curve (pcurve) is defined for each elementary
    	-- edge of the result. To attach such parametric curves to the
    	-- constructed edges you may use a constructor with the PerformNow
    	-- flag equal to false; then you use:
    	-- -      the function ComputePCurveOn1 to ask for
    	--    the additional computation of a pcurve in the parametric
    	--    space of the first shape,
    	-- -      the function ComputePCurveOn2 to ask for
    	--    the additional computation of a pcurve in the parametric
    	--    space of the second shape, in the end,
    	-- -      the function Build to construct the result.
    	--   Approximation of intersection edges
    	--   The underlying 3D geometry attached to each elementary edge
    	-- of the result is:
    	-- -       analytic where possible, provided the corresponding
    	--    geometry corresponds to a type of analytic curve
    	--    defined in the Geom package; for example, the intersection
    	--    of a cylindrical shape with a plane gives an ellipse or a    circle;
    	-- -       or elsewhere, given as a succession of points grouped
    	--    together in a BSpline curve of degree 1.
    	-- If you prefer to have an attached 3D geometry which is a
    	-- BSpline approximation of the computed set of points on
    	-- computed elementary intersection edges whose underlying geometry
    	-- is not analytic, you may use a constructor with the PerformNow
    	-- flag equal to false. Then you use:
    	-- -      the function Approximation to ask for this
    	--    computation option, and
    	-- -      the function Build to construct the result.
    	-- -      Note that as a result, approximations will only be
    	--    computed on edges built on new intersection lines.
    	-- -      Example
    	-- You may also combine these computation options. In the following example:
    	-- - each elementary edge of the computed intersection,
    	--   built on a new intersection line, which does not
    	--  correspond to an analytic Geom curve, will be approximated by
    	--   a BSpline curve whose degree is not greater than 8.
    	-- - each elementary edge built on a new intersection line, will have:
    	-- - a pcurve in the parametric space of the intersected face of shape S1,
    	-- - no pcurve in the parametric space of the intersected face of shape S2.
    	--       // TopoDS_Shape S1 = ... , S2 = ... ;
    	-- Standard_Boolean PerformNow = Standard_False;
    	-- BRepAlgoAPI_Section S ( S1, S2, PerformNow );
    	-- S.ComputePCurveOn1 (Standard_True);
    	-- S.Approximation (Standard_True);
    	-- S.Build();
    	-- TopoDS_Shape R = S.Shape();
	returns Section from BRepAlgoAPI;

    Init1(me : out;S1 : Shape from TopoDS);
    	---Purpose: initialize first part
    	---Level: Public
 
    Init1(me : out;Pl : Pln from gp);
    	---Purpose: initialize first part
    	---Level: Public
 
    Init1(me : out;Sf : Surface from Geom);
    	---Purpose: initialize first part
    	---Level: Public
 
    Init2(me : out;S2 : Shape from TopoDS);
    	---Purpose: initialize second part
    	---Level: Public
 
    Init2(me : out;Pl : Pln from gp);
    	---Purpose: initialize second part
    	---Level: Public
 
    Init2(me : out;Sf : Surface from Geom);
    	---Purpose: Reinitializes the first and the
    	-- second parts on which this algorithm is going to perform
    	-- the intersection computation. This is done with either: the
    	-- surface Sf, the plane Pl or the shape Sh.
    	-- You use the function Build to construct the result.
 
    Approximation(me : out;B : Boolean);
    	---Level: Public
    	---Purpose: Defines an option for computation
    	-- of further intersections. This computation will be performed by
    	-- the function Build in this framework.
    	-- By default, the underlying 3D geometry attached to each
    	-- elementary edge of the result of a computed intersection is:
    	-- - analytic where possible, provided the corresponding
    	--    geometry corresponds to a type of analytic curve defined in
    	--    the Geom package; for example the intersection of a
    	--    cylindrical shape with a plane gives an ellipse or a circle;
    	-- -      or elsewhere, given as a succession of points grouped
    	-- together in a BSpline curve of degree 1. If Approx equals
    	-- true, when further computations are performed in this framework
    	-- with the function Build, these edges will have an attached 3D
    	--    geometry which is a BSpline approximation of the computed
    	--    set of points.
    	--   Note that as a result, approximations will be computed
    	-- on edges built only on new intersection lines.
 
    ComputePCurveOn1(me : out;B : Boolean);
    	---Level: Public
    	---Purpose: 
    	-- Indicates if the Pcurve must be (or not) performed on first part. 

    ComputePCurveOn2(me : out;B : Boolean);
    	---Level: Public
    	---Purpose: Define options for the computation of further
    	-- intersections, which will be performed by the function Build
    	-- in this framework.
    	-- By default, no parametric 2D curve (pcurve) is defined for the
    	-- elementary edges of the result. If ComputePCurve1 equals true,
    	-- further computations performed in this framework with the function
    	-- Build will attach an additional pcurve in the parametric space of
    	-- the first shape to the constructed edges.
    	-- If ComputePCurve2 equals true, the additional pcurve will be
    	-- attached to the constructed edges in the parametric space of the
    	-- second shape.
    	-- These two functions may be used together.
 
    Build(me : in out)
    	---Purpose:  Performs the computation of
    	-- section lines between two parts defined at the time of
    	-- construction of this framework or reinitialized with the Init1 and
    	-- Init2 functions.
    	-- The constructed shape will be returned by the function Shape.
    	-- This is a compound object composed of edges. These
    	-- intersection edges may be built:
    	-- -      on new intersection lines, or
    	-- -      on coincident portions of edges in the two intersected shapes.
    	-- These intersection edges are independent: they are not chained
    	-- or grouped into wires.
    	-- If no intersection edge exists, the result is an empty compound object.
    	-- The shapes involved in the construction of section lines can
    	-- be retrieved with the function Shape1 or Shape2. Note that other
    	-- objects than TopoDS_Shape shapes given as arguments at the
    	-- construction time of this framework, or to the Init1 or
    	-- Init2 function, are converted into faces or shells before
    	-- performing the computation of the intersection.
    	-- Parametric 2D curves on intersection edges
    	-- No parametric 2D curve (pcurve) is defined for the elementary
    	-- edges of the result. To attach parametric curves like this to
    	-- the constructed edges you have to use:
    	-- -      the function
    	-- ComputePCurveOn1 to ask for the additional computation of a
    	-- pcurve in the parametric space of the first shape,
    	-- -      the function
    	--    ComputePCurveOn2 to ask for the additional computation of a
    	--    pcurve in the parametric space of the second shape.
    	-- This must be done before calling this function.
    	--   Approximation of intersection edges
    	-- The underlying 3D geometry attached to each elementary edge of the result is:
    	-- -      analytic (where possible) provided the corresponding
    	-- geometry corresponds to a type of analytic curve defined in
    	--    the Geom package; for example, the intersection of a
    	--    cylindrical shape with a plane gives an ellipse or a circle;    or
    	-- -      elsewhere, given as a succession of points grouped
    	--    together in a BSpline curve of degree 1.
    	--   If, on computed elementary intersection edges whose
    	-- underlying geometry is not analytic, you prefer to have an
    	-- attached 3D geometry which is a Bspline approximation of the
    	-- computed set of points, you have to use the function Approximation
    	-- to ask for this computation option before calling this function.
    	-- You may also have combined these computation options: look at the
    	-- example given above to illustrate the use of the constructors.
    	is redefined static;

    HasAncestorFaceOn1(me; E : Shape from TopoDS;
    	    	    	   F : out Shape from TopoDS)
    	returns Boolean;
    	---Level: Public
    	---Purpose:
    	-- get the face of the first part giving section edge <E>.
    	-- Returns True on the 3 following conditions :
    	-- 1/ <E> is an edge returned by the Shape() method. 
    	-- 2/ First part of section performed is a shape.
    	-- 3/ <E> is built on a intersection curve (i.e <E>
    	-- 	 is not the result of common edges)
    	-- When False, F remains untouched.

    HasAncestorFaceOn2(me; E : Shape from TopoDS;
 	    	    	   F : out Shape from TopoDS)
    	returns Boolean;
    	---Purpose:  Identifies the ancestor faces of
    	-- the intersection edge E resulting from the last
    	-- computation performed in this framework, that is, the faces of
    	-- the two original shapes on which the edge E lies:
    	-- -      HasAncestorFaceOn1 gives the ancestor face in the first shape, and
    	-- -      HasAncestorFaceOn2 gives the ancestor face in the second shape.
    	--   These functions return true if an ancestor face F is found, or false if not.
    	--   An ancestor face is identifiable for the edge E if the following
    	-- conditions are satisfied:
    	-- -  the first part on which this algorithm performed its
    	--    last computation is a shape, that is, it was not given as
    	-- a surface or a plane at the time of construction of this
    	-- algorithm or at a later time by the Init1 function,
    	-- - E is one of the elementary edges built by the
    	-- last computation of this section algorithm.
    	-- To use these functions properly, you have to test the returned
    	-- Boolean value before using the ancestor face: F is significant
    	-- only if the returned Boolean value equals true.

    PCurveOn1(me; E : Shape from TopoDS)
    	returns Curve from Geom2d;
    	---Level: Public
    	---Purpose: returns the PCurve connected to section edge <E>
    	-- and lying on first part of Section.
    	-- N.B : PCurve on first part is computed only if Section is performed
    	-- after setting ComputePCurveOn1(Standard_True).

    PCurveOn2(me; E : Shape from TopoDS)
    	returns Curve from Geom2d;
    	---Level: Public
    	---Purpose: returns the PCurve connected to section edge <E>
    	-- and lying on second part of Section.
    	-- N.B : PCurve on second part is computed only if Section is performed
    	-- after setting ComputePCurveOn2(Standard_True).
    	-- Warning No pcurve is attached to an elementary edge of the
    	--    resulting section, and the function returns a null
    	--    handle, unless the function ComputePCurveOn1 or
    	--    ComputePCurveOn2 was previously used to define
    	--    this sort of option of computation.
    	-- -      A null handle is also returned if the edge E does
    	--    not belong to the last computed intersection, that
    	--    is, if it is not one of the elementary edges of the
    	--    compound object returned by the function Shape.
        
    InitParameters(me: out)
    	---Level: Private
    	is private;

fields
    myshapeisnull       : Boolean from Standard;
    myparameterschanged : Boolean from Standard;
    myApprox            : Boolean from Standard;
    myComputePCurve1    : Boolean from Standard;
    myComputePCurve2    : Boolean from Standard;
    
end Section from BRepAlgoAPI;
