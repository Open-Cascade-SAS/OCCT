-- Created on: 1997-12-03
-- Created by: Yves FRICAUD
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

private class DeltaOnModification from TNaming inherits DeltaOnModification from TDF

	---Purpose: This class provides default services for an
	--          AttributeDelta on a MODIFICATION action.
	--          
	--          Applying this AttributeDelta means GOING BACK to
	--          the attribute previously registered state.

uses

    Attribute      from TDF,
    HArray1OfShape from TopTools,
    NamedShape     from TNaming

is

    Create (NS : NamedShape from TNaming)
    	returns mutable DeltaOnModification from TNaming;
	---Purpose: Initializes a TDF_DeltaOnModification.

    Apply (me : mutable)
    	is redefined virtual;
    	---Purpose: Applies the delta to the attribute.

fields
    
    myOld  : HArray1OfShape from TopTools;
    myNew  : HArray1OfShape from TopTools;

end DeltaOnModification;
