-- Created on: 1993-01-08
-- Created by: Philippe DAUTRY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



package Sweep

    ---Purpose: This package contains generic classes usefull to create
    --          swept 3D primitives.

uses

    Standard, 
    TCollection, 
    TColStd,
    TopAbs

is

    deferred generic class Tool;
    -- signature  class. Required by  the LinearRegularSweep, defining
    -- the indexation type analysis services uppon shapes.
    
    deferred generic class Iterator;
    -- signature  class. Required by  the LinearRegularSweep, defining
    -- the iteration services uppon shapes.
    
    deferred generic class Builder;
    -- signature class. Required by the LinearRegularSweep.
    
    deferred generic class LinearRegularSweep,
    	Array2OfShapes,
        SequenceOfShapes;
	
	
    --
    --     The following classes provides a directing topology for the
    --     LinearRegularSweep. This  is  the  topology of an  open  or
    --     closed loop of edges.
    --     

    class NumShape;
	---Purpose: A shape represented by an index.
    
    class NumShapeTool;
	---Purpose: Tool for NumShapes.
    
    class NumShapeIterator;
	---Purpose: Iterator for NumShapes.
    
end Sweep;


