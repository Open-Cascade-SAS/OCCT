-- File:	RWStepAP203_RWChangeRequest.cdl
-- Created:	Fri Nov 26 16:26:35 1999 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0
-- Copyright:	Matra Datavision 1999

class RWChangeRequest from RWStepAP203

    ---Purpose: Read & Write tool for ChangeRequest

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    ChangeRequest from StepAP203

is
    Create returns RWChangeRequest from RWStepAP203;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : ChangeRequest from StepAP203);
	---Purpose: Reads ChangeRequest

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: ChangeRequest from StepAP203);
	---Purpose: Writes ChangeRequest

    Share (me; ent : ChangeRequest from StepAP203;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWChangeRequest;
