-- File:	PGeom_ToroidalSurface.cdl
-- Created:	Tue Mar  2 10:54:42 1993
-- Author:	Philippe DAUTRY
--		<fid@phylox>
-- Copyright:	 Matra Datavision 1993


class ToroidalSurface from PGeom inherits ElementarySurface from PGeom

        ---Purpose : This class defines the complete toroidal surface.
        --
	---See Also : ToroidalSurface from Geom.


uses Ax3          from gp

is



  Create returns mutable ToroidalSurface from PGeom;
	---Purpose: Creates a ToroidalSurface with default values.
    	---Level: Internal 


  Create (aPosition : Ax3 from gp;
    	  aMajorRadius: Real from Standard;
    	  aMinorRadius: Real from Standard)
     returns mutable ToroidalSurface from PGeom;
	---Purpose: Creates a ToroidalSurface with these values.
    	---Level: Internal 


  MajorRadius (me: mutable; aMajorRadius: Real from Standard);
        ---Purpose : Set the field majorRadius with <aMajorRadius>.
    	---Level: Internal 


  MajorRadius (me) returns Real from Standard;
        ---Purpose : Returns the value of the field majorRadius.
    	---Level: Internal 
     
     
  MinorRadius (me: mutable; aMinorRadius: Real from Standard);
        ---Purpose : Set the field minorRadius with <aMinorRadius>.
    	---Level: Internal 


  MinorRadius (me) returns Real from Standard;
        ---Purpose : Returns the value of the field minorRadius.
    	---Level: Internal 
     
     
fields

  majorRadius : Real from Standard;
  minorRadius : Real from Standard;

end;
