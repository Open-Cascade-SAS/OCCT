-- Created on: 1998-09-07
-- Created by: Christian CAILLET
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ActorWrite from IGESControl
    inherits ActorOfFinderProcess  from Transfer

    ---Purpose : Actor to write Shape to IGES

uses

    Finder from Transfer,
    FinderProcess from Transfer,
    Binder from Transfer

is

    Create returns ActorWrite;

    Recognize (me : mutable; start : Finder from Transfer)  returns Boolean
    	is redefined;
    ---Purpose : Recognizes a ShapeMapper

    Transfer  (me : mutable; start : Finder from Transfer;
    	       FP : mutable FinderProcess)  returns Binder  is redefined;
    ---Purpose : Transfers Shape to IGES Entities
    --         
    --           ModeTrans may be : 0 -> groups of Faces
    --           or 1 -> BRep

end ActorWrite;
