-- Created on: 2000-07-03
-- Created by: Andrey BETENEV
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1

class PropertyDefinition from StepRepr
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity PropertyDefinition

uses
    HAsciiString from TCollection,
    CharacterizedDefinition from StepRepr

is
    Create returns PropertyDefinition from StepRepr;
	---Purpose: Empty constructor

    Init (me: mutable; aName: HAsciiString from TCollection;
                       hasDescription: Boolean;
                       aDescription: HAsciiString from TCollection;
                       aDefinition: CharacterizedDefinition from StepRepr);
	---Purpose: Initialize all fields (own and inherited)

    Name (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Name
    SetName (me: mutable; Name: HAsciiString from TCollection);
	---Purpose: Set field Name

    Description (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Description
    SetDescription (me: mutable; Description: HAsciiString from TCollection);
	---Purpose: Set field Description
    HasDescription (me) returns Boolean;
	---Purpose: Returns True if optional field Description is defined

    Definition (me) returns CharacterizedDefinition from StepRepr;
	---Purpose: Returns field Definition
    SetDefinition (me: mutable; Definition: CharacterizedDefinition from StepRepr);
	---Purpose: Set field Definition

fields
    theName: HAsciiString from TCollection;
    theDescription: HAsciiString from TCollection; -- optional
    theDefinition: CharacterizedDefinition from StepRepr;
    defDescription: Boolean; -- flag "is Description defined"

end PropertyDefinition;
