-- Created on: 1993-09-28
-- Created by: Bruno DUMORTIER
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Curved from GeomFill inherits Filling from GeomFill

uses
    Array1OfPnt  from TColgp,
    Array1OfReal from TColStd

is
    Create;
    
    Create(P1, P2, P3, P4 : Array1OfPnt from TColgp)
    returns Curved from GeomFill;
    
    Create(P1, P2, P3, P4 : Array1OfPnt  from TColgp;
    	   W1, W2, W3, W4 : Array1OfReal from TColStd)
    returns Curved from GeomFill;
    

    Create(P1, P2, P3 : Array1OfPnt from TColgp)
    returns Curved from GeomFill;
    
    Create(P1, P2, P3 : Array1OfPnt  from TColgp;
    	   W1, W2, W3 : Array1OfReal from TColStd)
    returns Curved from GeomFill;
    

    Create(P1, P2 : Array1OfPnt from TColgp)
    returns Curved from GeomFill;
    
    Create(P1, P2 : Array1OfPnt  from TColgp;
    	   W1, W2 : Array1OfReal from TColStd)
    returns Curved from GeomFill;
    

    Init(me : in out;
    	 P1, P2, P3, P4 : Array1OfPnt from TColgp)
    is static;

    Init(me : in out;
    	 P1, P2, P3, P4 : Array1OfPnt  from TColgp;
    	 W1, W2, W3, W4 : Array1OfReal from TColStd)
    is static;

    Init(me : in out;
    	 P1, P2, P3 : Array1OfPnt from TColgp)
    is static;

    Init(me : in out;
    	 P1, P2, P3 : Array1OfPnt  from TColgp;
    	 W1, W2, W3 : Array1OfReal from TColStd)
    is static;

    Init(me : in out;
    	 P1, P2 : Array1OfPnt from TColgp)
    is static;

    Init(me : in out;
    	 P1, P2 : Array1OfPnt  from TColgp;
    	 W1, W2 : Array1OfReal from TColStd)
    is static;

end Curved;
