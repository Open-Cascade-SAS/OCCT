-- Created on: 1993-03-02
-- Created by: Philippe DAUTRY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



deferred class SweptSurface from PGeom inherits Surface from PGeom

        ---Purpose : A  swept surface  is  one that is constructed  by
        --         sweeping a curve by another curve.
        --         
	---See Also : SweptSurface from Geom.


uses Dir         from gp,
     Curve       from PGeom,
     SurfaceForm from GeomAbs, 
     Shape       from GeomAbs

is


    Initialize;
	---Purpose: Initializes the field(s) with default value(s).
    	---Level: Internal 


    Initialize(aBasisCurve: Curve from PGeom;
    	       aDirection: Dir from gp);
	---Purpose: Initialize the fields with these values.
    	---Level: Internal 


  BasisCurve (me: mutable; aBasisCurve: Curve from PGeom);
        ---Purpose : Set the value of the field basisCurve with <aBasisCurve>.
    	---Level: Internal 


  BasisCurve (me) returns Curve from PGeom;
        ---Purpose : Returns the value of the field basisCurve.
    	---Level: Internal 


  Direction (me: mutable; aDirection: Dir from gp);
        ---Purpose : Set the value of the field direction with <aDirection>.
    	---Level: Internal 


  Direction (me) returns Dir from gp;
        ---Purpose : Returns the value of the field direction.
    	---Level: Internal 


fields

  basisCurve : Curve       from PGeom   is protected;
  direction  : Dir         from gp      is protected;

end;
