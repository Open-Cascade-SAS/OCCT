-- Created on: 2002-12-12
-- Created by: data exchange team
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class DataEnvironment from StepRepr
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity DataEnvironment

uses
    HAsciiString from TCollection,
    HArray1OfPropertyDefinitionRepresentation from StepRepr

is
    Create returns DataEnvironment from StepRepr;
	---Purpose: Empty constructor

    Init (me: mutable; aName: HAsciiString from TCollection;
                       aDescription: HAsciiString from TCollection;
                       aElements: HArray1OfPropertyDefinitionRepresentation from StepRepr);
	---Purpose: Initialize all fields (own and inherited)

    Name (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Name
    SetName (me: mutable; Name: HAsciiString from TCollection);
	---Purpose: Set field Name

    Description (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Description
    SetDescription (me: mutable; Description: HAsciiString from TCollection);
	---Purpose: Set field Description

    Elements (me) returns HArray1OfPropertyDefinitionRepresentation from StepRepr;
	---Purpose: Returns field Elements
    SetElements (me: mutable; Elements: HArray1OfPropertyDefinitionRepresentation from StepRepr);
	---Purpose: Set field Elements

fields
    theName: HAsciiString from TCollection;
    theDescription: HAsciiString from TCollection;
    theElements: HArray1OfPropertyDefinitionRepresentation from StepRepr;

end DataEnvironment;
