-- Created on: 1992-06-22
-- Created by: Gilles DEBARBOUILLE
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

private class Sentence from Units 

	---Purpose: This class describes all the methods to create and
	--          compute an expression contained in a string.

uses

    Token          from Units,
    TokensSequence from Units,
    Lexicon        from Units

--raises

is

    Create(alexicon : Lexicon from Units ; astring : CString)
    
    ---Level: Internal 
    
    ---Purpose: Creates and  returns  a   Sentence, by  analyzing  the
    --          string <astring> with the lexicon <alexicon>.
    
    returns Sentence from Units;
    
    SetConstants(me : in out)
    
    ---Level: Internal 
    
    ---Purpose: For each constant encountered, sets the value.
    
    is static;
    
    Sequence(me) returns any TokensSequence from Units
    
    ---Level: Internal 
    
    ---C++: inline
    
    ---Purpose: Returns <thesequenceoftokens>.
    
    is static;
    
    Sequence(me : in out ; asequenceoftokens : any TokensSequence from Units)
    
    ---Level: Internal 
    
    ---C++: inline
    
    ---Purpose: Sets the field <thesequenceoftokens> to <asequenceoftokens>.
    
    is static;
    
    Evaluate(me : in out)returns Token from Units
    
    ---Level: Internal 
    
    ---Purpose: Computes and  returns in a   token the result  of  the
    --          expression.
    
    is static;
    
    IsDone(me) returns Boolean from Standard
    ---Level: Internal 
    ---C++: inline
    ---Purpose: Return True if number of created tokens > 0
    --          (i.e creation of sentence is succesfull)
    is static;

    Dump(me)
    
    ---Level: Internal 
    
    ---C++: inline
    
    ---Purpose: Useful for debugging.
    
    is static;

fields

    thesequenceoftokens : TokensSequence from Units;

end Sentence;
