-- Created on: 2000-05-10
-- Created by: Andrey BETENEV
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1

class RepItemGroup from StepAP214
inherits Group from StepBasic

    ---Purpose: Representation of STEP entity RepItemGroup

uses
    HAsciiString from TCollection,
    RepresentationItem from StepRepr

is
    Create returns RepItemGroup from StepAP214;
	---Purpose: Empty constructor

    Init (me: mutable; aGroup_Name: HAsciiString from TCollection;
                       hasGroup_Description: Boolean;
                       aGroup_Description: HAsciiString from TCollection;
                       aRepresentationItem_Name: HAsciiString from TCollection);
	---Purpose: Initialize all fields (own and inherited)

    RepresentationItem (me) returns RepresentationItem from StepRepr;
	---Purpose: Returns data for supertype RepresentationItem
    SetRepresentationItem (me: mutable; RepresentationItem: RepresentationItem from StepRepr);
	---Purpose: Set data for supertype RepresentationItem

fields
    theRepresentationItem: RepresentationItem from StepRepr; -- supertype

end RepItemGroup;
