-- Created on: 1992-11-17
-- Created by: Christian CAILLET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



deferred class Selection  from IFSelect  inherits TShared

    ---Purpose : A Selection allows to define a set of Interface Entities.
    --           Entities to be put on an output file should be identified in
    --           a way as independant from such or such execution as possible.
    --           This permits to handle comprehensive criteria, and to replay
    --           them when a new variant of an input file has to be processed.
    --         
    --           Its input can be, either an Interface Model (the very source),
    --           or another-other Selection(s) or any other ouput. All list
    --           computations start from an input Graph (from IFGraph)

uses AsciiString from TCollection, EntityIterator, Graph, SelectionIterator

raises InterfaceError

is

    RootResult (me; G : Graph) returns EntityIterator
    	raises InterfaceError  is deferred;
    ---Purpose : Returns the list of selected entities, computed from Input
    --           given as a Graph. Specific to each class of Selection
    --           Note that uniqueness of each entity is not required here
    --           This method can raise an exception as necessary

    HasUniqueResult (me) returns Boolean  is virtual protected;
    ---Purpose : Returns True if RootResult guarantees uniqueness for each
    --           Entity. Called by UniqueResult.
    --           Default answer is False. Can be redefined.

    UniqueResult (me; G : Graph) returns EntityIterator;
    ---Purpose : Returns the list of selected entities, each of them beeing
    --           unique. Default definition works from RootResult. According
    --           HasUniqueResult, UniqueResult returns directly RootResult,
    --           or build a Unique Result from it with a Graph.

    CompleteResult (me; G : Graph) returns EntityIterator  is virtual;
    ---Purpose : Returns the list of entities involved by a Selection, i.e.
    --           UniqueResult plus the shared entities (directly or not)


    FillIterator (me; iter : in out SelectionIterator)  is deferred;
    ---Purpose : Puts in an Iterator the Selections from which "me" depends
    --           (there can be zero, or one, or a list).
    --           Specific to each class of Selection

    Label (me) returns AsciiString from TCollection  is deferred;
    ---Purpose : Returns a text which defines the criterium applied by a
    --           Selection (can be used to be printed, displayed ...)
    --           Specific to each class

end Selection;
