-- Created on: 1992-11-27
-- Created by: Isabelle GRIGNON
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Domain from BRepGProp 

	---Purpose: Arc iterator. Returns only Forward and Reversed edges from 
        --          the face in an undigested order.

uses Face     from TopoDS,
     Edge     from TopoDS,
     Explorer from TopExp
is
  
  Create returns Domain;
        --- Purpose : Empty constructor. 
	---C++: inline
  
  Create (F : Face from TopoDS) returns Domain;
        --- Purpose : Constructor. Initializes the domain with the face.
	---C++: inline
  
  Init(me : in out;F : Face from TopoDS);
        --- Purpose : Initializes the domain with the face.
	---C++: inline
  
  More(me : in out)  returns Boolean from Standard
        --- Purpose :
        --  Returns True if there is another arc of curve in the list.
  ---C++: inline
  is static;
  
  Init(me : in out)
        --- Purpose : Initializes the exploration with the face already set.
        ---C++: inline
  is static;
  
  Value(me : in out) returns Edge from TopoDS  
        ---Purpose: Returns the current edge.
        ---C++: return const &
	---C++: inline
  is static;
  
  Next(me : in out)  
        --- Purpose :
        --  Sets the index of the arc iterator to the next arc of
        --  curve.
  is static;

fields

    myExplorer : Explorer from TopExp;

end Domain;




