--
-- File:	AlienImage_SGIRGBAlienImage.cdl
-- Created:	23/03/93
-- Author:	BBL
-- Modified:	02-06-98 : FMN ; Suppression appel Clear (deja fait dans ALienData)
--
---Copyright:	Matravision 1993
--

class SGIRGBAlienImage from AlienImage inherits AlienUserImage from AlienImage

    	---Purpose: Defines an SGI .rgb Alien image, i.e. an image using
    	-- the image format for Silicon Graphics workstations.

uses
	File 			from OSD,
	AsciiString 		from TCollection,
	ColorImage 		from Image,
	PseudoColorImage 	from Image,
	Image			from Image,
	SGIRGBAlienData 	from AlienImage

is
	Create returns mutable SGIRGBAlienImage from AlienImage;
    	---Purpose: Constructs an empty SGI .rgb Alien image.
    
	Clear( me : in out mutable) ;
	---Level: Public
	---Purpose: Frees memory allocated by SGIRGBAlienImage

	SetName( me : in out mutable;
		 aName : in AsciiString from TCollection) ;
	---Level: Public
	---Purpose: Set Image name .

	Name( me : in immutable ) returns AsciiString from TCollection ;
		  ---C++: return const &
    		  ---Purpose: Reads the  Image name .

	ToImage( me : in immutable ) 
	  returns mutable Image from Image ;
	---Level: Public
	---Purpose : Converts a SGIRGBAlienImage object to a Image object.

	FromImage( me : in out mutable ; anImage : in Image from Image ) ;
	---Level: Public
	---Purpose : Converts a Image object to a SGIRGBAlienImage object.

	Read ( me : in out mutable; afile : in out File from OSD )
	  returns Boolean from Standard ;
	---Purpose: Reads content of a SGIRGBAlienImage object from a file
	--          Returns True if file is a XWD file .

	Write( me : in immutable; afile : in out File from OSD )
	  returns Boolean from Standard ;
	---Purpose: Writes content of a SGIRGBAlienImage object to a file

fields
	myData : SGIRGBAlienData  from  AlienImage;

end ;
 
