-- Created on: 1995-06-22
-- Created by: Christophe MARION
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class BiPoint from HLRAlgo

uses
    Address from Standard,
    Boolean from Standard,
    Integer from Standard
    
is
    Create
    returns BiPoint from HLRAlgo; 
    	---C++: inline
    
    Create(X1,Y1,Z1,X2,Y2,Z2       : Real    from Standard;
           XT1,YT1,ZT1,XT2,YT2,ZT2 : Real    from Standard;
           Index                   : Integer from Standard;
           reg1,regn,outl,intl     : Boolean from Standard)
    returns BiPoint from HLRAlgo; 
    
    Create(X1,Y1,Z1,X2,Y2,Z2       : Real    from Standard;
           XT1,YT1,ZT1,XT2,YT2,ZT2 : Real    from Standard;
           Index                   : Integer from Standard;
           flag                    : Boolean from Standard)
    returns BiPoint from HLRAlgo; 
    
    Create(X1,Y1,Z1,X2,Y2,Z2       : Real    from Standard;
           XT1,YT1,ZT1,XT2,YT2,ZT2 : Real    from Standard;
           Index,i1,i1p1,i1p2      : Integer from Standard;
           reg1,regn,outl,intl     : Boolean from Standard)
    returns BiPoint from HLRAlgo; 
    
    Create(X1,Y1,Z1,X2,Y2,Z2       : Real    from Standard;
           XT1,YT1,ZT1,XT2,YT2,ZT2 : Real    from Standard;
           Index,i1,i1p1,i1p2      : Integer from Standard;
           flag                    : Boolean from Standard)
    returns BiPoint from HLRAlgo; 
    
    Create(X1,Y1,Z1,X2,Y2,Z2               : Real    from Standard;
           XT1,YT1,ZT1,XT2,YT2,ZT2         : Real    from Standard;
           Index,i1,i1p1,i1p2,i2,i2p1,i2p2 : Integer from Standard;
           reg1,regn,outl,intl             : Boolean from Standard)
    returns BiPoint from HLRAlgo; 
    
    Create(X1,Y1,Z1,X2,Y2,Z2               : Real    from Standard;
           XT1,YT1,ZT1,XT2,YT2,ZT2         : Real    from Standard;
           Index,i1,i1p1,i1p2,i2,i2p1,i2p2 : Integer from Standard;
           flag                            : Boolean from Standard)
    returns BiPoint from HLRAlgo; 
    
    Rg1Line(me) returns Boolean from Standard
    	---C++: inline
    is static;

    Rg1Line(me : in out; B : Boolean from Standard)
    	---C++: inline
    is static;

    RgNLine(me) returns Boolean from Standard
    	---C++: inline
    is static;

    RgNLine(me : in out; B : Boolean from Standard)
    	---C++: inline
    is static;

    OutLine(me) returns Boolean from Standard
    	---C++: inline
    is static;

    OutLine(me : in out; B : Boolean from Standard)
    	---C++: inline
    is static;

    IntLine(me) returns Boolean from Standard
    	---C++: inline
    is static;

    IntLine(me : in out; B : Boolean from Standard)
    	---C++: inline
    is static;

    Hidden(me) returns Boolean from Standard
    	---C++: inline
    is static;

    Hidden(me : in out; B : Boolean from Standard)
    	---C++: inline
    is static;

    Indices(me) returns Address from Standard
    	---C++: inline
    is static;

    Coordinates(me) returns Address from Standard
    	---C++: inline
    is static;

fields
    myIndices     : Integer from Standard[10];
    myCoordinates : Real    from Standard[12];
    
end BiPoint;
