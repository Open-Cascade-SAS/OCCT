-- Created on: 1992-06-22
-- Created by: Gilles DEBARBOUILLE
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

private class UnitSentence from Units

	---Purpose: This   class describes   all    the  facilities to
	--          manipulate and compute units contained in a string
	--          expression.

inherits

    Sentence from Units

uses

    QuantitiesSequence from Units

--raises

is

    Create(astring : CString)
    
    ---Level: Internal 
    
    ---Purpose: Creates   and   returns a   UnitSentence.   The string
    --          <astring> describes in natural  language the  unit  or
    --          the composed unit to be analysed.
    
    returns UnitSentence from Units;
    
    Create(astring : CString ; aquantitiessequence : QuantitiesSequence from Units)
    
    ---Level: Internal 
    
    ---Purpose: Creates  and returns    a  UnitSentence.  The   string
    --          <astring> describes in natural language the unit to be
    --          analysed.   The    sequence     of physical quantities
    --          <asequenceofquantities>   describes    the   available
    --          dictionary of units you want to use.
    
    returns UnitSentence from Units;
    
    Analyse(me : in out)
    
    ---Level: Internal 
    
    ---Purpose: Analyzes   the sequence  of   tokens  created  by  the
    --          constructor to  find  the true significance   of  each
    --          token.
    
    is static;
    
    SetUnits(me : in out ; aquantitiessequence : QuantitiesSequence from Units)
    
    ---Level: Internal 
    
    ---Purpose: For each token which  represents a unit, finds  in the
    --          sequence    of    physical   quantities      all   the
    --          characteristics of the unit found.
    
    is static;

--fields

end UnitSentence;
