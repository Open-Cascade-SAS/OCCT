-- Created on: 1992-09-28
-- Created by: Remi GILET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class MakeConicalSurface from GC inherits Root from GC

    	---Purpose : This class implements the following algorithms used 
    	--           to create a ConicalSurface from Geom.
    	--           * Create a ConicalSurface parallel to another and passing 
    	--             through a point.
    	--           * Create a ConicalSurface parallel to another at a distance
    	--             <Dist>.
    	--           * Create a ConicalSurface by 4 points.
    	--           * Create a ConicalSurface by its axis and 2 points.
    	--           * Create a ConicalSurface by 2 points and 2 radius.
        --  The local coordinate system of the ConicalSurface is defined
        --  with an axis placement (see class ElementarySurface).
        -- 
        --  The "ZAxis" is the symmetry axis of the ConicalSurface, 
        --  it gives the direction of increasing parametric value V.
        --  The apex of the surface is on the negative side of this axis.
        -- 
        --  The parametrization range is  :
        --     U [0, 2*PI],  V ]-infinite, + infinite[
        --     
        --  The "XAxis" and the "YAxis" define the placement plane of the 
        --  surface (Z = 0, and parametric value V = 0)  perpendicular to 
        --  the symmetry axis. The "XAxis" defines the origin of the 
        --  parameter U = 0.  The trigonometric sense gives the positive 
        --  orientation for the parameter U.
        -- 
        --  When you create a ConicalSurface the U and V directions of
        --  parametrization are such that at each point of the surface the
        --  normal is oriented towards the "outside region".

uses Pnt            from gp,
     Ax1            from gp,
     Ax2            from gp,
     Lin            from gp,
     Cone           from gp,
     ConicalSurface from Geom,
     Real           from Standard

raises NotDone from StdFail

is

Create (A2     : Ax2  from gp      ; 
    	Ang    : Real from Standard; 
    	Radius : Real from Standard) returns MakeConicalSurface;
    	--- Purpose :
    	--  A2 defines the local coordinate system of the conical surface.
    	--  Ang is the conical surface semi-angle ]0, PI/2[.
    	--  Radius is the radius of the circle Viso in the placement plane 
    	--  of the conical surface defined with "XAxis" and "YAxis".
    	--  The "ZDirection" of A2 defines the direction of the surface's
    	--  axis of symmetry.
    	--  If the location point of A2 is the apex of the surface 
    	--  Radius = 0 .
    	--  At the creation the parametrization of the surface is defined
    	--  such that the normal Vector (N = D1U ^ D1V) is oriented towards
    	-- the "outside region" of the surface. 
	--  Status is "NegativeRadius" if Radius < 0.0 or "BadAngle" if
    	--  Ang < Resolution from gp or Ang >= PI/ - Resolution

Create (C : Cone from gp) returns MakeConicalSurface;
    	--- Purpose : Creates a ConicalSurface from a non persistent Cone from package gp.

Create(Cone  : Cone from gp;
       Point : Pnt  from gp) returns MakeConicalSurface;
    	---Purpose : Make a ConicalSurface from Geom <TheCone> parallel to another 
    	--           ConicalSurface <Cone> and passing through a Pnt <Point>.

Create(Cone : Cone  from gp      ;
       Dist : Real  from Standard) returns MakeConicalSurface;
    	---Purpose : Make a ConicalSurface from Geom <TheCone> parallel to another 
    	--           ConicalSurface <Cone> at the distance <Dist> which can 
    	--           be greater or lower than zero.

Create(P1     :     Pnt from gp;
       P2     :     Pnt from gp;
       P3     :     Pnt from gp;
       P4     :     Pnt from gp) returns MakeConicalSurface;
    	---Purpose : Make a ConicalSurface from Geom <TheCone> passing through 3
    	--           Pnt <P1>,<P2>,<P3>.
    	--           Its axis is <P1P2> and the radius of its base is
    	--           the distance between <P3> and <P1P2>.
    	--           The distance between <P4> and <P1P2> is the radius of 
    	--           the section passing through <P4>.
    	--           An error iss raised if <P1>,<P2>,<P3>,<P4> are 
    	--           colinear or if <P3P4> is perpendicular to <P1P2> or 
    	--           <P3P4> is colinear to <P1P2>.

Create(Axis   : Ax1  from gp;
       P1,P2  : Pnt  from gp) returns MakeConicalSurface;
    	---Purpose: Make a ConicalSurface by its axis <Axis> and and two points.

Create(Axis   : Lin  from gp;
       P1,P2  : Pnt  from gp) returns MakeConicalSurface;
    	---Purpose: Make a ConicalSurface by its axis <Axis> and and two points.

Create(P1     :     Pnt  from gp      ;
       P2     :     Pnt  from gp      ;
       R1     :     Real from Standard;
       R2     :     Real from Standard) returns MakeConicalSurface;
    	---Purpose: Make a ConicalSurface with two points and two radius.
    	--          The axis of the solution is the line passing through 
    	--          <P1> and <P2>.
    	--          <R1> is the radius of the section passing through <P1> 
    	--          and <R2> the radius of the section passing through <P2>.

Value(me) returns ConicalSurface from Geom
    raises NotDone
    is static;
    	---Purpose: Returns the constructed cone.
    	-- Exceptions
    	-- StdFail_NotDone if no cone is constructed.
    	---C++: return const&

Operator(me) returns ConicalSurface from Geom
    is static;
    	---C++: return const&
    	---C++: alias "Standard_EXPORT operator Handle_Geom_ConicalSurface() const;"

fields

    TheCone : ConicalSurface from Geom;
    --The solution from Geom.
    
end MakeConicalSurface;
