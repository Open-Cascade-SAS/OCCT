-- Created on: 1997-10-02
-- Created by: Xuan Trang PHAM PHU
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ShellToSolid from TopOpeBRepBuild

---Purpose: 
-- This class builds solids from a set of shells SSh and a solid F. 

uses

    Shell from TopoDS,
    Solid from TopoDS,
    ListOfShape from TopTools

is

    Create returns ShellToSolid;
     
    Init(me : in out)
    is static;
    
    AddShell(me : in out; Sh : Shell from TopoDS)
    is  static;
     	
    MakeSolids(me : in out; 
    	       So : Solid from TopoDS;
    	       LSo : in out ListOfShape from TopTools)
    is static;

fields 

    myLSh : ListOfShape from TopTools;
    
end ShellToSolid;
