-- Created on: 1997-02-12
-- Created by: Alexander BRIVIN
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Transform from Vrml 

	---Purpose:  defines a Transform of VRML specifying transform
	---          properties.
    	--  This  node  defines  a  geometric  3D  transformation   consisting   of  (in  order) 
    	--  a  (possibly)  non-uniform  scale  about  an  arbitrary  point,  a  rotation  about 
    	--  an arbitrary point  and  axis  and  translation. 
    	--  By  default  : 
	--    myTranslation (0,0,0) 
	--    myRotation  (0,0,1,0)
	--    myScaleFactor (1,1,1)
	--    myScaleOrientation (0,0,1,0)
	--    myCenter (0,0,0)

uses
 
   Vec         from  gp, 
   SFRotation  from  Vrml

is
 
    Create returns  Transform from Vrml; 
 
    Create ( aTranslation      : Vec         from  gp; 
    	     aRotation         : SFRotation  from  Vrml; 
    	     aScaleFactor      : Vec         from  gp; 
    	     aScaleOrientation : SFRotation  from  Vrml; 
             aCenter           : Vec         from  gp )
    	returns  Transform from Vrml; 

    SetTranslation ( me : in out;  aTranslation : Vec  from  gp );
    Translation ( me )  returns Vec  from  gp;

    SetRotation ( me : in out;  aRotation : SFRotation  from  Vrml );
    Rotation ( me )  returns  SFRotation  from  Vrml;

    SetScaleFactor ( me : in out;  aScaleFactor : Vec  from  gp );
    ScaleFactor ( me )  returns Vec  from  gp;

    SetScaleOrientation ( me : in out;  aScaleOrientation : SFRotation  from  Vrml );
    ScaleOrientation ( me  )  returns  SFRotation  from  Vrml;

    SetCenter ( me : in out;  aCenter : Vec  from  gp );
    Center ( me )  returns Vec  from  gp;

    Print  ( me;  anOStream: in out OStream from Standard) returns OStream from Standard;
    ---C++:  return  & 

fields
 
    myTranslation      : Vec         from  gp;   -- Translation vector
    myRotation         : SFRotation  from  Vrml; -- Rotation
    myScaleFactor      : Vec         from  gp;   -- Scale factors
    myScaleOrientation : SFRotation  from  Vrml; -- Defines rotational space for scale
    myCenter           : Vec         from  gp;   -- Center point for scale and rotate

end Transform;
