-- Created on: 1993-02-22
-- Created by: Philippe DAUTRY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class BezierCurve from PGeom inherits BoundedCurve from PGeom

        ---Purpose : Defines a rational or non rational Bezier curve.
        --         
	---See Also : BezierCurve from Geom.

uses  HArray1OfReal from PColStd,
      HArray1OfPnt  from PColgp

is 


  Create returns mutable BezierCurve from PGeom;
        ---Purpose : Creates a non rational  Bezier curve with default
        --         values.
    	---Level: Internal 

  Create(aPoles    : HArray1OfPnt;
         aWeights  : HArray1OfReal;
	 aRational : Boolean from Standard)
     returns mutable BezierCurve from PGeom;
        ---Purpose : Creates a non rational Bezier curve with a set of
        --         poles aCurvePoles and a set of weights aPoleWeight.
    	---Level: Internal 


  Rational (me: mutable; aRational: Boolean from Standard);
        ---Purpose : Set the value of the field rational with <aRational>.
    	---Level: Internal 


  Rational (me) returns Boolean;
        ---Purpose : Returns the value of the field rational.
    	---Level: Internal 


  Poles (me: mutable; aPoles : HArray1OfPnt from PColgp);
        ---Purpose : Set the value of the field poles with <aPoles>.
    	---Level: Internal 


  Poles (me) returns HArray1OfPnt from PColgp;
        ---Purpose : Returns the value of the field poles.
    	---Level: Internal 


  Weights (me: mutable; aWeights : HArray1OfReal from PColStd);
        ---Purpose : Set the value of the field weights.
    	---Level: Internal 


  Weights (me)returns HArray1OfReal from PColStd;
        ---Purpose : Returns the value of the field weights.
    	---Level: Internal 


fields

   rational : Boolean from Standard;
   poles    : HArray1OfPnt  from PColgp;
   weights  : HArray1OfReal from PColStd;

end;
