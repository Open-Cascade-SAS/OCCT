-- File:	IntTools_ShrunkRange.cdl
-- Created:	Sun Mar 11 10:31:46 2001
-- Author:	Peter KURNEV
--		<pkv@irinox>
---Copyright:	 Matra Datavision 2001


class ShrunkRange from IntTools 

	---Purpose:  
	---  The class provides the computation of 
	---  a working (shrunk) range [t1, t2] for 
    	---  the 3D-curve of the edge. 
	 
uses
 
    Edge from TopoDS, 
    Vertex from TopoDS, 
    Range from IntTools, 
    Box from Bnd, 
    Context from IntTools 

--raises

is 
    Create 
    	returns ShrunkRange from IntTools;
	---Purpose:
	--- Empty constructor
	---
	
    Create (aE  : Edge from TopoDS; 
	    aV1 : Vertex from TopoDS;              
	    aV2 : Vertex from TopoDS;              
    	    aR  : Range from IntTools; 
    	    ICtx: Context from IntTools)   
	returns ShrunkRange from IntTools;
	---Purpose:
	---
    SetContext(me:out; 
    	  aContext : Context from IntTools); 
    ---Purpose:
	--- Sets the intersecton context
	--- 
    Context(me) 
    	returns Context from IntTools; 
    ---C++:  return const &   
     ---Purpose:
	--- Gets the intersecton context
	---
 
 
    SetShrunkRange(me:out;  aR:Range from IntTools);
    	---Purpose:
	--- Sets an shrunk range
	---

    ShrunkRange(me) 
    	returns Range from IntTools; 
    	---C++:  return  const& 
	---Purpose:
	--- Returns shrunk range
	---
  
    BndBox  (me) 
    	returns Box from Bnd; 
    	---C++:  return  const& 
	---Purpose:
	--- Returns bounding box for edge restricted
	--- by shrunk range
	---
     
    Edge  (me) 
    	returns Edge from TopoDS; 
    	---C++:  return  const&	 
	---Purpose:
	--- Returns edge for which 
	--- the shrunk range is computed
	---
	     
    Perform(me:out); 
    	---Purpose:
	--- Computes shrunk range for
	--- an edge given in constructor
	--- 
    	
	 
    IsDone (me) 
	returns Boolean from Standard; 
	---Purpose:
	--- Returns true if no error occured
	--- during shrunk range computation
	---
	 
    ErrorStatus(me) 
    	returns Integer from Standard;  
	---Purpose:
	--- Returns code of computing shrunk range
	--- completion
	--- 0 - means successful completion
	--- 1 - nothing has been done
	--- 2 - initial range is out of edge's range
	--- 3 - first boundary of initial range is more than
	---     last boundary
	--- 4 - projection of first vertex failed
	--- 5 - projection of second vertex failed
	--- 6 - shrunk range can not be computed
	---     shrunk range is setted to initial range
	---

fields
    myEdge        :  Edge from TopoDS; 
    myV1          :  Vertex from TopoDS;
    myV2          :  Vertex from TopoDS; 
    myRange       :  Range from IntTools; 
    myShrunkRange :  Range from IntTools; 
    myBndBox      :  Box from Bnd;  
    myContext     :  Context from IntTools;
    myIsDone      :  Boolean from Standard; 
    myErrorStatus :  Integer from Standard;   
     
end ShrunkRange;
