-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class FIR from TopOpeBRepDS 

---Purpose: FaceInterferenceReducer

uses

    DataMapOfShapeListOfShapeOn1State from TopOpeBRepDS,
    HDataStructure from TopOpeBRepDS

is

    Create(HDS : HDataStructure) returns FIR from TopOpeBRepDS;
    ProcessFaceInterferences(me:out;M:DataMapOfShapeListOfShapeOn1State);
    ProcessFaceInterferences(me:out;I:Integer;M:DataMapOfShapeListOfShapeOn1State);

fields

    myHDS : HDataStructure from TopOpeBRepDS;
    
end FIR from TopOpeBRepDS;
