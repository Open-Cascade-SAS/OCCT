-- Created on: 1993-10-18
-- Created by: Christophe MARION
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class EdgeFaceTool from HLRBRep

	---Purpose: The EdgeFaceTool computes the  UV coordinates at a
	--          given parameter on a Curve and a Surface.  It also
	--          compute the signed  curvature value in a direction
	--          at a given u,v point on a surface.

uses
    Address  from Standard,
    Boolean  from Standard,
    Real     from Standard,
    Dir      from gp

is
    CurvatureValue(myclass;
                   F  : Address from Standard; -- as Surface from HLRBRep
                   U  : Real    from Standard;
                   V  : Real    from Standard;
                   Tg : Dir     from gp)       -- as tangent of the  edge
    returns Real from Standard;                -- at U,V point.
    
    UVPoint(myclass;
            Par :     Real    from Standard;
            E   :     Address from Standard; -- as Curve   from HLRBRep
            F   :     Address from Standard; -- as Surface from HLRBRep
	    U,V : out Real    from Standard)
    	---Purpose: return True if U and V are found.
    returns Boolean from Standard;
    
end EdgeFaceTool;
