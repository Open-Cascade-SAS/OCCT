-- Created on: 1995-12-21
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class SolidBuilder from TopOpeBRepBuild 

uses

    Shape from TopoDS,
    
    ShapeSet from TopOpeBRepBuild,
    LoopSet from TopOpeBRepBuild,
    BlockIterator from TopOpeBRepBuild,
    BlockBuilder from TopOpeBRepBuild,

    ShellFaceSet from TopOpeBRepBuild,
    SolidAreaBuilder from TopOpeBRepBuild
    
is

    Create returns SolidBuilder;

    Create(FS : in out ShellFaceSet; ForceClass : Boolean = Standard_False)  
    returns SolidBuilder;
    ---Purpose: Create a SolidBuilder to build the areas on
    -- the shapes (shells, blocks of faces) described by <LS>.

    InitSolidBuilder(me : in out; 
    	    	     FS : in out ShellFaceSet;
    	    	     ForceClass : Boolean) is static;
    
    -- Output methods 
    InitSolid(me : in out) returns Integer from Standard;
    MoreSolid(me) returns Boolean from Standard is static;
    NextSolid(me : in out) is static;
    
    -- Exploration of the wires of the current Solid
    InitShell(me : in out) returns Integer from Standard;
    MoreShell(me) returns Boolean from Standard is static;
    NextShell(me : in out) is static;
    IsOldShell(me) returns Boolean from Standard is static;
    OldShell(me) returns Shape from TopoDS is static;
    ---Purpose: Returns current shell
    -- This shell may be : 
    -- * an old shell OldShell(), which has not been reconstructed;
    -- * a new shell made of faces described by ...NewFace() methods.
    ---C++: return const &

    -- Exploration of the faces of current shell when IsOldShell = False
    InitFace(me : in out) returns Integer from Standard;
    MoreFace(me) returns Boolean from Standard is static;
    NextFace(me : in out) is static;
    Face(me) returns Shape from TopoDS is static;
    ---Purpose: Returns current new face of current new shell.
    ---C++: return const &

    --- private
    MakeLoops(me : in out; SS : in out ShapeSet from TopOpeBRepBuild) 
    is static private;
    
fields

    myLoopSet : LoopSet from TopOpeBRepBuild;
    myBlockIterator : BlockIterator from TopOpeBRepBuild;
    myBlockBuilder : BlockBuilder from TopOpeBRepBuild;

    mySolidAreaBuilder : SolidAreaBuilder from TopOpeBRepBuild;
    
end SolidBuilder;
