-- Created on: 1999-06-17
-- Created by: Vladislav ROMASHKO
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class TreeNode from PDataStd inherits Attribute from PDF 

uses 
     
    Attribute from PDF, 
    GUID      from Standard 

is

    Create returns TreeNode from PDataStd;
        
    First(me) returns TreeNode from PDataStd;
	 
    SetFirst(me : mutable; F : TreeNode from PDataStd);    
    
    Next(me) returns TreeNode from PDataStd;
        
    SetNext(me : mutable; F : TreeNode from PDataStd);    
    
    SetTreeID(me : mutable; GUID : GUID from Standard);

    GetTreeID(me) returns GUID from Standard;

fields

    myFirst  : TreeNode from PDataStd;  
    myNext   : TreeNode from PDataStd;  
    myTreeID : GUID     from Standard;

end TreeNode;
 
