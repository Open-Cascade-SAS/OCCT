-- Created on: 1992-07-21
-- Created by: Laurent PAINNOT
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.





generic class CurveLocator from Extrema 
    (Curve1 as any;
     Tool1  as any;   -- as ToolCurve(Curve1)
     Curve2 as any;
     Tool2  as any;   -- as ToolCurve(Curve2)
     POnC   as any;
     Pnt    as any)
					
     
is

    Locate (myclass; P: Pnt; C: Curve1; NbU: Integer; Papp: out POnC);
    ---Purpose: Among a set of points {C(ui),i=1,NbU}, locate the point
    --          P=C(uj) such that:
    --           distance(P,C) = Min{distance(P,C(ui))}


    Locate (myclass; P: Pnt; C: Curve1; NbU: Integer; Umin, Usup: Real;Papp: out POnC);
    ---Purpose: Among a set of points {C(ui),i=1,NbU}, locate the point
    --          P=C(uj) such that:
    --           distance(P,C) = Min{distance(P,C(ui))}
    --           The research is done between umin and usup.


   Locate (myclass; C1: Curve1; C2: Curve2; NbU, NbV: Integer; Papp1, Papp2: out POnC);
    ---Purpose: Among two sets of points {C1(ui),i=1,NbU} and
    --          {C2(vj),j=1,NbV}, locate the two points P1=C1(uk) and 
    --          P2=C2(vl) such that:
    --           distance(P1,P2) = Min {distance(C1(ui),C2(vj))}.


end CurveLocator;
