-- Copyright (c) 2003-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class Modification from ShapeCustom inherits Modification from BRepTools

        ---Purpose: A base class of Modification's from ShapeCustom.
	--          Implements message sending mechanism.

uses
    Shape from TopoDS,
    Msg from Message,
    Gravity from Message,
    BasicMsgRegistrator from ShapeExtend

is

    SetMsgRegistrator (me:mutable; msgreg: BasicMsgRegistrator from ShapeExtend) is virtual;
	---Purpose: Sets message registrator

    MsgRegistrator (me) returns BasicMsgRegistrator from ShapeExtend;
    	---Purpose: Returns message registrator

    SendMsg (me; shape  : Shape from TopoDS;
                 message: Msg from Message;
                 gravity: Gravity from Message = Message_Info);
    	---Purpose: Sends a message to be attached to the shape.
	--          Calls corresponding message of message registrator.

fields

    myMsgReg: BasicMsgRegistrator from ShapeExtend;

end SweptToElementary;
