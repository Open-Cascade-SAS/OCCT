-- Created on: 1996-01-22
-- Created by: Philippe MANGIN
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class GaussSetIntegration from math
    ---Purpose: -- This class implements the integration of a set of N
    --              functions of M  variables variables between the
    --              parameter bounds Lower[a..b] and Upper[a..b].
    --  Warning: - The case M>1 is not implemented.


uses Vector from math,
     IntegerVector from math, 
     FunctionSet from math,
     OStream from Standard,
     NotDone from StdFail

raises NotDone, NotImplemented

is

     Create(F: in out FunctionSet; Lower, Upper: Vector;
     	    Order: IntegerVector)
     ---Purpose:
     -- The Gauss-Legendre integration with Order = points of 
     -- integration for each unknow, is done on the function F 
     -- between the bounds Lower and Upper.
     returns GaussSetIntegration     
     raises  NotImplemented;
     
     IsDone(me)
     	---Purpose: returns True if all has been correctly done.
    	---C++: inline

     returns Boolean
     is static;
     
     Value(me)
     	---Purpose: returns the value of the integral.
    	---C++: inline
    	---C++: return const&

     returns Vector
     raises NotDone
     is static;


    Dump(me; o: in out OStream)
    	---Purpose: Prints information on the current state of the object.
    is static;




fields

Val: Vector;
Done: Boolean;

end GaussSetIntegration;
