-- Created on: 1994-02-14
-- Created by: model
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

generic class GenHSurface from Adaptor3d
    (TheSurface as Surface from Adaptor3d)
 
inherits HSurface from Adaptor3d 
    
	---Purpose: Generic class used to create a surface manipulated
      	--          with Handle from a surface described by the class Surface. 
	
uses

     Surface      from Adaptor3d


raises

    OutOfRange          from Standard,
    NoSuchObject        from Standard,
    DomainError         from Standard


is

    Create
    
	---Purpose: Creates an empty GenHSurface.
    	returns mutable GenHSurface from Adaptor3d; 
    

    Create(S: TheSurface)
    
	---Purpose: Creates a GenHSurface from a Surface.
    	returns mutable GenHSurface from Adaptor3d; 


    Set(me: mutable; S: TheSurface)
    
	---Purpose: Sets the field of the GenHSurface.
    	is static;

    --
    --  Access to the surface
    --  
    
    Surface(me) returns Surface from Adaptor3d;
	---Purpose: Returns a reference to the Surface inside the HSurface.
	--          This is redefined from HSurface, cannot be inline.
	--          
	---C++: return const &

    ChangeSurface(me : mutable)
    
	---Purpose: Returns the surface used to create the GenHSurface.
	--          
	---C++: return &
	---C++: inline

    	returns TheSurface;


fields

    mySurf: TheSurface is protected;

end GenHSurface;
