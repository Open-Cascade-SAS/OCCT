-- File:      HLRAppli_ReflectLines.cdl
-- Created:   05.12.12 15:53:35
-- Created by: Julia GERASIMOVA
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ReflectLines from HLRAppli

        ---Purpose : This class builds reflect lines on a shape
        --         according to the axes of view defined by user.
        --         Reflect lines are represented by edges in 3d.


uses
    Shape from TopoDS,
    Projector from HLRAlgo
    
is 
    Create(aShape : Shape from TopoDS)
    ---Purpose: Constructor
    --
    returns ReflectLines from HLRAppli;
    
    SetAxes(me: in out;
    	    Nx,  Ny,  Nz  : Real from Standard;
    	    XAt, YAt, ZAt : Real from Standard;
	    XUp, YUp, ZUp : Real from Standard);
	---Purpose: Sets the normal to the plane of visualisation,
	--          the coordinates of the view point and
	--          the coordinates of the vertical direction vector.

    Perform(me: in out);
    
    GetResult(me)
    returns Shape from TopoDS;
	---Purpose: returns resulting compound of reflect lines
	--          represented by edges in 3d
   
fields

    myProjector : Projector from HLRAlgo;
    myShape     : Shape     from TopoDS;
    myCompound  : Shape     from TopoDS;
    
end ReflectLines;
