-- Created by: Robert COUBLANC
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class SensitiveText2d from StdSelect inherits SensitiveEntity from 
Select2D

	---Purpose:  A framework to define a sensitive text entity for 2D views.
        
uses
    ExtendedString  from TCollection,
    EntityOwner     from SelectBasics,
    ListOfBox2d     from SelectBasics,
    Projector       from Select2D,
    Array1OfPnt2d   from TColgp,
    Box2d from Bnd
    
is

    Create(anOwnerId : EntityOwner from SelectBasics;
    	   aString   : ExtendedString from TCollection;
    	   XPox,YPos : Real from Standard;
    	   Angle     : Real = 0;
    	   aFontIndex: Integer = -1)
    returns mutable SensitiveText2d from StdSelect;
    	---Purpose: Constructs a sensitive 2D text object defined by the
    	-- owner anOwnerId, the string aString, the point
    	-- defined by the parameters XPos and YPos, the angle
    	-- Angle and the font index aFontIndex. 

    NeedsConversion (me) returns Boolean is redefined static;
    	---Purpose: returns Standard_True 
    	---Level: Public 
    	---C++: inline

    Convert(me:mutable; aTextProj : Projector from Select2D) is redefined virtual;
    	---Purpose: gets the size of the text in the 2d view 
    	---Level: Public 


    Areas(me:mutable; aresult : in out ListOfBox2d from SelectBasics) is redefined static;  
    	---Level: Public 
    	---Purpose: to be implemented specifically by each type of
    	--          sensitive  primitive .
    	--          
    
    Matches (me  :mutable; 
             X,Y : Real from Standard;
             aTol: Real from Standard;
             DMin: out Real from Standard) 
    returns Boolean
    is redefined static;

    Matches (me  :mutable; 
             XMin,YMin,XMax,YMax : Real from Standard;
             aTol: Real from Standard)
    returns Boolean
    is redefined static;

    Matches (me  :mutable; 
             Polyline:Array1OfPnt2d from TColgp;
	     aBox:Box2d from Bnd;
             aTol: Real from Standard)
    returns Boolean
    is redefined static;

fields

    mytext : ExtendedString from TCollection;
    myxpos : Real;
    myypos : Real;
    myangle: Real;
    myfont : Integer;

    myinitbox: Box2d from Bnd; --box before rotation...

end SensitiveText2d;
