-- Created on: 1991-02-21
-- Created by: Isabelle GRIGNON
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class   ExtPElS from Extrema
    	---Purpose: It calculates all the extremum distances
    	--          between a point and a surface.
    	--          These distances can be minimum or maximum.

uses   	POnSurf  from Extrema,
    	Cone     from gp,
	Pln      from gp,
    	Cylinder from gp,
    	Pnt      from gp,
    	Sphere   from gp,
    	Torus    from gp

raises  NotDone from StdFail,
    	OutOfRange

is
    Create returns ExtPElS;
    
    Create (P: Pnt; S: Cylinder; Tol: Real) returns ExtPElS;
      	---Purpose: It calculates all the distances between a point 
      	--          and a cylinder from gp.
      	--          Tol is used to test if the point is on the axis.

    Perform(me: in out; P: Pnt; S: Cylinder; Tol: Real) 
    is static;

    Create (P: Pnt; S: Pln; Tol: Real) returns ExtPElS;
      	---Purpose: It calculates all the distances between a point 
      	--          and a plane from gp.
      	--          Tol is used to test if the point is on the plane.

    Perform(me: in out; P: Pnt; S: Pln; Tol: Real) 
    is static;


    Create (P: Pnt; S: Cone; Tol: Real) returns ExtPElS;
      	---Purpose: It calculates all the distances between a point 
      	--          and a cone from gp.
      	--          Tol is used to test if the point is at the apex or
      	--          on the axis.

    Perform(me: in out;P: Pnt; S: Cone; Tol: Real)
    is static;
    
    Create (P: Pnt; S: Torus; Tol: Real) returns ExtPElS;
      	---Purpose: It calculates all the distances between a point 
      	--          and a torus from gp.
      	--          Tol is used to test if the point is on the axis.
    
    Perform(me: in out; P: Pnt; S: Torus; Tol: Real)
    is static;

    Create (P: Pnt; S: Sphere; Tol: Real) returns ExtPElS;
      	---Purpose: It calculates all the distances between a point 
      	--          and a sphere from gp.
      	--          Tol is used to test if the point is at the center.
    
    Perform(me: in out; P: Pnt; S: Sphere; Tol: Real)
    is static;


    IsDone (me) returns Boolean
    	---Purpose: Returns True if the distances are found.
    	is static;
    
    NbExt (me) returns Integer
    	---Purpose: Returns the number of extremum distances.
    	raises  NotDone from StdFail
	    	-- if IsDone(me)=False.
    	is static;

    SquareDistance (me; N: Integer) returns Real
    	---Purpose: Returns the value of the Nth resulting square distance.
    	raises  NotDone from StdFail,
    	    	-- if IsDone(me)=False.
    	        OutOfRange
		-- if N < 1 or N > NbPoints(me).
    	is static;

    Point (me; N: Integer) returns POnSurf
        ---C++: return const &
    	---Purpose: Returns the point of the Nth resulting distance.
    	raises  NotDone from StdFail,
    	    	-- if IsDone(me)=False.
    	        OutOfRange
		-- if N < 1 or N > NbPoints(me).
    	is static;

fields
    myDone : Boolean;
    myNbExt: Integer;
    mySqDist: Real [4];
    myPoint: POnSurf from Extrema [4];

end ExtPElS;
