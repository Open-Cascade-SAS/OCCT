-- File:	StepFEA_FeaTangentialCoefficientOfLinearThermalExpansion.cdl
-- Created:	Thu Dec 12 17:51:06 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class FeaTangentialCoefficientOfLinearThermalExpansion from StepFEA
inherits FeaMaterialPropertyRepresentationItem from StepFEA

    ---Purpose: Representation of STEP entity FeaTangentialCoefficientOfLinearThermalExpansion

uses
    HAsciiString from TCollection,
    SymmetricTensor23d from StepFEA

is
    Create returns FeaTangentialCoefficientOfLinearThermalExpansion from StepFEA;
	---Purpose: Empty constructor

    Init (me: mutable; aRepresentationItem_Name: HAsciiString from TCollection;
                       aFeaConstants: SymmetricTensor23d from StepFEA);
	---Purpose: Initialize all fields (own and inherited)

    FeaConstants (me) returns SymmetricTensor23d from StepFEA;
	---Purpose: Returns field FeaConstants
    SetFeaConstants (me: mutable; FeaConstants: SymmetricTensor23d from StepFEA);
	---Purpose: Set field FeaConstants

fields
    theFeaConstants: SymmetricTensor23d from StepFEA;

end FeaTangentialCoefficientOfLinearThermalExpansion;
