-- File:	RWStepShape_RWConnectedEdgeSet.cdl
-- Created:	Fri Dec 28 16:02:00 2001 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class RWConnectedEdgeSet from RWStepShape

    ---Purpose: Read & Write tool for ConnectedEdgeSet

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    ConnectedEdgeSet from StepShape

is
    Create returns RWConnectedEdgeSet from RWStepShape;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : ConnectedEdgeSet from StepShape);
	---Purpose: Reads ConnectedEdgeSet

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: ConnectedEdgeSet from StepShape);
	---Purpose: Writes ConnectedEdgeSet

    Share (me; ent : ConnectedEdgeSet from StepShape;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWConnectedEdgeSet;
