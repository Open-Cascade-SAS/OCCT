-- File:	StepRepr_CompositeShapeAspect.cdl
-- Created:	Tue Apr 24 13:43:49 2001
-- Author:	Christian CAILLET
--		<cky@photox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 2001

class CompositeShapeAspect  from StepRepr    inherits ShapeAspect from StepRepr

    ---Purpose : Added for Dimensional Tolerances

uses
    Integer

is

    Create returns mutable CompositeShapeAspect;

end CompositeShapeAspect;
