-- Created on: 1996-12-17
-- Created by: Yves FRICAUD
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



private class RefShape from TNaming 

uses
   Label       from TDF,
   NamedShape  from TNaming, 	
   Shape       from TopoDS,
   PtrNode     from TNaming     

is
    Create returns RefShape from TNaming;
	---C++: inline    
    
    Create (S : Shape from TopoDS) returns RefShape from TNaming;
	---C++: inline    
    
    Shape    (me : in out; S    : Shape    from TopoDS);
    	---C++: inline
    
    FirstUse (me : in out; aPtr : PtrNode from TNaming);
	---C++: inline

    ---Category: Querying

    FirstUse (me) returns PtrNode from TNaming;
	---C++: inline    
    
    Shape (me) returns Shape    from TopoDS;
	---C++: return const&
    	---C++: inline

    Label (me) returns Label from TDF;
    
    NamedShape (me) returns NamedShape from TNaming;

	    
fields

    myShape      : Shape    from TopoDS;
    myFirstUse   : PtrNode  from TNaming;	

end RefShape;
