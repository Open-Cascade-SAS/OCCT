-- Created on: 1993-12-02
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




generic class PointOnRst from Blend
    (TheArc    as any)


	---Purpose: Definition of an intersection point between a line
	--          and a restriction on a surface.
	--          Such a point is contains geometrical informations (see
	--          the Value method) and logical informations.


uses Transition from IntSurf
     
raises DomainError from Standard

is


    Create
    
	---Purpose: Empty constructor.

    	returns PointOnRst from Blend;


    Create( A: TheArc; Param: Real from Standard;
            TLine, TArc: Transition from IntSurf)

	---Purpose: Creates the PointOnRst on the arc A, at parameter Param,
	--          with the transition TLine on the walking line, and
	--          TArc on the arc A.

    	returns PointOnRst from Blend;



    SetArc(me: in out; A: TheArc; Param: Real from Standard;
                       TLine, TArc: Transition from IntSurf)

	---Purpose: Sets the values of a point which is on the arc
	--          A, at parameter Param.


    	is static;



    Arc(me)
    
	---Purpose: Returns the arc of restriction containing the
	--          vertex.

    	returns any TheArc
	---C++: return const&
	---C++: inline
	
	is static;


    TransitionOnLine(me)
    
	---Purpose: Returns the transition of the point on the
	--          line on surface.

    	returns Transition from IntSurf
	---C++: return const&
	---C++: inline
	
	is static;


    TransitionOnArc(me)
    
	---Purpose: Returns the transition of the point on the arc
	--          returned by Arc().

    	returns Transition from IntSurf
	---C++: return const&
	---C++: inline
	
	is static;


    ParameterOnArc(me)
    
	---Purpose: Returns the parameter of the point on the
	--          arc returned by the method Arc().

    	returns Real from Standard
	---C++: inline
	
	is static;


fields

    arc       : TheArc;
    traline   : Transition from IntSurf;
    traarc    : Transition from IntSurf;
    prm       : Real       from Standard;

end PointOnRst;
