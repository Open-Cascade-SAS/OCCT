-- Created on: 1993-11-10
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class WPointInter from TopOpeBRep 

  -- as WPointTool from TopOpeLine
  -- 	 (PntOn2S from IntSurf)
  -- 	 

	---Purpose: 

uses

  PntOn2S from IntSurf,
  PPntOn2S from TopOpeBRep,
  Pnt2d from gp,
  Pnt from gp
  
is

  Create returns WPointInter from TopOpeBRep;
  
  Set(me : in out; P : PntOn2S from IntSurf) is static;

  ParametersOnS1(me; U,V : out Real from Standard) is static;
		  
  ParametersOnS2(me; U,V : out Real from Standard) is static;
		  
  Parameters(me; U1,V1,U2,V2 : out Real from Standard) is static;
	    
  ValueOnS1(me) returns Pnt2d from gp is static;
	
  ValueOnS2(me) returns Pnt2d from gp is static;
	
  Value(me) returns Pnt from gp is static;
   ---C++: return const &

  PPntOn2SDummy(me) returns PPntOn2S from TopOpeBRep;

fields

    myPP2S : PPntOn2S from TopOpeBRep;

end WPointInter;
