-- Created on: 1992-08-27
-- Created by: Christophe MARION
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DrawablePolyEdgeTool from HLRTest inherits Drawable3D from Draw

	---Purpose: Used to display the results.

uses
    Boolean      from Standard,
    Integer      from Standard,
    Display      from Draw,
    PolyAlgo     from HLRBRep,
    ListOfBPoint from HLRBRep

is
    Create(Alg    : PolyAlgo from HLRBRep;
           ViewId : Integer  from Standard;
           Debug  : Boolean  from Standard = Standard_False)
    returns DrawablePolyEdgeTool from HLRTest;
    
    Show(me : mutable)
    	---C++: inline
    is static;

    Hide(me : mutable)
    	---C++: inline
    is static;

    DisplayRg1Line(me : mutable; B : Boolean from Standard)
	---C++: inline
    is static;
    
    DisplayRg1Line(me) returns Boolean from Standard
	---C++: inline
    is static;
    
    DisplayRgNLine(me : mutable; B : Boolean from Standard)
	---C++: inline
    is static;
    
    DisplayRgNLine(me) returns Boolean from Standard
	---C++: inline
    is static;
    
    DisplayHidden(me : mutable; B : Boolean from Standard)
	---C++: inline
    is static;
    
    DisplayHidden(me) returns Boolean from Standard
	---C++: inline
    is static;
    
    DrawOn(me; D : in out Display from Draw);
    
    Debug(me) returns Boolean from Standard
	---C++: inline
    is static;
    
    Debug(me : mutable; B : Boolean from Standard)
	---C++: inline
    is static;
    
fields
    myAlgo     : PolyAlgo     from HLRBRep;
    myDispRg1  : Boolean      from Standard;
    myDispRgN  : Boolean      from Standard;
    myDispHid  : Boolean      from Standard;
    myViewId   : Integer      from Standard;
    myBiPntVis : ListOfBPoint from HLRBRep;
    myBiPntHid : ListOfBPoint from HLRBRep;
    myDebug    : Boolean      from Standard;
    myHideMode : Boolean      from Standard;

end DrawablePolyEdgeTool;
