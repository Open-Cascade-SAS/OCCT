-- Created on: 1993-06-17
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package TopOpeBRepBuild 

---Purpose: 
--  This package describes algorithms and dedicated tools
--  involved in topological operation on BRep shapes.
--  These "builders" works on a data structure that must have been
--  previously filled (by a "filler") according to the
--  topological operation rules defined in class DataStructure
--  from TopOpeBRepDS.
--  The DSFiller must be considered as a "linking" tool
--  dealing with geometric data as an input and a DS as an
--  output.
--  These geometric data may be seen as the result of 3D 
--  intersection between BRep shapes.

uses

    Standard, MMgt, TCollection, TColStd, 
    gp, Geom, Geom2d, Geom2dInt,
    TopAbs, TopoDS, TopTools, TopExp,
    BRepClass, BRep,
    TopOpeBRepDS, TopOpeBRepTool,  
    --modified by NIZNHY-PKV Thu Feb 10 11:51:54 2000  f
    Bnd 
    --modified by NIZNHY-PKV Thu Feb 10 11:51:57 2000  t
    
is
    
    class Loop;
    imported ListOfLoop;
    imported ListIteratorOfListOfLoop;
    class LoopSet;
    deferred class LoopClassifier;
    enumeration LoopEnum is ANYLOOP,BOUNDARY,BLOCK end LoopEnum;
    imported ListOfListOfLoop;
    imported ListIteratorOfListOfListOfLoop;
    class AreaBuilder;

    class Pave;
    imported ListOfPave;
    imported ListIteratorOfListOfPave;
    class PaveSet;
    class PaveClassifier;
    class Area1dBuilder;
    class EdgeBuilder;

    --modified by NIZHNY-MZV  Mon Sep 20 15:43:24 1999 
    class  Tools;
--    class  LoopTreeNode; 
--    class  ListOfLoopTreeNode  instantiates  List  from  TCollection  (LoopTreeNode); 
--    class  IndexedDataMapOfLoopListOfLoop  instantiates  IndexedDataMap  from  TCollection 
--    (Transient  from  Standard,  ListOfLoop  from  TopOpeBRepBuild,  MapTransientHasher  from  TColStd);


    class ShapeSet;
    class WireEdgeSet;pointer PWireEdgeSet to WireEdgeSet from TopOpeBRepBuild;
    class ShellFaceSet;

    class BlockIterator;
    class BlockBuilder;

    deferred class CompositeClassifier;
    class WireEdgeClassifier;
    class ShellFaceClassifier;

    class Area2dBuilder;
    class FaceAreaBuilder;
    class FaceBuilder;

    class Area3dBuilder;
    class SolidAreaBuilder;
    class SolidBuilder;
    
    class ShapeListOfShape;
    imported ListOfShapeListOfShape;
    imported ListIteratorOfListOfShapeListOfShape;
    imported DataMapOfShapeListOfShapeListOfShape;
    imported DataMapIteratorOfDataMapOfShapeListOfShapeListOfShape;

    class GTopo; pointer PGTopo to GTopo from TopOpeBRepBuild;
    class GIter;
    class GTool;
    
    class Builder; pointer PBuilder to Builder from TopOpeBRepBuild;  
    --modified by NIZHNY-MZV  Wed Sep 29 09:33:20 1999
    class Builder1;
    class BuilderON;
    
    class HBuilder;
    class WireToFace;
    class ShellToSolid;
    class FuseFace;

--modified by NIZNHY-PKV Thu Feb 10 11:25:15 2000  from 
    class  CorrectFace2d; 
    class  VertexInfo; 
    class  Tools2d;	     
    imported IndexedDataMapOfShapeVertexInfo;  
   		 
--modified by NIZNHY-PKV Thu Feb 10 11:25:19 2000  to

end TopOpeBRepBuild;
