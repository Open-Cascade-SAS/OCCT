-- Created on: 2002-12-12
-- Created by: data exchange team
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class NodeGroup from StepFEA
inherits FeaGroup from StepFEA

    ---Purpose: Representation of STEP entity NodeGroup

uses
    HAsciiString from TCollection,
    FeaModel from StepFEA,
    HArray1OfNodeRepresentation from StepFEA

is
    Create returns NodeGroup from StepFEA;
	---Purpose: Empty constructor

    Init (me: mutable; aGroup_Name: HAsciiString from TCollection;
                       aGroup_Description: HAsciiString from TCollection;
                       aFeaGroup_ModelRef: FeaModel from StepFEA;
                       aNodes: HArray1OfNodeRepresentation from StepFEA);
	---Purpose: Initialize all fields (own and inherited)

    Nodes (me) returns HArray1OfNodeRepresentation from StepFEA;
	---Purpose: Returns field Nodes
    SetNodes (me: mutable; Nodes: HArray1OfNodeRepresentation from StepFEA);
	---Purpose: Set field Nodes

fields
    theNodes: HArray1OfNodeRepresentation from StepFEA;

end NodeGroup;
