-- Created on: 1996-12-16
-- Created by: Christian CAILLET
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class SelectNamed  from StepData    inherits SelectMember

    ---Purpose : This select member can be of any kind, and be named
    --           But its takes more memory than some specialised ones
    --           This class allows one name for the instance

uses CString, Logical, AsciiString from TCollection,  Field from StepData

is

    Create  returns mutable SelectNamed;

    HasName (me) returns Boolean  is redefined;

    Name (me) returns CString  is redefined;

    SetName (me : mutable; name : CString)  returns Boolean  is redefined;
    -- redefined to accept any name

    Field (me) returns Field;
    ---C++ : return const &

    CField (me : mutable) returns Field;
    ---C++ : return &


    Kind (me) returns Integer  is redefined;
    --  see Field for Kind (same codes)

    SetKind  (me : mutable; kind : Integer)  is redefined;
    --  called by various Set*

    Int (me) returns Integer  is redefined;
    ---Purpose : This internal method gives access to a value implemented by an
    --           Integer (to read it)

    SetInt (me : mutable; val : Integer)  is redefined;
    ---Purpose : This internal method gives access to a value implemented by an
    --           Integer (to set it)

    Real (me) returns Real  is redefined;

    SetReal (me : mutable; val : Real)  is redefined;

    String (me) returns CString  is redefined;

    SetString (me : mutable; val : CString)  is redefined;

fields

    thename : AsciiString;
    theval  : Field from StepData;

end SelectNamed;
