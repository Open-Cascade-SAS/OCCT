-- Created on: 1998-07-31
-- Created by: Christian CAILLET
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SignTransferStatus  from XSControl    inherits Signature  from IFSelect

    ---Purpose : This Signatures gives the Transfer Status of an entity, as
    --           recorded in a TransferProcess. It can be :
    --           - Void : not recorded, or recorded as void with no message
    --             (attributes are not taken into account)
    --           - Warning : no result, warning message(s), no fail
    --           - Fail : no result, fail messages (with or without warning)
    --           - Result.. : result, no message (neither warning nor fail)
    --             Result.. i.e. Result:TypeName of the result
    --           - Result../Warning : result, with warning but no fail
    --           - Result../Fail : result, with fail (.e. bad result)
    --           - Fail on run : no result yet recorded, no message, but
    --             an exception occurred while recording the result
    --             (this should not appear and indicates a programming error)

uses CString, Transient, InterfaceModel,
     TransientProcess, TransferReader

is

    Create returns mutable SignTransferStatus;
    ---Purpose : Creates a SignTransferStatus, not initialised
    --           it gives nothing (empty string)

    Create (TR : TransferReader) returns mutable SignTransferStatus;
    ---Purpose : Creates a SignTransferStatus, which will work on the current
    --           TransientProcess brought by the TransferReader (its MapReader)

    SetReader (me : mutable; TR : TransferReader);
    ---Purpose : Sets a TransferReader to work

    SetMap (me : mutable; TP : TransientProcess);
    ---Purpose : Sets a precise map to sign entities
    --           This definition oversedes the creation with a TransferReader

    Map    (me) returns TransientProcess;
    ---Purpose : Returns the TransientProcess used as precised one
    --           Returns a Null Handle for a creation from a TransferReader
    --           without any further setting

    Reader (me) returns TransferReader;
    ---Purpose : Returns the Reader (if created with a Reader)
    --           Returns a Null Handle if not created with a Reader


    Value (me; ent : any Transient; model : InterfaceModel) returns CString;
    ---Purpose : Returns the Signature for a Transient object, as its transfer
    --           status

fields
 
    theTR : TransferReader;
    theTP : TransientProcess;
 
end SignTransferStatus;
