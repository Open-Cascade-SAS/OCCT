-- Created on: 1993-06-03
-- Created by: Bruno DUMORTIER
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package Geom2dAdaptor 

	---Purpose: this package  contains the geometric definition of
	--          2d  curves compatible  with  the  Adaptor  package
	--          templates.

uses
    Geom2d,
    GeomAbs,
    Adaptor2d,
    gp,
    Standard,
    TColStd,
    TColgp

is

 
      class Curve; 

      private class GHCurve instantiates GenHCurve2d from Adaptor2d
    	    (Curve from Geom2dAdaptor);

      class HCurve;
	---Purpose: Inherited  from    GHCurve.   Provides a  curve
	--          handled by reference.

      --
      --   Package methods
      --   
      
      MakeCurve(HC : Curve2d from Adaptor2d) returns Curve from Geom2d
	    ---Purpose: Creates  a 2d  curve  from  a  HCurve2d.  This
	    --          cannot process the OtherCurves.
      raises
      	DomainError from Standard; -- if GeomAbs_OtherCurve

end Geom2dAdaptor;



