-- Created on: 2000-05-25
-- Created by: Peter KURNEV
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class DrawableShape from BOPTest inherits DrawableShape from DBRep

    ---Purpose: 

uses  

    Shape           from TopoDS,
    Color           from Draw,
    Display         from Draw,
    Text3D          from Draw,
    Marker3D        from Draw,
    CString         from Standard,
    Pnt             from gp

is

    Create (S         : Shape from TopoDS;
    	    FreeCol   : Color from Draw;    -- color for free edges
    	    ConnCol   : Color from Draw;    -- color for shared edges
	    EdgeCol   : Color from Draw;    -- color for other edges
	    IsosCol   : Color from Draw;    -- color for Isos
	    size      : Real;               -- size for infinite isos
	    nbisos    : Integer;            -- # of isos on each face
	    discret   : Integer;            -- # of points on curves
    	    Text      : CString from Standard; 
    	    TextColor : Color from Draw
    	    )
    	returns mutable DrawableShape from BOPTest;

    Create (S         : Shape from TopoDS;
    	    Text      : CString from Standard; 
    	    TextColor : Color from Draw
    	    )
    	returns mutable DrawableShape from BOPTest; 
	
    Pnt(me) returns Pnt from gp  is private;
  
    DrawOn(me; dis : in out Display from Draw)
    is redefined;
    
fields

    myText : Text3D from Draw;
    myTextColor : Color from Draw;

end DrawableShape;
