-- Created by: Tanya COOL
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Drawer from Prs2d inherits TShared from MMgt

  --- Purpose: Graphic attributes management
  --           Qualifies how the presentation algorithms compute
  --           the presentation of a specific kind of object. 
  --           This includes for example color, width and type
  --           of lines...

uses

    NameOfColor         from Quantity,
    TypeOf2DObject      from Prs2d,
    AspectRoot          from Prs2d,
    AspectName          from Prs2d,
    DataMapOfAspectRoot from Prs2d
    
is
    Create returns mutable Drawer from Prs2d;
    ---Purpose: Initializes graphic attribute manager

    FindAspect( me; anAspectName: AspectName from Prs2d )
      returns AspectRoot from Prs2d is virtual;
    ---Level: Public
    ---Purpose: Returns a link with Prs2d_Drawer AspectName, 
    --          which provides settings for object "anAspectName" 
    --          used to display "anAspectName"
  	
    SetAspect( me: mutable;
               anAspectRoot: AspectRoot from Prs2d;
               anAspectName: AspectName from Prs2d );
    ---Level: Public
    ---Purpose: Sets the Aspect <anAspectRoot> of the Drawer
    
    InitAspectRootMap( me: mutable ) is private;
    ---Level: Internal
    ---Purpose: Initializes Aspect classes data map

   --******************************************************

    SetMaxParameterValue( me: mutable; Value: Real from Standard ) is virtual;
    ---Level: Public
    ---Purpose: defines the maximum value allowed for the first and last
    --          parameters of an infinite line.
    --          Default value: 500000. 
    
    MaxParameterValue( me ) returns Real from Standard is virtual;
    ---Level: Public
    ---Purpose: Indicates the maximum value allowed for the first and last
    --          parameters of an infinite line.


fields

    myDataMapAspectRoot: DataMapOfAspectRoot from Prs2d is protected;
    myMaxParameterValue: Real from Standard is protected;
   
end Drawer;
