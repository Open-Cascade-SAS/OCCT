-- File:	RWStepRepr_RWMakeFromUsageOption.cdl
-- Created:	Mon Jul  3 20:13:36 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class RWMakeFromUsageOption from RWStepRepr

    ---Purpose: Read & Write tool for MakeFromUsageOption

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    MakeFromUsageOption from StepRepr

is
    Create returns RWMakeFromUsageOption from RWStepRepr;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : MakeFromUsageOption from StepRepr);
	---Purpose: Reads MakeFromUsageOption

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: MakeFromUsageOption from StepRepr);
	---Purpose: Writes MakeFromUsageOption

    Share (me; ent : MakeFromUsageOption from StepRepr;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWMakeFromUsageOption;
