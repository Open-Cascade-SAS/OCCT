
-- File:	MFT_FontManager.cdl
-- Created:	Tue Mar 3 09:14:42 1997
-- Author:	Gerard GRAS
--		<gg@photox>
---Copyright:	 Matra Datavision 1993

class FontManager from MFT inherits TShared from MMgt

        ---Purpose: This class permits to manage MDTV fonts.
	--  Warning: A FontManager is associated to a xxx.mft font file 
	-- 	    The coordinates of the outline vectors of each character
	-- 	    must be given in the space defined by the font bounding box


uses

	TextManager		from MFT,
	TypeOfCommand		from MFT,
        TypeOfValue 		from MFT,
	CommandDescriptor	from MFT,
	FileRecord		from MFT,
	FileHandle		from MFT,
	FilePosition		from MFT,
	FontStyle		from Aspect,
	AsciiString		from TCollection,
	Length			from Quantity,
	Factor			from Quantity,
	PlaneAngle		from Quantity,
	OpenMode 		from OSD

raises

	FontManagerDefinitionError	from MFT,
	FontManagerError		from MFT,
	OutOfRange			from Standard,
	OutOfMemory			from Standard,
	TypeMismatch			from Standard

is

	-------------------------
	-- Category: Constructors
	-------------------------

	Create (anAliasName: CString from Standard)
	returns mutable FontManager from MFT
	---Level: Public
	---Purpose: Gives access to the font <anAliasName> associated
	--	    to the file $CSF_MDTVFontDirectory/<anAliasName>.mft  
	--	    in ReadOnly access mode.
	--  Warning: If the symbol CSF_MDTVFontDirectory is not defined
	--	    try to reads or writes in $PWD directory.
	--  Example: myFontManager = new MFT_FontManager("Helvetica-Bold")
	--	    permits to access to the file 
	--	    $CSF_MDTVFontDirectory/"helvetica-bold.mft" 
	--  Trigger: If the font file don't exist or if the file 
	--	    don't have an MFT signature.

	raises FontManagerDefinitionError from MFT;

	Create (aFont: FontStyle from Aspect;
		aFileMode: OpenMode from OSD = OSD_ReadOnly;
		isComposite: Boolean from Standard = Standard_False)
	returns mutable FontManager from MFT
	---Level: Public
	---Purpose: Gives access to the font <aFont> associated
	--	    to the file $CSF_MDTVFontDirectory/<aFont.AliasName()>.mft  
	--	    with the open mode <aFileMode> and the composite
	--	    flag <isComposite>.
	--  Example: The flag must be sets to TRUE for KANJI extended fonts.
	--  Warning: If the symbol CSF_MDTVFontDirectory is not defined
	--	    try to reads or writes in $PWD directory.	 
--  Trigger: If <aFileMode> is ReadOnly or ReadWrite and
	--	    the font file don't exist or if the file 
	--	    don't have an MFT signature.

	raises FontManagerDefinitionError from MFT;

	-------------------------
	-- Category: Destructors
	-------------------------

        Destroy ( me : mutable);
        ---Level: Internal
        ---Purpose: Save the font file when the open mode is
	--	   Write or ReadWrite and Close it in all the case.
        ---C++: alias ~

	---------------------------------------------
	-- Category: Methods to updates the .mft files
	---------------------------------------------

	SetFont (me : mutable;
		aFont: FontStyle from Aspect)
	---Level: Advanced
	---Purpose: Updates the font name. 
	--  Trigger: If the font file is not opened
	--	    in WriteOnly or ReadWrite mode
		
	raises FontManagerError from MFT;

	SetChar (me: mutable;
		aChar: Character from Standard)
	---Level: Advanced
	---Purpose: Defines and Enable the char <aChar> for writing.	 
--  Trigger: If the font file is not opened
	--	    in WriteOnly or ReadWrite mode
	--	    or the char is already defined.
	raises FontManagerError from MFT;


	SetAccentChar (me: mutable;
		aChar: Character from Standard)
	---Level: Advanced
	---Purpose: Defines and Enable the accent char <aChar> for writing.	 
--  Trigger: If the font file is not opened
	--	    in WriteOnly or ReadWrite mode
	--	    or the char is already defined.

	raises FontManagerError from MFT;

	SetChar (me: mutable;
		aChar: ExtCharacter from Standard)
	---Level: Advanced
	---Purpose: Defines and Enable the char <aChar> for writing.
	--	    This char being current for adding command.
	--  Warning: The char must have an UNICODE UCS2 encoding. 
	--  Trigger: If the font file is not opened
	--	    in WriteOnly or ReadWrite mode
	--	    or if the font is not a composite font.

	raises FontManagerError from MFT;

	SetEncoding (me: mutable;
		aPosition: Integer from Standard;
		anEncoding: CString from Standard)
	---Purpose: Changes the default encoding of the char position
	--	   <aPosition>.
        --  Example: SetEncoding(233,"eacute")
	--	   change the default encoding of the char position 233
	--	   from "Oslash" to "eacute". 
	raises FontManagerError from MFT;
	---Purpose:  Trigger  - If the font file is not opened
	--	    in WriteOnly or ReadWrite mode.
	--	    or if the char encoding is not defined.

	DelChar (me: mutable;
		aChar: Character from Standard)
	---Level: Advanced
	---Purpose: Remove the definition of the char <aChar>
	raises FontManagerError from MFT;
	---Purpose:  Trigger  - If the font file is not opened
	--	    in WriteOnly or ReadWrite mode.

	DelChar (me: mutable;
		aChar: ExtCharacter from Standard)
	---Level: Advanced
	---Purpose: Remove the definition of the char <aChar>
	--	    This char being current for adding command.
	--Warning: The char must have an UNICODE UCS2 encoding.
	raises FontManagerError from MFT;
	---Purpose:  Trigger  - If the font file is not opened
	--	    in WriteOnly or ReadWrite mode
	--	    or if the font is not a composite font.

	AddCommand (me : mutable;
		aCommand: TypeOfCommand from MFT)
	---Level: Advanced
	---Purpose: Adds the command <aCommand> of <aNumberOfValues>
	--	    to describe the current char.
	--	    This command being current for adding parameters if any.
	raises FontManagerError from MFT;
	---Purpose  Trigger - If the font file is not opened
	--	    in WriteOnly or ReadWrite mode
	--	    or if a current char don't have being defined.
	--  Warning: the last command of the char descriptor
	--	   must have a type MFC_TOC_ENDCHAR.

	AddValue (me : mutable;
		aValue: Integer from Standard)
	---Level: Advanced
	---Purpose: Adds the integer parameter <aValue> to fill
	--	    the current command.
	raises FontManagerError from MFT;
	---Purpose:  Trigger - If the font file is not opened
	--	    in WriteOnly or ReadWrite mode
	--	    or if a current command don't have being defined,
	--	    or if the number of values is > MaxCommandValues()

	AddValue (me : mutable;
		aValue: Real from Standard)
	---Level: Advanced
	---Purpose: Adds the float parameter <aValue> to fill
	--	    the current command.
	raises FontManagerError from MFT;
	---Purpose:  Trigger - If the font file is not opened
	--	    in WriteOnly or ReadWrite mode
	--	    or if a current command don't have being defined
	--	    or if the number of values is > MaxCommandValues()

	AddValue (me : mutable;
		aValue: CString from Standard)
	---Level: Advanced
	---Purpose: Adds the string parameter <aValue> to fill
	--	    the current command.
	raises FontManagerError from MFT;
	---Purpose:  Trigger - If the font file is not opened
	--	    in WriteOnly or ReadWrite mode
	--	    or if a current command don't have being defined,
	--	    or if the number of values is > MaxCommandValues()
	--  Warning: The max length of a string must be < MaxCommandValues()*4-1

	SetBoundingBox (me : mutable;
		aMinX: Integer from Standard = 0;
		aMinY: Integer from Standard = 0;
		aMaxX: Integer from Standard = 1000;
		aMaxY: Integer from Standard = 1000)
	---Level: Advanced
	---Purpose: Sets the bounding box of the font. 
	raises FontManagerError from MFT;
	---Purpose:  Trigger - If the font file is not opened
	--	    in WriteOnly or ReadWrite mode
	--	    or if the bounding box has a wrong value.
	--  Warning: The bounding box coordinates default are :
	--	    0,0,1000,1000 

	SetFontMatrix (me : mutable;
		M1: Real from Standard = 0.001;
		M2: Real from Standard = 0.0;
		M3: Real from Standard = 0.0;
		M4: Real from Standard = 0.001;
		M5: Real from Standard = 0.0;
		M6: Real from Standard = 0.0)
	---Level: Advanced
	---Purpose: Sets the font matrix. 
	raises FontManagerError from MFT;
	---Purpose:  Trigger - If the font file is not opened
	--	    in WriteOnly or ReadWrite mode
	--  Warning: The font matrix default are :
	--	    0.001,0,0,0.001,0,0 

	SetPaintType (me : mutable;
		aValue: Integer from Standard = 0)
	---Level: Advanced
	---Purpose: Sets the paint type of the font. 
	raises FontManagerError from MFT;
	---Purpose:  Trigger - If the font file is not opened
	--	    in WriteOnly or ReadWrite mode
	--	    or if the value is not a Type 1 font value.
	--  Warning: The paint type <aValue> must be one of Type 1 font
	--	   value 0 for FILL , 1 for STROKE or 2 for OUTLINE.

	SetFixedPitch (me : mutable;
		aFlag: Boolean from Standard = Standard_False)
	---Level: Advanced
	---Purpose: Sets the fixed pitch flag of the font
	--  as TRUE if the font must have an fixed char width 
	--  or FALSE if the font must have a proportionnal char width.
	raises FontManagerError from MFT;
	---Purpose:  Trigger - If the font file is not opened
	--	    in WriteOnly or ReadWrite mode

	SetItalicAngle (me : mutable;
		anAngle: PlaneAngle from Quantity = 0.0)
	---Level: Advanced
	---Purpose: Sets the italic angle of the font given in RAD
	--		clock-wise from vertical.
	raises FontManagerError from MFT;
	---Purpose:    Trigger - If the font file is not opened
	--	    in WriteOnly or ReadWrite mode

	ComputeBoundingBox (me: mutable)
	---Level: Advanced
	---Purpose: Computes the bounding box of the font from the
	--	    min-max of all chars of the font. 
	--  Warning: this must be call after all characters has been defined.
	raises FontManagerError from MFT;
	---Purpose:  Trigger - If the font file is not opened
	--	    in WriteOnly or ReadWrite mode.

	---------------------------------------------------------------
	-- Category: Methods to sets the current interpretor attributes 
	---------------------------------------------------------------

	SetFontAttribs (me: mutable;
		aWidth,aHeight: Length from Quantity;
		aSlant: PlaneAngle from Quantity = 0.0;
		aPrecision: Factor from Quantity = 0.02;
		aCapsHeight: Boolean from Standard = Standard_False);
	---Level: Public
	---Purpose: Sets the current font attributes.
	--  <aWidth> : the maximum width of one character.
	--  <aHeight> : the maximum height of one character
	--		according to the <aCapsHeight> parameter.
	--  <aSlant> : the slant of one character given in RAD
	--		clock-wise from vertical.
	--  <aPrecision> : the relative interpolator precision is
	--	the maximum flatness error deflection for the curves.
	--  <aCapsHeight> : if TRUE the font height is apply only
	--  	        on the ascent component of the characters;
	--		    if FALSE the font height is apply both
	--		on the ascent and descent  components of the characters.

	----------------------------------------------------------------
	-- Category: Methods to retrieve current attributes informations. 
	----------------------------------------------------------------

	DrawText (me: mutable;
		aTextManager: TextManager from MFT;
		aString: CString from Standard;
		anX,anY: Length from Quantity;
		anOrientation: PlaneAngle from Quantity = 0.0);
	---Level: Public
	---Purpose: Drawn an ANSI text 
	--  <aTextManager> : the draw manager to call for each vertex of the string.
	--  <aString> : the string to interpret 
	--  <anX>,<anY> : the position of the text
	--  <anOrientation> : the orientation angle in RAD from horizontal. 

	DrawText (me: mutable;
		aTextManager: TextManager from MFT;
		aString: ExtString from Standard;
		anX,anY: Length from Quantity;
		anOrientation: PlaneAngle from Quantity = 0.0)
	---Level: Public
	---Purpose: Drawn an EXTENDED text 
	--  <aTextManager> : the draw manager to call for each vertex of the string.
	--  <aString> : the string to interpret 
	--  <anX>,<anY> : the position of the text
	--  <anOrientation> : the orientation angle in RAD from horizontal. 
	raises FontManagerError from MFT;
	---Purpose:  Trigger - If the font is not a composite font and
	--	   the string is not ASCII.

	BoundingBox (me ;
		aMinX,aMinY,aMaxX,aMaxY: out Integer from Standard);
	---Level: Advanced
	---Purpose: Retrieves the bounding box of the font. 

	CharBoundingBox (me : mutable ;
		aPosition: Integer from Standard;
		aMinX,aMinY,aMaxX,aMaxY: out Integer from Standard)
	---Level: Advanced
	---Purpose: Retrieves the bounding box of a character. 
	raises FontManagerError from MFT;
	---Purpose:  Trigger - If the position <aPosition> is < 0 or > MaxCharPosition(). 

	PaintType (me)
		returns Integer from Standard;
	---Level: Advanced
	---Purpose: Retrieves the paint type of the font. 

	FixedPitch (me)
		returns Boolean from Standard;
	---Level: Advanced
	---Purpose: Retrieves the fixed pitch flag of the font

	ItalicAngle (me)
		returns PlaneAngle from Quantity;
	---Level: Advanced
	---Purpose: Retrieves the italic angle of the font

	FontAttribs (me : mutable;
		aWidth,aHeight,aDescent: out Length from Quantity;
		aSlant: out PlaneAngle from Quantity;
		aPrecision: out Factor from Quantity;
		aCapsHeight: out Boolean from Standard)
		returns CString from Standard;
	---Level: Public
	---Purpose: Runs the interpretor with the current attributes setting
	--	   (font and text attributes)
	--	   and returns :
	--	   The max char width of the font CharSet <aWidth>.
	--	   The max char height of the font CharSet <aHeight>.
	--	   The max char descent value below the baseline <aDescent>
	--	   The slant angle of the font <aSlant>
	--	   The interpolator precision of the font <aPrecision>
	--  	   The caps height flag <aCapsHeight>
	--	   The FULL font name.

	TextSize (me : mutable;
		aString: CString from Standard;
		aWidth,anAscent,aLbearing,aDescent: out Length from Quantity);
	---Level: Public
	---Purpose: Runs the interpretor on the ASCII text <aString> 
	--	   with the current font attributes setting and returns :
	--	   The string width <aWidth>.
	--	   The string ascent <anAscent>.
	--	   The string left bearing value from the origine <aLbearing>
	--	   The string descent value below the baseline <aDescent>

	TextSize (me : mutable;
		aString: ExtString from Standard;
		aWidth,anAscent,aLbearing,aDescent: out Length from Quantity)
	---Level: Public
	---Purpose: Runs the interpretor on the EXTENDED text <aString> 
	--	   with the current font attributes setting and returns :
	--	   The string width <aWidth>.
	--	   The string ascent <anAscent>.
	--	   The string left bearing value from the origine <aLbearing>
	--	   The string descent value below the baseline <aDescent>
	raises FontManagerError from MFT;
	---Purpose:  Trigger - If the font is not a composite font and
	--	   the string is not ASCII.

	CharSize (me : mutable;
		aChar: Character from Standard;
		aWidth,aLbearing,aRbearing: out Length from Quantity;
		anAscent,aDescent: out Length from Quantity)
		returns Boolean from Standard;
	---Level: Public
	---Purpose: Runs the interpretor with the current attributes setting
	--	   (font attributes)
	--	   and returns :
	--	   The char width <aWidth>.
	--	   The char left bearing <aLbearing>.
	--	   The char right bearing <aRbearing>.
	--	   The char ascent <anAscent>.
	--	   The char descent value below the baseline <aDescent>
	--	And returns TRUE if the character is defined.

	CharSize (me : mutable;
		aChar: ExtCharacter from Standard;
		aWidth,aLbearing,aRbearing: out Length from Quantity;
		anAscent,aDescent: out Length from Quantity)
		returns Boolean from Standard
	---Level: Public
	---Purpose: Runs the interpretor with the current attributes setting
	--	   (font attributes)
	--	   and returns :
	--	   The extended char width <aWidth>.
	--	   The extended char left bearing <aLbearing>.
	--	   The extended char right bearing <aRbearing>.
	--	   The extended char ascent <anAscent>.
	--	   The extended char descent value below the baseline <aDescent>
	--	And returns TRUE if the character is defined.
	raises FontManagerError from MFT;
	---Purpose:  Trigger - If the font is not a composite font and
	--	   the char is not ASCII.

	----------------------------
	-- Category: Inquire methods
	----------------------------

	Font (me)
		returns FontStyle from Aspect;
	---Level: Public
	---Purpose: Retrieves the font descriptor of this font

        IsComposite (me)
                returns Boolean from Standard;
        ---Level: Public
        ---Purpose: Returns TRUE if the font is composite.
        --  Example: KANJI fonts returns TRUE.

	IsKnown (myclass;
		anAliasName: CString from Standard)
		returns Boolean from Standard;
	---Purpose: Returns TRUE if the font
	--	    $CSF_MDTVFontDirectory/<anAliasName>.mft does exist.

	Font (myclass;
		anAliasName: CString from Standard)
		returns FontStyle from Aspect
	---Level: Public
	---Purpose: Retrieves the font descriptor from an existing font
	raises FontManagerError from MFT;
	---Purpose: Trigger - If the font does not exist.

	FontNumber (myclass;
		aFilter: CString from Standard = "*")
		returns Integer from Standard;
	---Level: Public
	---Purpose: Returns the MFT font number available
	--	    in the directory $CSF_MDTVFontDirectory
	--	    according to the filter :
        -- "-foundry-family-weight-slant-swidth-adstyl-pixelsize-pointsize-
        --  resx-resy-spacing-avdWidth-registry-encoding"
	--  Examples: number = MFT_FontMAnager::FontNumber("-euclid3");
	--	    returns only the euclid3 fonts.
	--          number = MFT_FontMAnager::FontNumber(
	--			"-*-*-*-*-*-*-*-*-*-*-*-*-japanese");
	--	    returns only the japanese fonts.

	Font (myclass;
		aRank: Integer from Standard)
		returns FontStyle from Aspect
	---Level: Public
	---Purpose: Retrieves the font descriptor of index <aRank>
	--	   from the directory $CSF_MDTVFontDirectory
	raises OutOfRange from Standard;
	---Purpose:  Trigger - If the font rank <aRank> is < 1 or > FontNumber().

	MaxCommandValues (myclass)
		returns Integer from Standard;
	---Purpose: Returns the max values of any defined command

	Encoding (me: mutable;
		aPosition: Integer from Standard)
		returns CString from Standard
	---Purpose: Returns the encoding of the char position
	--	   <aPosition>.
	raises FontManagerError from MFT;
	---Purpose:  Trigger -  If the char is not defined

	Encoding (me: mutable;
		anEncoding: CString from Standard)
		returns Integer from Standard
	---Purpose: Returns the char position
	--	   from the encoding <anEncoding>.
	raises FontManagerError from MFT;
	---Purpose:  Trigger - If the char is not defined

	Dump (me : mutable);
	---Level: Public
	---Purpose: Dumps the font descriptor of all characters.

	Dump (me : mutable; aChar: Character from Standard);
	---Level: Public
	---Purpose: Dumps the font descriptor of the character <aChar>.

	Dump (me : mutable; aChar: ExtCharacter from Standard)
	---Level: Public
	---Purpose: Dumps the font descriptor of the extended character <aChar>.
	raises FontManagerError from MFT;
	---Purpose:  Trigger - If the font is not a composite font.

	Save (me : mutable) returns Boolean from Standard;
	---Level: Public
	---Purpose: Saves the entire MFT font in an ASCII format
	--	    readable by the Restore() method. 
	--	    to the file $CSF_MDTVFontDirectory/<anAliasName>.dat  
	--	    And returns TRUE if the file have been saves correctly.

	Restore (myclass; anAliasName: CString from Standard) returns Boolean from Standard;
	---Level: Public 
	---Purpose: Restores the entire MFT font
	--	    from the file $CSF_MDTVFontDirectory/<anAliasName>.dat  
	--	    And returns TRUE if the file have been restores correctly.

	UnderlinePosition (me) returns Length from Quantity;
	---Level: Public 
	---Purpose: Returns the Underline descent position from the origin 
	--	   of the text according to the current font attributes.

	----------------------------
	-- Category: Private methods
	----------------------------

	Open (myclass;
		aFileName: AsciiString from TCollection;
		aFileMode: OpenMode from OSD)
		returns FileHandle from MFT is private;
	---Purpose: Open the file ,load and verify the header
	--	   and returns a file handle >= 0

	Close (myclass; aFileHandle: FileHandle from MFT)
		returns Boolean from Standard is private;
	---Purpose: Close the file.
	--	   Returns TRUE if the file was successfully closed.

	Close (me: mutable)
		returns Boolean from Standard is private;
	---Purpose: Saves updated records and Close this file.
	--	   Returns TRUE if the file was successfully closed.

	Read (myclass; aRecord: in out FileRecord from MFT)
		returns Boolean from Standard is private;
	---Purpose: Reads a record from the file.
	--	   Returns TRUE if the file was successfully read.

	Write (myclass; aRecord: in out FileRecord from MFT)
		returns Boolean from Standard is private;
	---Purpose: Writes a record to the file.
	--	   Returns TRUE if the file was successfully written.

	Locate (myclass; aRecord: in out FileRecord from MFT;
		aFilePosition: FilePosition from MFT)
		returns Address from Standard is private;
	---Purpose: Locates an information from the file record.
	--	   and returns the info address.
	--  Warning: May read or write the current record
	--	   from/to the file and reload an other record
	--	   according the file position info.

	Path (myclass;
		aFileName: AsciiString from TCollection;
		anExtension: CString from Standard = ".mft")
		returns CString from Standard is private;
	---Purpose: Computes the full path of the font file name
	--	    $CSF_MDTVFontDirectory/<aFileName><anExtension>  

	MaxCharPosition (me)
		returns Integer from Standard is private;
	---Purpose: Returns the max position of any defined char
	--	   in the header of the file according with the
	--	   type of the font.

	SetTextAttribs (me : mutable;
		aString: CString from Standard;
		anOrientation: PlaneAngle from Quantity = 0.0) is private;
	---Purpose: Sets the text attributes.
	--  <aString> : the string to interpret 
	--  <anOrientation> : the orientation angle in RAD from horizontal. 

	SetTextAttribs (me : mutable;
		aString: ExtString from Standard;
		anOrientation: PlaneAngle from Quantity = 0.0)
	---Purpose: Sets the extended text attributes.
	--  <aString> : the string to interpret 
	--  <anOrientation> : the orientation angle in RAD from horizontal. 
	raises FontManagerError from MFT is private;
	---Purpose:  Trigger - If the font is not a composite font and
	--	   the string is not ASCII.

	IsDefinedChar (me;
		aPosition: Integer from Standard)
		returns Boolean from Standard
	---Purpose: Returns TRUE if the char at position <aPosition> is defined
	--	    in the header of the file.
	raises FontManagerError from MFT is private;
	---Purpose:  Trigger - If the position <aPosition> is < 0 or > MaxCharPosition(). 

	FirstDefinedChar (me)
		returns Integer from Standard is private;
	---Purpose: Returns the first defined char position 
	--	    in the header of the file..

	LastDefinedChar (me)
		returns Integer from Standard is private;
	---Purpose: Returns the last defined char position 
	--	    in the header of the file..

	SetChar (me: mutable;
		aPosition: Integer from Standard) is private;
	---Purpose: Enable the char at position <aPosition> for reading.

	DrawChar (me: mutable;
		aTextManager: TextManager from MFT;
		aPosition: Integer from Standard) 
		returns Boolean from Standard is private;
	---Purpose: Drawn the char at position <aPosition> 
	--   with the draw manager <aTextManager>.
	--   and returns FALSE if the drawing must be ended.

	ComputeBoundingBox (me: mutable;
		aPosition: Integer from Standard) is private;
	---Purpose: Computes the bounding box of the char position <aPosition>.

	NextCommand (myclass; aRecord: in out FileRecord from MFT)
		returns CommandDescriptor from MFT is private;
	---Purpose: Returns the next command descriptor
	--	    from the current char (see SetChar()).
	--  Warning: the last command of the char descriptor
	--	   has a type MFC_TOC_ENDCHAR.

        Value(myclass;
		aDescriptor: CommandDescriptor from MFT;
                aRank: Integer from Standard)
                returns TypeOfValue from MFT
        ---Purpose: Returns the value type at position <aRank>
        --          from the descriptor command.
        raises FontManagerError from MFT is private;
        ---Purpose:  Trigger - If the position <aRank> is < 1 or > the command length.

	IValue (myclass; aRecord: in out FileRecord from MFT;
		aRank: Integer)
		returns Integer from Standard
	---Purpose: Returns the integer parameter at position <aRank>
	--	    of the current command.
	raises TypeMismatch from Standard is private;
	---Purpose:  Trigger --If the position <aRank> is < 1 or > the command length. 
	--	    or if the value is not an INT value.

	FValue (myclass; aRecord: in out FileRecord from MFT;
		aRank: Integer)
		returns ShortReal from Standard
	---Purpose: Returns the float parameter at position <aRank>
	--	    of the current command.
	raises TypeMismatch from Standard is private;
	---Purpose:  Trigger  - If the position <aRank> is < 1 or > the command length. 
	--	    or if the value is not a FLOAT value.

	SValue (myclass; aRecord: in out FileRecord from MFT;
		aRank: Integer)
		returns CString from Standard
	---Purpose: Returns the string parameter at position <aRank>
	--	    of the current command.
	raises TypeMismatch from Standard is private;
	---Purpose:  Trigger - If the position <aRank> is < 1 or > the command length. 
	--	    or if the value is not a STRING value.

	Dump (me : mutable; aPosition: Integer from Standard) is private;
	---Purpose: Dumps the font descriptor of the character at
	--    	    position <aPosition>.

fields

	myFileName:		AsciiString from TCollection;
	myFileMode:		OpenMode from OSD;
	myFileHandle:		FileHandle from MFT;
	myIsComposite:		Boolean from Standard;
	myIsFixedPitch:		Boolean from Standard;
	myItalicAngle:		ShortReal from Standard;
	myPaintType:		Integer from Standard;
	myCharWidth:		ShortReal from Standard;
	myCharHeight:		ShortReal from Standard;
	myCharSlant:		ShortReal from Standard;
	myCharPrecision:	ShortReal from Standard;
	myCharCapsHeight:	Boolean from Standard;
	myFileHeader:		FileRecord from MFT;
	myCharEntries:		FileRecord from MFT;
	myCommandBuffer:	FileRecord from MFT;

end FontManager from MFT;
