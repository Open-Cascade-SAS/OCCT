-- Created on: 2002-10-29
-- Created by: Michael SAZONOV
-- Copyright (c) 2002-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


package BinMDF

        ---Purpose: This package provides classes and methods to
        --          translate a transient DF into a persistent one and
        --          vice versa.
        --          
        --          Driver
        --          
        --          A driver is a tool used to translate a transient
        --          attribute into a persistent one and vice versa.
        --          
        --          Driver Table
        --          
        --          A driver table is an object building links between
        --          object types and object drivers. In the
        --          translation process, a driver table is asked to
        --          give a translation driver for each current object
        --          to be translated.

uses
    TCollection,
    TColStd,
    TDF,
    CDM,
    BinObjMgt

is

    deferred class ADriver; -- Attribute Storage/Retrieve Driver.

    class ReferenceDriver;  -- Driver for reference

    class TagSourceDriver;  -- Driver for TDF_TagSource

    private alias StringIdMap is DataMapOfAsciiStringInteger from TColStd;

    -- Map (Type, ADriver)
    class TypeADriverMap instantiates DataMap from TCollection
        (Type from Standard,
         ADriver from BinMDF,
         MapTransientHasher from TColStd);

    -- Double Map (Type, Integer ID)
    class TypeIdMap instantiates DoubleMap from TCollection
        (Type from Standard,
         Integer from Standard,
         MapTransientHasher from TColStd,
         MapIntegerHasher from TColStd);

    -- Attribute Storage Driver Table.
    class ADriverTable;

    AddDrivers (aDriverTable : ADriverTable  from BinMDF;
                aMsgDrv      : MessageDriver from CDM);
        ---Purpose: Adds the attribute storage drivers to <aDriverTable>.

end BinMDF;
