-- Created on: 1993-02-02
-- Created by: Christian CAILLET
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



deferred class GeneralModule  from Interface  inherits TShared

    ---Purpose : This class defines general services, which must be provided
    --           for each type of Entity (i.e. of Transient Object processed
    --           by an Interface) : Shared List, Check, Copy, Delete, Category
    --           
    --           To optimise processing (e.g. firstly bind an Entity to a Module
    --           then calls  Module), each recognized Entity Type corresponds
    --           to a Case Number, determined by the Protocol each class of
    --           GeneralModule belongs to.

uses Transient, HAsciiString from TCollection,
     InterfaceModel, ShareTool, Check, EntityIterator, CopyTool

is

    FillShared (me; model : InterfaceModel; CN : Integer; ent : Transient;
    	iter : in out EntityIterator)  is virtual;
    ---Purpose : Specific filling of the list of Entities shared by an Entity
    --           <ent>, according a Case Number <CN> (formerly computed by
    --           CaseNum), considered in the context of a Model <model>
    --           Default calls FillSharedCase (i.e., ignores the model)
    --           Can be redefined to use the model for working

    FillSharedCase (me; CN : Integer; ent : Transient;
    	iter : in out EntityIterator)  is deferred;
    ---Purpose : Specific filling of the list of Entities shared by an Entity
    --           <ent>, according a Case Number <CN> (formerly computed by
    --           CaseNum). Can use the internal utility method Share, below

    Share (me; iter : in out EntityIterator; shared : Transient);
    ---Purpose : Adds an Entity to a Shared List (uses GetOneItem on <iter>)

    ListImplied (me; model : InterfaceModel; CN : Integer; ent : Transient;
    	iter : in out EntityIterator)  is virtual;
    ---Purpose : List the Implied References of <ent> considered in the context
    --           of a Model <model> : i.e. the Entities which are Referenced
    --           while not considered as Shared (not copied if <ent> is,
    --           references not renewed by CopyCase but by ImpliedCase, only
    --           if referenced Entities have been Copied too)
    --           FillShared + ListImplied give the complete list of References
    --           Default calls ListImpliedCase (i.e. ignores the model)
    --           Can be redefined to use the model for working

    ListImpliedCase (me; CN : Integer; ent : Transient;
    	iter : in out EntityIterator)  is virtual;
    ---Purpose : List the Implied References of <ent> (see above)
    --           are Referenced while not considered as Shared (not copied if
    --           <ent> is, references not renewed by CopyCase but by
    --           ImpliedCase, only if referenced Entities have been Copied too)
    --           FillSharedCase + ListImpliedCase give the complete list of
    --           Referenced Entities
    --           The provided default method does nothing (Implied References
    --           are specific of a little amount of Entity Classes).


    CheckCase (me; CN : Integer; ent : Transient; shares : ShareTool;
    	       ach    : in out Check)  is deferred;
    ---Purpose : Specific Checking of an Entity <ent>
    --           Can check context queried through a ShareTool, as required


    CanCopy (me; CN : Integer; ent : Transient) returns Boolean  is virtual;
    ---Purpose : Specific answer to the question "is Copy properly implemented"
    --           Remark that it should be in phase with the implementation of
    --           NewVoid+CopyCase/NewCopyCase
    --           Default returns always False, can be redefined

    Dispatch (me; CN : Integer;
    	      entfrom : Transient; entto : out mutable Transient;
    	      TC : in out CopyTool)  returns Boolean  is virtual;
    ---Purpose : Dispatches an entity
    --           Returns True if it works by copy, False if it just duplicates
    --           the starting Handle
    --           
    --           Dispatching means producing a new entity, image of the
    --           starting one, in order to be put into a new Model, this Model
    --           being itself the result of a dispatch from an original Model
    --           
    --           According to the cases, dispatch can either
    --           * just return <entto> as equating <entfrom>
    --             -> the new model designates the starting entity : it is
    --             lighter, but the dispatched entity being shared might not be
    --             modified for dispatch
    --           * copy <entfrom> to <entto>
    --             by calling NewVoid+CopyCase (two steps) or NewCopiedCase (1)
    --             -> the dispatched entity is a COPY, hence it can be modified
    --             
    --           The provided default just duplicates the handle without
    --           copying, then returns False. Can be redefined


    NewVoid (me; CN : Integer; entto : out mutable Transient)
    	returns Boolean  is deferred;
    ---Purpose : Creates a new void entity <entto> according to a Case Number
    --           This entity remains to be filled, by reading from a file or
    --           by copying from another entity of same type (see CopyCase)

    CopyCase (me; CN : Integer;
    	      entfrom : Transient; entto : mutable Transient;
    	      TC : in out CopyTool)  is deferred;
    ---Purpose : Specific Copy ("Deep") from <entfrom> to <entto> (same type)
    --           by using a CopyTool which provides its working Map.
    --           Use method Transferred from CopyTool to work

    NewCopiedCase (me; CN : Integer;
    	    	   entfrom : Transient; entto : out mutable Transient;
    	    	   TC : in out CopyTool)  returns Boolean  is virtual;
    ---Purpose : Specific operator (create+copy) defaulted to do nothing.
    --           It can be redefined : When it is not possible to work in two
    --           steps (NewVoid then CopyCase). This can occur when there is
    --           no default constructor : hence the result <entto> must be
    --           created with an effective definition.
    --           Remark : if NewCopiedCase is defined, CopyCase has nothing to do
    --           Returns True if it has produced something, false else

    RenewImpliedCase (me; CN : Integer;
    	         entfrom : Transient; entto : mutable Transient;
    	         TC : CopyTool)  is virtual;
    ---Purpose : Specific Copying of Implied References
    --           A Default is provided which does nothing (must current case !)
    --           Already copied references (by CopyFrom) must remain unchanged
    --           Use method Search from CopyTool to work

    WhenDeleteCase (me; CN : Integer;
    	    	ent : mutable Transient; dispatched : Boolean)  is virtual;
    ---Purpose : Prepares an entity to be deleted. What does it mean :
    --           Basically, any class of entity may define its own destructor
    --           By default, it does nothing but calling destructors on fields
    --           With the Memory Manager, it is useless to call destructor,
    --           it is done automatically when the Handle is nullified(cleared)
    --           BUT this is ineffective in looping structures (whatever these
    --           are "Implied" references or not).
    --           
    --           THUS : if no loop may appear in definitions, a class which
    --           inherits from TShared is correctly managed by automatic way
    --           BUT if there can be loops (or simply back pointers), they must
    --           be broken, for instance by clearing fields of one of the nodes
    --           The default does nothing, to be redefined if a loop can occur
    --           (Implied generally requires WhenDelete, but other cases can
    --           occur)
    --           
    --  Warning : <dispatched> tells if the entity to be deleted has been
    --           produced by Dispatch or not. Hence WhenDelete must be in
    --           coherence with Dispatch
    --           Dispatch can either copy or not.
    --           If it copies the entity, this one should be deleted
    --           If it doesnt (i.e. duplicates the handle) nothing to do
    --           
    --           If <dispatch> is False, normal deletion is to be performed

    CategoryNumber (me; CN : Integer; ent : Transient; shares : ShareTool)
    	returns Integer  is virtual;
    ---Purpose : Returns a category number which characterizes an entity
    --           Category Numbers are managed by the class Category
    --           <shares> can be used to evaluate this number in the context
    --           Default returns 0 which means "unspecified"

    Name  (me; CN : Integer; ent : Transient; shares : ShareTool)
    	returns HAsciiString from TCollection  is virtual;
    ---Purpose : Determines if an entity brings a Name (or widerly, if a Name
    --           can be attached to it, through the ShareTool
    --           By default, returns a Null Handle (no name can be produced)
    --           Can be redefined
    --           
    --  Warning : While this string may be edited on the spot, if it is a read
    --           field, the returned value must be copied before.

end GeneralModule;
