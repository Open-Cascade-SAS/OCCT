-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class AutoDesignGroupAssignment from StepAP214 

inherits GroupAssignment from StepBasic

uses

	HArray1OfAutoDesignGroupedItem from StepAP214, 
	AutoDesignGroupedItem from StepAP214, 
	Group from StepBasic
is

	Create returns AutoDesignGroupAssignment;
	---Purpose: Returns a AutoDesignGroupAssignment


	Init (me : mutable;
	      aAssignedGroup : Group from StepBasic;
	      aItems : HArray1OfAutoDesignGroupedItem from StepAP214) is virtual;

	-- Specific Methods for Field Data Access --

	SetItems(me : mutable; aItems : HArray1OfAutoDesignGroupedItem);
	Items (me) returns HArray1OfAutoDesignGroupedItem;
	ItemsValue (me; num : Integer) returns AutoDesignGroupedItem;
	NbItems (me) returns Integer;

fields

	items : HArray1OfAutoDesignGroupedItem from StepAP214; -- a SelectType

end AutoDesignGroupAssignment;
