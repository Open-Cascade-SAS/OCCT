-- Created on: 1993-08-04
-- Created by: Martine LANGLOIS
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MakeVectorWithMagnitude2d from StepToGeom

    ---Purpose: This class implements the mapping between classes 
    --          Vector from StepGeom which describes a VectorWithMagnitude 
    --          from Prostep and VectorWithMagnitude from Geom2d.
  
uses 
     VectorWithMagnitude from Geom2d,
     Vector from StepGeom

is 

    Convert ( myclass; SV : Vector from StepGeom;
                       CV : out VectorWithMagnitude from Geom2d )
    returns Boolean from Standard;

end MakeVectorWithMagnitude2d;
