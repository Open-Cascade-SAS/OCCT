-- File:	ShapeAnalysis_WireOrder.cdl
-- Created:	Wed Jun  3 12:06:27 1998
-- Author:	data exchange team
--		<det@nnov.matra-dtv.fr>
---Copyright:	 Matra Datavision 1998


class WireOrder from ShapeAnalysis 

	---Purpose: This class is intended to control and, if possible, redefine
    	--          the order of a list of edges which define a wire
    	--          Edges are not given directly, but as their bounds (start,end)
    	--           
    	--          This allows to use this tool, either on existing wire, or on
    	--          data just taken from a file (coordinates are easy to get)
    	--           
    	--          It can work, either in 2D, or in 3D, but not miscible
    	--          Warning about tolerance : according to the mode (2D/3D), it
        --          must be given as 2D or 3D (i.e. metric) tolerance, uniform
        --          on the whole list
        --           
        --          Two phases : firstly add the couples (start,end)
        --          secondly perform then get the result

uses
    XY from gp,
    XYZ from gp,
    HSequenceOfXYZ from TColgp,
    HArray1OfInteger from TColStd

raises
    TypeMismatch from Standard

is

    Create returns WireOrder from ShapeAnalysis;
    	---Purpose: Empty constructor

    Create(mode3d: Boolean; tol: Real) returns WireOrder from ShapeAnalysis;
    	---Purpose : Creates a WireOrder in 3D (if mode3d is True) or 2D (if False)
    	--           with a tolerance

    SetMode(me : in out; mode3d: Boolean; tol    : Real);
    	---Purpose : Sets new values. Clears the connexion list
    	--           If <mode3d> changes, also clears the edge list (else, doesnt)

    Tolerance(me) returns Real;
    	---Purpose : Returns the working tolerance

    Clear(me: in out);
    	---Purpose : Clears the list of edges, but not mode and tol

    Add(me: in out; start3d, end3d: XYZ from gp)
    	---Purpose : Adds a couple of points 3D (start,end)
    raises TypeMismatch;
    	--           Error if initial mode was 2D

    Add(me: in out; start2d, end2d: XY from gp)
    	---Purpose : Adds a couple of points 2D (start,end)
    raises TypeMismatch;
    	--           Error if initial mode was 3D

    NbEdges(me) returns Integer;
    	---Purpose : Returns the count of added couples of points (one per edges)
	
    KeepLoopsMode(me: in out) returns Boolean;
        ---C++: return&
	---Purpose : If this mode is True method perform does not sort edges of
	--           different loops. The resulting order is first loop, second
	--           one etc...
	
    Perform(me: in out; closed: Boolean = Standard_True);
    	---Purpose : Computes the better order
    	--           If <closed> is True (D) considers also closure
    	--           Optimised if the couples were already in order
    	--           The criterium is : two couples in order if distance between
    	--           end-prec and start-cur is less then starting tolerance <tol>
    	--           Else, the smallest distance is reached
    	--           Gap corresponds to a smallest distance greater than <tol>

    IsDone(me) returns Boolean;
    	---Purpose : Tells if Perform has been done
   	--           Else, the following methods returns original values

    Status(me) returns Integer;
    	---Purpose : Returns the status of the order (0 if not done) :
    	--            0 : all edges are direct and in sequence
    	--            1 : all edges are direct but some are not in sequence
    	--            2 : in addition, unresolved gaps remain
    	--           -1 : some edges are reversed, but no gap remain
    	--           -2 : some edges are reversed and some gaps remain
    	--           -10 : COULD NOT BE RESOLVED, Failure on Reorder
    	--           gap : regarding starting <tol>

    Ordered(me; n: Integer) returns Integer;
    	---Purpose : Returns the number of original edge which correspond to the
    	--           newly ordered number <n>
    	--  Warning : the returned value is NEGATIVE if edge should be reversed

    XYZ(me; num: Integer; start3d, end3d : out XYZ from gp);
    	---Purpose : Returns the values of the couple <num>, as 3D values

    XY(me; num: Integer; start2d, end2d: out XY from gp);
    	---Purpose : Returns the values of the couple <num>, as 2D values

    Gap(me; num : Integer = 0) returns Real;
    	---Purpose : Returns the gap between a couple and its preceeding
    	--           <num> is considered ordered
    	--           If <num> = 0 (D), returns the greatest gap found

    SetChains(me : in out; gap : Real);
    	---Purpose : Determines the chains inside which successive edges have a gap
    	--           less than a given value. Queried by NbChains and Chain

    NbChains(me) returns Integer;
    	---Purpose : Returns the count of computed chains

    Chain(me; num: Integer; n1,n2: out Integer);
    	---Purpose : Returns, for the chain n0 num, starting and ending numbers of
    	--           edges. In the list of ordered edges (see Ordered for originals)

    SetCouples(me: in out; gap: Real);
    	---Purpose : Determines the couples of edges for which end and start fit
    	--           inside a given gap. Queried by NbCouples and Couple

    NbCouples(me) returns Integer;
    	---Purpose : Returns the count of computed couples

    Couple(me; num: Integer; n1, n2: out Integer);
    	---Purpose : Returns, for the couple n0 num, the two implied edges
    	--           In the list of ordered edges

fields

    myKeepLoops : Boolean from Standard;
    myOrd     : HArray1OfInteger from TColStd;
    myChains  : HArray1OfInteger from TColStd;
    myCouples : HArray1OfInteger from TColStd;
    myXYZ     : HSequenceOfXYZ   from TColgp;
    myTol     : Real;
    myGap     : Real;
    myStat    : Integer;
    myMode    : Boolean;

end WireOrder;
