-- Created on: 2002-10-29
-- Created by: Michael SAZONOV
-- Copyright (c) 2002-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



package BinObjMgt 

---Purpose: This package defines services to manage the storage
--          grain of data produced by applications.

uses
    TDF,
    Standard,
    TCollection,
    TColStd

is

        -- Storage Relocation Table
    alias SRelocationTable is IndexedMapOfTransient from TColStd;

        -- Retrieval Relocation Table
    alias RRelocationTable is DataMapOfIntegerTransient from TColStd;

    primitive PChar;            -- pointer to Character from Standard;
    primitive PByte;            -- pointer to Byte from Standard;
    primitive PExtChar;         -- pointer to ExtCharacter from Standard;
    primitive PInteger;         -- pointer to Integer from Standard;
    primitive PReal;            -- pointer to Real from Standard;
    primitive PShortReal;       -- pointer to ShortReal from Standard;

    class Persistent;

end BinObjMgt;
