-- Created on: 1991-01-14
-- Created by: Arnaud BOUZY
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class UnaryFunction from Expr

inherits UnaryExpression from Expr  

    ---Purpose: Defines the use of an unary function in an expression 
    --          with a given argument.

uses NamedUnknown from Expr,
    AsciiString from TCollection,
    Array1OfNamedUnknown from Expr,
    Array1OfReal from TColStd,
    GeneralFunction from Expr,
    GeneralExpression from Expr

raises InvalidFunction from Expr, 
    NumericError from Standard,
    NotEvaluable from Expr

is

    Create(func : GeneralFunction; exp : GeneralExpression)
    ---Purpose: Creates me as <func>(<exp>).
    --          Raises exception if <func> is not unary.
    returns mutable UnaryFunction
    raises InvalidFunction;

    Function(me)
    ---Purpose: Returns the function defining <me>.
    returns GeneralFunction;
    
    ShallowSimplified(me) 
    ---Purpose: Returns a GeneralExpression after a simplification 
    --          of the arguments of <me>.
    returns any GeneralExpression
    raises NumericError;

    Copy(me)
    ---Purpose: Returns a copy of <me> having the same unknowns and functions.
    returns mutable like me;
    
    IsIdentical(me; Other : GeneralExpression)
    ---Purpose: Tests if <me> and <Other> define the same expression.
    --          This method does not include any simplification before
    --          testing.
    returns Boolean;

    IsLinear(me)
    returns Boolean;

    Derivative(me; X : NamedUnknown)
    ---Purpose: returns the derivative on <X> unknown of <me>. 
    returns any GeneralExpression;

    Evaluate(me; vars : Array1OfNamedUnknown; vals : Array1OfReal)
    ---Purpose: Returns the value of <me> (as a Real) by 
    --          replacement of <vars> by <vals>.
    --          Raises NotEvaluable if <me> contains NamedUnknown not 
    --          in <vars> or NumericError if result cannot be computed.
    returns Real
    raises NotEvaluable,NumericError;

    String(me)
    ---Purpose: returns a string representing <me> in a readable way.
    returns AsciiString;

fields

    myFunction : GeneralFunction;

end UnaryFunction;
