-- Created on: 1993-09-22
-- Created by: Didier PIFFAULT
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Edge from BRepMesh 

  ---Purpose: 


uses    Boolean from Standard,
        Integer from Standard,
        DegreeOfFreedom from BRepMesh


is            Create
              returns Edge from BRepMesh;
    	          ---C++: inline
    	          
              Create       (vDebut    : Integer from Standard;
                            vFin      : Integer from Standard;
                            canMove   : DegreeOfFreedom from BRepMesh)
              ---Purpose: Contructs a link beetween to vertices.
              returns Edge from BRepMesh;


            FirstNode      (me)
              ---Purpose: Give the index of first node of the Link.
              ---C++: inline
              returns Integer from Standard
              is static;


            LastNode       (me)
              ---Purpose: Give the index of Last node of the Link.
              ---C++: inline
              returns Integer from Standard
              is static;


            Movability     (me)
              ---C++: inline
              returns DegreeOfFreedom from BRepMesh
              is static;


            SetMovability  (me   : in out;
                            Move : DegreeOfFreedom from BRepMesh)
              is static;

       HashCode       (me;
                       Upper : Integer from Standard)
          returns Integer from Standard
          ---C++: function call
          is static;


        SameOrientation(me; Other : Edge from BRepMesh)
          returns Boolean from Standard
          is static;


        IsEqual        (me; Other : Edge from BRepMesh)
          returns Boolean from Standard
          ---C++: alias operator ==
          is static;


        fields  myFirstNode  : Integer from Standard;
                myLastNode   : Integer from Standard;
                myMovability : DegreeOfFreedom from BRepMesh;

        end Edge;
