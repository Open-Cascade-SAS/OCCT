-- Created on: 2001-08-28
-- Created by: data exchange team
-- Copyright (c) 2001-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Curve from ShapeCustom 

	---Purpose: Converts BSpline curve to periodic

uses

    Curve from Geom

is

    Create returns Curve from ShapeCustom;
    
    Create (C: Curve from Geom) returns Curve from ShapeCustom;
    
    Init (me: in out; C: Curve from Geom);
    
    ConvertToPeriodic (me: in out; substitute: Boolean; preci: Real = -1)
    returns Curve from Geom;
        ---Purpose: Tries to convert the Curve to the Periodic form
    	--          Returns the resulting curve
    	--          Works only if the Curve is BSpline and is closed with 
        --          Precision::Confusion()
    	--          Else, or in case of failure, returns a Null Handle
fields

    myCurve: Curve from Geom;

end Curve;
