-- Created on: 2008-01-21
-- Created by: Galina KULIKOVA
-- Copyright (c) 2008-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ParamList from Interface inherits TShared from MMgt

	---Purpose: 

uses
    FileParameter from Interface,VectorOfFileParameter from Interface

raises  RangeError from Standard,
    	OutOfRange from Standard,
	OutOfMemory from Standard 
is

    Create( theIncrement : Integer = 256) returns ParamList from Interface;
    ---Purpose: Creates an vector with size of memmory blok equal to theIncrement
    
    
    Length (me) returns Integer from Standard;
    	---Purpose: Returns the number of elements of <me>.
    	--           
        ---C++: inline

    Lower (me) returns Integer from Standard;
    	---Purpose:  Returns the lower bound.
    	-- Warning
    	--Client programs of the Array1 class must be independent of the first item range.--          
    	---C++: inline
	
    Upper (me) returns Integer from Standard;
    	---Purpose: Returns the upper bound.
    	-- Warning
    	--Client programs of the Array1 class must be independent of the first item range.--          
    	---C++: inline

    SetValue (me : mutable; Index: Integer from Standard; Value: FileParameter from Interface) 
    	---Purpose: Assigns the value <Value> to the <Index>-th item of this array.
    raises OutOfRange from Standard;

    Value (me; Index:Integer from Standard) returns FileParameter from Interface
    	---Purpose: Return the value of  the  <Index>th element of the
    	--          array.
    	---C++: alias operator ()
    	---C++: return const &
    raises OutOfRange from Standard;
    
    ChangeValue (me: mutable; Index:Integer from Standard) returns FileParameter from Interface
    	---Purpose: return the value  of the <Index>th element  of the
    	--          array.
    	--
    	---C++: alias operator ()
    	---C++: return &
    raises OutOfRange from Standard;
    
    Clear(me: mutable);
    

    
    
fields

    	
  myVector : VectorOfFileParameter;

end ParamList;
