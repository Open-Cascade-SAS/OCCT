-- Created on: 1996-01-29
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class WireToFace from TopOpeBRepBuild

---Purpose: 
-- This class builds faces from a set of wires  SW and a face F.
-- The face must have and underlying surface, say S.
-- All of the edges of all of the wires must have a 2d representation 
-- on surface S (except if S is planar)

uses

    Wire from TopoDS,
    Face from TopoDS,
    ListOfShape from TopTools

is

    Create returns WireToFace;
     
    Init(me : in out)
    is static;
    
    AddWire(me : in out; W : Wire from TopoDS)
    is  static;
     	
    MakeFaces(me : in out; 
    	      F : Face from TopoDS;
    	      LF : in out ListOfShape from TopTools)
    is static;

fields 

    myLW : ListOfShape from TopTools;
    
end WireToFace;
