-- Created on: 1996-09-04
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Pipe from LocOpe 

	---Purpose: Defines a  pipe  (near from   Pipe from BRepFill),
	--          with modifications provided for the Pipe feature.

uses Pipe from BRepFill,

     ListOfShape               from TopTools,
     DataMapOfShapeListOfShape from TopTools,
     Curve                     from  Geom,      
     Shape                     from TopoDS,
     Wire                      from TopoDS,     
     SequenceOfPnt             from TColgp,
     SequenceOfCurve           from TColGeom
     

raises NoSuchObject from Standard,
       DomainError  from Standard

is

    Create (Spine   : Wire from TopoDS;
    	    Profile : Shape from TopoDS)
	    
    	returns Pipe from LocOpe;


    Spine(me)
    
    	returns Shape from TopoDS
	---C++: inline
	---C++: return const &
	is static;


    Profile(me)
    
    	returns Shape from TopoDS
	---C++: inline
	---C++: return const &
	is static;


    FirstShape(me)
    
    	returns Shape from TopoDS
	---C++: inline
	---C++: return const &
	is static;


    LastShape(me)
    
    	returns Shape from TopoDS
	---C++: inline
	---C++: return const &
	is static;


    Shape(me)
    
    	returns Shape from TopoDS
	---C++: return const &
	is static;


    Shapes(me: in out; S: Shape from TopoDS)
    
    	returns ListOfShape from TopTools
	---C++: return const &
    	raises NoSuchObject from Standard,
	       -- The exception is raised if S is not a subshape of the profile
               DomainError  from Standard
	       -- The exception is raised if S is neither a vertex nor
	       -- an edge
	is static;


    Curves(me: in out; Spt: SequenceOfPnt from TColgp)

	---C++: return const &
    	returns SequenceOfCurve from TColGeom
	is static;

    BarycCurve(me: in out) 
     
    	returns  Curve  from  Geom 
	is  static;

fields

    myPipe : Pipe                      from BRepFill;
    myMap  : DataMapOfShapeListOfShape from TopTools;
    myRes  : Shape                     from TopoDS;
    myGShap: ListOfShape               from TopTools;
    myCrvs : SequenceOfCurve           from TColGeom;
    myFirstShape : Shape             from TopoDS;
    myLastShape  : Shape             from TopoDS;

end Pipe;
