-- Created on: 1993-08-10
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


package HLRTopoBRep

	---Purpose: This     Package  provides  some       topological
	--          reconstruction services needed  by the Hidden Line
	--          Removal Algorithms   using OutLine  and    IsoLine
	--          facilities, applied  to an object represented by a
	--          BRep data structure.

uses
    Standard,
    MMgt,
    TCollection,
    TColStd,
    TopoDS,
    TopTools,
    TopExp,
    gp,
    Geom2d,
    IntSurf,
    BRepAdaptor,
    BRepTopAdaptor,
    Contap,
    HLRAlgo
    
is
    class VData;

    class ListOfVData            instantiates List    from TCollection 
    	(VData from HLRTopoBRep);

    class MapOfShapeListOfVData  instantiates DataMap from TCollection
    	(Shape          from TopoDS,
         ListOfVData    from HLRTopoBRep,
         ShapeMapHasher from TopTools);

    class FaceData;

    class DataMapOfShapeFaceData instantiates DataMap from TCollection
    	(Shape          from TopoDS,
	 FaceData       from HLRTopoBRep,
	 ShapeMapHasher from TopTools);
					
    class Data;

    class FaceIsoLiner;
    
    class OutLiner;

    class DSFiller;

end HLRTopoBRep;
