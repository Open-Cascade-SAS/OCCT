-- Created on: 1993-06-23
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ShapeData from TopOpeBRepDS

uses 
    
    ListOfInterference from TopOpeBRepDS,
    ListOfShape from TopTools,
    Config from TopOpeBRepDS,
    Orientation from TopAbs
    
is  
    
    Create returns ShapeData;
    Interferences(me) returns ListOfInterference;
    ---C++:return const & 
    ChangeInterferences(me:in out) returns ListOfInterference;
    ---C++:return &
    
    Keep(me) returns Boolean from Standard
    is static;
    ChangeKeep(me : in out; B : Boolean from Standard)
    is static;

fields

    myInterferences : ListOfInterference from TopOpeBRepDS;
    mySameDomain    : ListOfShape from TopTools;
    mySameDomainRef : Integer from Standard;
    mySameDomainOri : Config from TopOpeBRepDS;
    mySameDomainInd : Integer;
    myOrientation : Orientation from TopAbs;
    myOrientationDef : Boolean;
    myAncestorRank : Integer; -- 1 or 2
    myKeep      : Boolean from Standard;

friends 
    
    class DataStructure from TopOpeBRepDS

end ShapeData from TopOpeBRepDS;
