-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PresentationStyleAssignment from StepVisual 

inherits TShared from MMgt

uses

	HArray1OfPresentationStyleSelect from StepVisual, 
	PresentationStyleSelect from StepVisual
is

	Create returns PresentationStyleAssignment;
	---Purpose: Returns a PresentationStyleAssignment

	Init (me : mutable;
	      aStyles : HArray1OfPresentationStyleSelect from StepVisual) is virtual;

	-- Specific Methods for Field Data Access --

	SetStyles(me : mutable; aStyles : HArray1OfPresentationStyleSelect);
	Styles (me) returns HArray1OfPresentationStyleSelect;
	StylesValue (me; num : Integer) returns PresentationStyleSelect;
	NbStyles (me) returns Integer;

fields

	styles : HArray1OfPresentationStyleSelect from StepVisual; -- a SelectType

end PresentationStyleAssignment;
