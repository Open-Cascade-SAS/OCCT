-- Created on: 1993-01-09
-- Created by: CKY / Contract Toubro-Larsen ( Anand NATRAJAN )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ExternalRefFile from IGESBasic  inherits IGESEntity

        ---Purpose: defines ExternalRefFile, Type <416> Form <1>
        --          in package IGESBasic
        --          Used when entire reference file is to be instanced

uses

        HAsciiString from TCollection

is

        Create returns ExternalRefFile;

        -- Specific Methods pertaining to the class

        Init (me : mutable; aFileIdent : HAsciiString);
        ---Purpose : This method is used to set the field of the class
        --           ExternalRefFile
        --       - aFileIdent : External Reference File Identifier

        FileId (me) returns HAsciiString from TCollection;
        ---Purpose : returns External Reference File Identifier

fields

--
-- Class    : IGESBasic_ExternalRefFile
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class ExternalRefFile.
--
-- Reminder : A ExternalRefFile instance is defined by :
--            - an External Reference File Identifier

        theExtRefFileIdentifier : HAsciiString from TCollection;

end ExternalRefFile;
