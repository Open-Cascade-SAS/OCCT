-- Created by: Peter Kurnev
-- Copyright (c) 2010-2014 OPEN CASCADE SAS
-- Copyright (c) 2007-2010 CEA/DEN, EDF R&D, OPEN CASCADE
-- Copyright (c) 2003-2007 OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN, CEDRAT,
--                         EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

--
class CheckerSI from BOPAlgo 
    inherits PaveFiller from BOPAlgo  
    
    ---Purpose: Checks shape on self-interference.

is
    Create 
    	returns CheckerSI from BOPAlgo;  
    ---C++: alias "Standard_EXPORT virtual ~BOPAlgo_CheckerSI();"  
    

    Perform(me:out) 
    	is redefined;   
  

    Init  (me:out) 
    	is redefined protected;

    SetLevelOfCheck(me:out; 
      theLevel: Integer from Standard); 
    ---Purpose:  Sets the level of checking shape on self-interference.
    --           It defines which interferferences will be checked: 
    --           0 - only V/V; 
    --           1 - V/V and V/E; 
    --           2 - V/V, V/E and E/E; 
    --           3 - V/V, V/E, E/E and V/F;
    --           4 - V/V, V/E, E/E, V/F and E/F; 
    --           5 - all interferences, default value. 
 

    PostTreat  (me:out)  
    	is protected;       
    ---Purpose: Provides post-tratment actions 	 
    
    PerformVZ(me:out) 
      is virtual protected; 
       --Purpose: Computes Vertex/Solid interferences 
       
    PerformEZ(me:out) 
      is virtual protected;  
      --Purpose: Computes Edge/Solid interferences 
     
    PerformFZ(me:out) 
      is virtual protected;   
      --Purpose: Computes Face/Solid interferences 
    PerformZZ(me:out) 
      is virtual protected;  
      --Purpose: Computes Solid/Solid interferences 
 
 
fields
    myLevelOfCheck: Integer from Standard is protected;
    
end CheckerSI;
