-- Created on: 1996-09-05
-- Created by: Yves FRICAUD
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MakeLoops from BRepOffset 

	---Purpose: 

uses
    ListOfShape from TopTools,
    AsDes       from BRepAlgo,
    Analyse     from BRepOffset,
    Image       from BRepAlgo,
    DataMapOfShapeShape from TopTools
    
is
    Create;
    
    Build         (me: in out; LF    :        ListOfShape from TopTools;
    	 	    	       AsDes :        AsDes       from BRepAlgo;
		    	       Image : in out Image       from BRepAlgo);	 

    BuildOnContext(me: in out; LContext :        ListOfShape from TopTools;
    	    	    	       Analyse  :        Analyse     from BRepOffset;
    	    	    	       AsDes    :        AsDes       from BRepAlgo;
		    	       Image    : in out Image       from BRepAlgo; 
    	    	    	       InSide   :        Boolean     from Standard);

    BuildFaces    (me: in out; LF    :        ListOfShape from TopTools;
    	    	    	       AsDes :        AsDes       from BRepAlgo;
		    	       Image : in out Image       from BRepAlgo);

fields 
    myVerVerMap  : DataMapOfShapeShape from TopTools; 
		     	
end MakeLoops;
