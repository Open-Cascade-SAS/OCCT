-- Created on: 2002-12-12
-- Created by: data exchange team
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class MaterialPropertyRepresentation from StepRepr
inherits PropertyDefinitionRepresentation from StepRepr

    ---Purpose: Representation of STEP entity MaterialPropertyRepresentation

uses
    RepresentedDefinition from StepRepr,
    Representation from StepRepr,
    DataEnvironment from StepRepr

is
    Create returns MaterialPropertyRepresentation from StepRepr;
	---Purpose: Empty constructor

    Init (me: mutable; aPropertyDefinitionRepresentation_Definition: RepresentedDefinition from StepRepr;
                       aPropertyDefinitionRepresentation_UsedRepresentation: Representation from StepRepr;
                       aDependentEnvironment: DataEnvironment from StepRepr);
	---Purpose: Initialize all fields (own and inherited)

    DependentEnvironment (me) returns DataEnvironment from StepRepr;
	---Purpose: Returns field DependentEnvironment
    SetDependentEnvironment (me: mutable; DependentEnvironment: DataEnvironment from StepRepr);
	---Purpose: Set field DependentEnvironment

fields
    theDependentEnvironment: DataEnvironment from StepRepr;

end MaterialPropertyRepresentation;
