-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class FaceBound from StepShape 

inherits TopologicalRepresentationItem from StepShape 

uses

	Loop from StepShape, 
	Boolean from Standard, 
	HAsciiString from TCollection
is

	Create returns mutable FaceBound;
	---Purpose: Returns a FaceBound


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aBound : mutable Loop from StepShape;
	      aOrientation : Boolean from Standard) is virtual;

	-- Specific Methods for Field Data Access --

	SetBound(me : mutable; aBound : mutable Loop);
	Bound (me) returns mutable Loop;
	SetOrientation(me : mutable; aOrientation : Boolean);
	Orientation (me) returns Boolean;

fields

	bound : Loop from StepShape;
	orientation : Boolean from Standard;

end FaceBound;
