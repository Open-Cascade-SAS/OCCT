-- Created on: 1993-10-21
-- Created by: Jean-Louis FRENKEL
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Modified by  rob 09-oct-96



class Presentation3d from PrsMgr inherits Presentation from PrsMgr

uses
    PresentationManager from PrsMgr,
    Presentation from Prs3d,
    NameOfColor from Quantity,
    Transformation from Geom,
    Length from Quantity,
    ShadingAspect from Prs3d,
    TypeOfPresentation3d from PrsMgr,
    DataStructureManager from Graphic3d,
    Structure from Graphic3d,
    PresentableObjectPointer from PrsMgr,PresentableObject from PrsMgr,
    Prs from PrsMgr,
    Projector from Prs3d,
    KindOfPrs from PrsMgr
is
    Create(aPresentationManager: PresentationManager from PrsMgr;
           aPresentableObject: PresentableObject from PrsMgr)
    returns mutable Presentation3d  from  PrsMgr
    is private;

    KindOfPresentation(me) returns KindOfPrs from PrsMgr is redefined static;

    Destroy(me: mutable) is redefined;
    ---Level: Public
    ---Purpose: Destructor
    ---C++:     alias ~

    Display(me: mutable) 
    is redefined static private;
    
    Display (me: mutable;
             theIsHighlight: Boolean from Standard)
    is static private;
    ---Level: Private;
    ---Purpose: displays myStructure and sets myDisplayReason to theIsHighlight value if
    -- myStructure was not displayed or was invisible
    
    Erase(me: mutable) is redefined static private;

    SetVisible (me: mutable; theValue: Boolean from Standard) is redefined static private;

    Highlight(me: mutable) is redefined static private;
    
    Unhighlight (me) is redefined static private;
    
    IsDisplayed (me) returns Boolean from Standard
    is redefined static private;

    IsHighlighted (me) returns Boolean from Standard
    is redefined static private;


    DisplayPriority(me) returns Integer from Standard
    is redefined static private;
    
    SetDisplayPriority(me:mutable;aNewPrior:Integer from Standard)
    is redefined static private;

    SetZLayer ( me : mutable;
                theLayerId : Integer from Standard )
      is redefined static private;
    ---Purpose: Set Z layer ID for the presentation

    GetZLayer ( me )
      returns Integer from Standard is redefined static private;
    ---Purpose: Get Z layer ID for the presentation

    Clear(me:mutable)
    ---Purpose: removes the whole content of the presentation.
    --          Does not remove the other connected presentations.
    --          
    is redefined static private;


    Color(me:mutable; aColor: NameOfColor from Quantity)
    is static private;
    
    BoundBox(me)
    is static private;
    
---Category: references to other presentation.

    Connect(me; anOtherPresentation: Presentation3d from PrsMgr)
    is static private;
    
---Category: Transformation methods.

    Transform (me; aTransformation: Transformation from Geom)
    is static private;

    Place (me; X,Y,Z: Length from Quantity)
    is static private;

    Multiply (me; aTransformation: Transformation from Geom)
    is static private;

    Move (me; X,Y,Z: Length from Quantity)
    is static private;
    	
 ---Category: Global Aspect methods

    SetShadingAspect(me;
    	             aShadingAspect: ShadingAspect from Prs3d)
    is static private;

    Presentation (me) returns mutable Presentation from Prs3d
    is static;


	    ---Category:  Computed Structures

    Compute(me : mutable; theStructure: Structure from Graphic3d)
    is static private;

    Compute(me : mutable; aProjector: DataStructureManager from Graphic3d)
    returns Structure from Graphic3d
    is static private;

    Compute(me           : mutable; 
    	    aProjector   : DataStructureManager from Graphic3d;
	    TheTrsf      : Transformation from Geom)
    returns Structure from Graphic3d
    is static private;

    Compute(me           :  mutable; 
    	    aProjector   :  DataStructureManager from Graphic3d;
    	    aGivenStruct :  Structure from Graphic3d)
    is static private;

    Compute(me           : mutable; 
    	    aProjector   : DataStructureManager from Graphic3d;
	    TheTrsf      : Transformation from Geom;
    	    aGivenStruct : Structure from Graphic3d)
    is static private;



    Projector(myclass; aProjector: DataStructureManager from Graphic3d)
    returns Projector from Prs3d
    is private;
    
fields

    myStructure: Prs from PrsMgr;
    myDisplayReason: Boolean from Standard;
    myPresentableObject: PresentableObjectPointer from PrsMgr;
friends 
    class PresentationManager from PrsMgr,
    class PresentableObject from PrsMgr,
    class Prs from PrsMgr
end Presentation3d from PrsMgr;
