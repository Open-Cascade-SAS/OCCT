-- Created on: 1993-12-02
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package Blend

uses IntSurf, 
    TColgp, 
    TColStd, 
    Adaptor2d, 
    gp, 
    TopAbs, 
    math, 
    TCollection, 
    MMgt, 
    StdFail,  
    GeomAbs

is

--    deferred generic class SurfaceTool;
    
    generic class Iterator;          -- template class

    deferred class AppFunction;      -- inherits FunctionSetWithDerivatives from math

    deferred class Function;         -- inherits AppFunction from Blend

    deferred class FuncInv;          -- inherits FunctionSetWithDerivatives from math

    deferred class CSFunction;       -- inherits AppFunction from Blend

    deferred class SurfRstFunction;  -- inherits AppFunction from Blend

    deferred class SurfPointFuncInv; -- inherits FunctionSetWithDerivatives from math

    deferred class SurfCurvFuncInv;  -- inherits FunctionSetWithDerivatives from math

    deferred class RstRstFunction;  -- inherits AppFunction from Blend

    deferred class CurvPointFuncInv; -- inherits FunctionSetWithDerivatives from math



    class Point;
    
    generic class Extremity;
    
    generic class PointOnRst;
    
    generic class Line;

    generic class Walking;

    generic class CSWalking;


    class SequenceOfPoint instantiates Sequence from TCollection
    	(Point from Blend);
	
    enumeration Status is 
    	StepTooLarge,
	StepTooSmall,
	Backward,
	SamePoints,
	OnRst1,
	OnRst2,
	OnRst12,
	OK
    end Status;


    enumeration DecrochStatus is 
    	NoDecroch,
	DecrochRst1,
	DecrochRst2,
	DecrochBoth
    end Status;



end Blend;
