-- File:	IGESGeom_ToolCopiousData.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolCopiousData  from IGESGeom

    ---Purpose : Tool to work on a CopiousData. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses CopiousData from IGESGeom,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolCopiousData;
    ---Purpose : Returns a ToolCopiousData, ready to work


    ReadOwnParams (me; ent : mutable CopiousData;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : CopiousData;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : CopiousData;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a CopiousData <ent>, from
    --           its specific (own) parameters

    DirChecker (me; ent : CopiousData) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : CopiousData;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : CopiousData; entto : mutable CopiousData;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : CopiousData;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolCopiousData;
