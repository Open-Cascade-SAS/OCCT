-- File:	IGESData_DefaultGeneral.cdl
-- Created:	Wed Sep  8 16:41:51 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class DefaultGeneral  from IGESData  inherits  GeneralModule  from IGESData

    ---Purpose : Processes the specific case of UndefinedEntity from IGESData
    --           (Case Number 1)

uses OStream, Transient,
     InterfaceModel, Check, ShareTool, EntityIterator, CopyTool,
     IGESEntity, DirChecker

is

    Create returns mutable DefaultGeneral;
    ---Purpose : Creates a DefaultGeneral and puts it into GeneralLib,
    --           bound with a Protocol from IGESData

    OwnSharedCase  (me; CN : Integer; ent : IGESEntity;
    	    	    iter : in out EntityIterator);
    ---Purpose : Lists the Entities shared by an IGESEntity, which must be
    --           an UndefinedEntity


    DirChecker (me; CN : Integer; ent : IGESEntity) returns DirChecker;
    ---Purpose : Returns a DirChecker, specific for each type of Entity
    --           Here, Returns an empty DirChecker (no constraint to check)

    OwnCheckCase (me; CN : Integer; ent : IGESEntity; shares : ShareTool;
    	          ach    : in out Check);
    ---Purpose : Performs Specific Semantic Check for each type of Entity
    --           Here, does nothing (no constraint to check)


    NewVoid (me; CN : Integer; entto : out mutable Transient)
    	returns Boolean;
    ---Purpose : Specific creation of a new void entity (UndefinedEntity only)

    OwnCopyCase (me; CN : Integer;
    	         entfrom : IGESEntity; entto : mutable IGESEntity;
    	         TC : in out CopyTool);
    ---Purpose : Copies parameters which are specific of each Type of Entity

end DefaultGeneral;
