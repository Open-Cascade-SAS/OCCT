-- File:	Translation.cdl
-- Created:	Wed Aug 26 14:32:08 1992
-- Author:	Remi GILET
--		<reg@topsn3>
---Copyright:	 Matra Datavision 1992

class MakeTranslation

from gce

    ---Purpose: This class implements elementary construction algorithms for a
    -- translation in 3D space. The result is a gp_Trsf transformation.
    -- A MakeTranslation object provides a framework for:
    -- -   defining the construction of the transformation,
    -- -   implementing the construction algorithm, and
    -- -   consulting the result.

uses Pnt  from gp,
     Trsf from gp,
     Vec  from gp,
     Real from Standard
     
is

Create(Vect : Vec from gp) returns MakeTranslation;
    --- Purpose: Constructs a translation along the vector " Vect"
    
Create(Point1 : Pnt from gp;
       Point2 : Pnt from gp) returns MakeTranslation;
    ---Purpose: Constructs a translation along the vector
    --   (Point1,Point2) defined from the point Point1 to the point Point2.
        
Value(me) returns Trsf from gp
    is static;
    ---C++: return const&
    ---Purpose:
    -- Returns the constructed transformation.

Operator(me) returns Trsf from gp
    is static;
    ---C++: return const&
    ---C++: alias "Standard_EXPORT operator gp_Trsf() const;"

fields

    TheTranslation : Trsf from gp;

end MakeTranslation;

