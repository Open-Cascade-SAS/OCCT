-- Created on: 1993-01-11
-- Created by: CKY / Contract Toubro-Larsen ( Anand NATRAJAN )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Flow from IGESAppli  inherits IGESEntity

        ---Purpose: defines Flow, Type <402> Form <18>
        --          in package IGESAppli
        --          Represents a single signal or a single fluid flow path
        --          starting from a starting Connect Point Entity and
        --          including additional intermediate connect points.

uses

        ConnectPoint                 from IGESDraw,
        TextDisplayTemplate          from IGESGraph,
        HAsciiString                 from TCollection,
        HArray1OfHAsciiString        from Interface,
        HArray1OfIGESEntity          from IGESData,
        HArray1OfConnectPoint        from IGESDraw,
        HArray1OfTextDisplayTemplate from IGESGraph

raises OutOfRange

is

        Create returns mutable Flow;

        -- Specific Methods pertaining to the class

        Init (me                : mutable;
              nbContextFlags    : Integer;
              aFlowType         : Integer;
              aFuncFlag         : Integer;
              allFlowAssocs     : HArray1OfIGESEntity;
              allConnectPoints  : HArray1OfConnectPoint;
              allJoins          : HArray1OfIGESEntity;
              allFlowNames      : HArray1OfHAsciiString;
              allTextDisps      : HArray1OfTextDisplayTemplate;
              allContFlowAssocs : HArray1OfIGESEntity);
        ---Purpose : This method is used to set the fields of the class Flow
        --       - nbContextFlags    : Count of Context Flags, always = 2
        --       - aFlowType         : Type of Flow, default = 0
        --       - aFuncFlag         : Function Flag, default = 0
        --       - allFlowAssocs     : Flow Associativity Entities
        --       - allConnectPoints  : Connect Point Entities
        --       - allJoins          : Join Entities
        --       - allFlowNames      : Flow Names
        --       - allTextDisps      : Text Display Template Entities
        --       - allContFlowAssocs : Continuation Flow Associativity Entities

    	OwnCorrect (me : mutable) returns Boolean;
	---Purpose : forces NbContextFalgs to 2, returns True if changed

        NbContextFlags (me) returns Integer;
        ---Purpose : returns number of Count of Context Flags, always = 2

        NbFlowAssociativities (me) returns Integer;
        ---Purpose : returns number of Flow Associativity Entities

        NbConnectPoints (me) returns Integer;
        ---Purpose : returns number of Connect Point Entities

        NbJoins (me) returns Integer;
        ---Purpose : returns number of Join Entities

        NbFlowNames (me) returns Integer;
        ---Purpose : returns number of Flow Names

        NbTextDisplayTemplates (me) returns Integer;
        ---Purpose : returns number of Text Display Template Entities

        NbContFlowAssociativities (me) returns Integer;
        ---Purpose : returns number of Continuation Flow Associativity Entities

        TypeOfFlow (me) returns Integer;
        ---Purpose : returns Type of Flow = 0 : Not Specified (default)
        --                                  1 : Logical
        --                                  2 : Physical

        FunctionFlag (me) returns Integer;
        ---Purpose : returns Function Flag = 0 : Not Specified (default)
        --                                   1 : Electrical Signal
        --                                   2 : Fluid Flow Path

        FlowAssociativity (me; Index : Integer) returns IGESEntity
        raises OutOfRange;
        ---Purpose : returns Flow Associativity Entity
        -- raises exception if Index <= 0 or Index > NbFlowAssociativities()

        ConnectPoint (me; Index : Integer) returns ConnectPoint
        raises OutOfRange;
        ---Purpose : returns Connect Point Entity
        -- raises exception if Index <= 0 or Index > NbConnectPoints()

        Join (me; Index : Integer) returns IGESEntity
        raises OutOfRange;
        ---Purpose : returns Join Entity
        -- raises exception if Index <= 0 or Index > NbJoins()

        FlowName (me; Index : Integer) returns HAsciiString from TCollection
        raises OutOfRange;
        ---Purpose : returns Flow Name
        -- raises exception if Index <= 0 or Index > NbFlowNames()

        TextDisplayTemplate (me; Index : Integer) returns TextDisplayTemplate
        raises OutOfRange;
        ---Purpose : returns Text Display Template Entity
        -- raises exception if Index <= 0 or Index > NbTextDisplayTemplates()

        ContFlowAssociativity (me; Index : Integer) returns IGESEntity
        raises OutOfRange;
        ---Purpose : returns Continuation Flow Associativity Entity
        -- raises exception if Index <= 0 or Index > NbContFlowAssociativities()

fields

--
-- Class    : IGESAppli_Flow
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class Flow.
--
-- Reminder : A Flow instance is defined by :
--            - Count of Context Flags, always = 2
--            - Type of Flow, default = 0
--            - Function Flag, default = 0
--            - Flow Associativity Entities
--            - Connect Point Entities
--            - Join Entities
--            - Flow Names
--            - Text Display Template Entities
--            - Continuation Flow Associativity Entities

        theNbContextFlags          : Integer;
        theTypeOfFlow              : Integer;
        theFunctionFlag            : Integer;
        theFlowAssociativities     : HArray1OfIGESEntity;
        theConnectPoints           : HArray1OfConnectPoint;
        theJoins                   : HArray1OfIGESEntity;
        theFlowNames               : HArray1OfHAsciiString;
        theTextDisplayTemplates    : HArray1OfTextDisplayTemplate;
        theContFlowAssociativities : HArray1OfIGESEntity;

end Flow;
