-- Created on: 1991-10-04
-- Created by: Remi GILET
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class BPoint from GccInt  

inherits Bisec from GccInt 
     ---Purpose: Describes a point as a bisecting object between two 2D geometric objects.
        
uses Pnt2d from gp,
     IType  from GccInt


is

Create(Point : Pnt2d) returns mutable BPoint;
    ---Purpose: Constructs a bisecting object whose geometry is the 2D point Point.
    
Point(me) returns Pnt2d from gp
    is redefined;
    ---Purpose: Returns a 2D point which is the geometry of this bisecting object.
    
ArcType(me) returns IType from GccInt
    is static;
    --- Purpose: Returns GccInt_Pnt, which is the type of any GccInt_BPoint bisecting object.
    
fields

    pnt : Pnt2d from gp;
    ---Purpose: The bisecting line.

end BPoint;    

