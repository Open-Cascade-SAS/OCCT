-- Created on: 2003-03-20
-- Created by: Michael KLOKOV
-- Copyright (c) 2003-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


deferred class HistoryCollector from BOP inherits TShared from MMgt
uses
    Shape from TopoDS,
    Operation from BOP,
    ListOfShape from TopTools,
    DataMapOfShapeListOfShape from TopTools,
    PDSFiller from BOPTools

is
    Initialize;
    
    Initialize(theShape1   : Shape from TopoDS;
    	       theShape2   : Shape from TopoDS;
	       theOperation: Operation from BOP);

    Generated (me: mutable; S : Shape from TopoDS)
    	returns ListOfShape from TopTools
	is virtual;
    	---C++:  return const & 
	
    SetResult(me: mutable; theResult: Shape from TopoDS;
    	    	    	   theDSFiller: PDSFiller from BOPTools)
    	is virtual;

    Modified (me: mutable; S : Shape from TopoDS)
    	returns ListOfShape from TopTools
	is virtual;
	---C++:  return const & 

    IsDeleted (me: mutable; S : Shape from TopoDS)
    	returns Boolean from Standard
	is virtual;

    HasGenerated (me)
    	returns Boolean from Standard
	is virtual;

    HasModified (me)
    	returns Boolean from Standard
	is virtual;

    HasDeleted (me)
    	returns Boolean from Standard
	is virtual;

fields
    myEmptyList: ListOfShape from TopTools is protected;
    myOp      : Operation from BOP is protected;
    myGenMap  : DataMapOfShapeListOfShape from TopTools is protected;
    myModifMap: DataMapOfShapeListOfShape from TopTools is protected;
    myS1         : Shape from TopoDS is protected;
    myS2         : Shape from TopoDS is protected;
    myResult     : Shape from TopoDS is protected;
    myHasDeleted : Boolean from Standard is protected;

end HistoryCollector from BOP;
