-- Created on: 1993-01-14
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package TopTools 

	---Purpose: The  TopTools package provides   utilities for the
	--          topological data structure.
	--          
	--          * ShapeMapHasher. Hash a  Shape base on the TShape
	--          and the Location. The Orientation is not used.
	--          
	--          * OrientedShapeMapHasher. Hash a Shape base on the
	--          TShape ,the Location and the Orientation.
	--          
	--          * Instantiations of TCollection for Shapes :
	--             MapOfShape
	--             IndexedMapOfShape
	--             DataMapOfIntegerShape
	--             DataMapOfShapeInteger
	--             DataMapOfShapeReal
	--             Array1OfShape
	--             HArray1OfShape
	--             SequenceOfShape
	--             HSequenceOfShape
	--             ListOfShape
	--             Array1OfListShape
	--             HArray1OfListShape
	--             DataMapOfIntegerListOfShape
	--             DataMapOfShapeListOfShape
	--             DataMapOfShapeListOfInteger
	--             IndexedDataMapOfShapeShape
	--             IndexedDataMapOfShapeListOfShape
	--             DataMapOfShapeShape
	--             IndexedMapOfOrientedShape
	--             DataMapOfShapeSequenceOfShape
	--             IndexedDataMapOfShapeAddress
        --             DataMapOfOrientedShapeShape
	--             
	--          * LocationSet : to write sets of locations.
	--          
	--          * ShapeSet : to writes sets of TShapes.
	--          
	--          Package Methods :
	--          
	--            Dump : To dump the topology of a Shape.
	--          

        --- Level : Public  
        --  All methods of all  classes will be public.


uses

    MMgt,
    TCollection,
    TColStd,
    TopLoc,
    TopAbs,
    TopoDS,
    Message

is

    ----------------------------------------------------------
    -- TCollections for Shapes
    ----------------------------------------------------------

    class ShapeMapHasher;
    
    class OrientedShapeMapHasher;
    
    imported MapOfShape;
    
    imported MapIteratorOfMapOfShape;

    imported MapOfOrientedShape;

    imported MapIteratorOfMapOfOrientedShape;

    imported IndexedMapOfShape;
				    
    imported DataMapOfIntegerShape;
				    
    imported DataMapIteratorOfDataMapOfIntegerShape;
    
    imported DataMapOfOrientedShapeInteger;
    
    imported DataMapIteratorOfDataMapOfOrientedShapeInteger;

    imported DataMapOfShapeInteger;

    imported DataMapIteratorOfDataMapOfShapeInteger;

    imported DataMapOfShapeReal;

    imported DataMapIteratorOfDataMapOfShapeReal;

    imported Array1OfShape;
	
    imported transient class HArray1OfShape; 
				  
    imported Array2OfShape;
	
    imported transient class HArray2OfShape;			 
	
    imported SequenceOfShape;
	
    imported transient class HSequenceOfShape;
	
    imported ListOfShape;
	
    imported ListIteratorOfListOfShape;
	
    imported Array1OfListOfShape;
	
    imported transient class HArray1OfListOfShape;
	
    imported DataMapOfIntegerListOfShape;
	
    imported DataMapIteratorOfDataMapOfIntegerListOfShape;
	
    imported DataMapOfShapeListOfShape;
	
    imported DataMapIteratorOfDataMapOfShapeListOfShape;
				 
    imported DataMapOfShapeListOfInteger;
				 
    imported DataMapIteratorOfDataMapOfShapeListOfInteger;
				 
    imported IndexedDataMapOfShapeShape;				
    imported IndexedDataMapOfShapeListOfShape;
					
    imported DataMapOfShapeShape;
					
    imported DataMapIteratorOfDataMapOfShapeShape;

    imported IndexedMapOfOrientedShape;

    imported DataMapOfShapeSequenceOfShape;

    imported DataMapIteratorOfDataMapOfShapeSequenceOfShape;

    imported IndexedDataMapOfShapeAddress;	  

     imported DataMapOfOrientedShapeShape;

     imported DataMapIteratorOfDataMapOfOrientedShapeShape;			    

    ----------------------------------------------------------
    -- Tools for writing and reading Locations and Shapes
    ----------------------------------------------------------

    class LocationSet;
  
    pointer LocationSetPtr to LocationSet from TopTools;

    class ShapeSet;
	---Purpose: A set of Shapes. Can be dump, wrote or read.
	
    --
    --     Package methods
    --   

    imported MutexForShapeProvider;
    
    Dump(Sh : Shape from TopoDS; S : in out OStream);
	  ---Purpose: Dumps the topological structure  of <Sh>  on the
	  --          stream <S>.

    Dummy(I : Integer);
	---Purpose: This is to bypass an extraction bug. It will force
	--          the  inclusion    of  Standard_Integer.hxx  itself
	--          including Standard_OStream.hxx  at   the   correct
	--          position.
    
end TopTools;


