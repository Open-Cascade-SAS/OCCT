-- Created on: 1994-06-07
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class SurfaceIterator from TopOpeBRepDS 
    inherits InterferenceIterator from TopOpeBRepDS

uses

    State               from TopAbs,
    Orientation         from TopAbs,
    ListOfInterference  from TopOpeBRepDS
    
is
    Create(L : ListOfInterference from TopOpeBRepDS) 
    returns SurfaceIterator;
    ---Purpose: Creates an  iterator on the  Surfaces on solid
    --          described by the interferences in <L>.
    
    Current(me) returns Integer from Standard
    ---Purpose: Index of the surface in the data structure.
    is static;
    
    Orientation(me; S : State from TopAbs) 
    returns Orientation from TopAbs
    is static;
    
end SurfaceIterator from TopOpeBRepDS;
