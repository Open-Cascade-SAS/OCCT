-- Created on: 1993-03-23
-- Created by: BBL
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class Pixel from Aspect inherits Storable

	---Version: 0.0

	---Purpose: This class defines a Pixel.
	---Keywords:
	---Warning:
	---References:
is

	Initialize;
	---Level: Public

	Print( me ; s : in out OStream ) is deferred ;
	---Level: Public
	---Purpose : Prints the contents of <me> on the stream <s>
	---C++: alias "friend Standard_EXPORT Standard_OStream& operator << (Standard_OStream&,const Aspect_Pixel& );"

end Pixel from Aspect;
