-- Created on: 1995-01-23
-- Created by: Didier Piffault
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

--		Full Copy of Select_Rectangle (Didier Piffault 94)


class SortAlgo from SelectBasics 

	---Purpose: Quickly selection of a rectangle in a set of rectangles


uses    Integer from Standard,
    	Real    from Standard,
	MapIteratorOfMapOfInteger from TColStd,
	MapOfInteger from TColStd,
	ListIteratorOfListOfInteger from TColStd,
	Box2d          from Bnd,
	HArray1OfBox2d from Bnd,
	BoundSortBox2d from Bnd


is      Create 
	---Purpose: Empty rectangle selector.
	    returns SortAlgo from SelectBasics;

	Create     (ClippingRectangle    : Box2d from Bnd;
    	    	    sizeOfSensitiveArea  : Real from Standard;
    	    	    theRectangles        : HArray1OfBox2d from Bnd)
	---Purpose: Creates a initialized selector.
	    returns SortAlgo from SelectBasics;

	Initialize (me                   : in out;
    	    	    ClippingRectangle    : Box2d from Bnd;
    	    	    sizeOfSensitiveArea  : Real from Standard;
    	    	    theRectangles        : HArray1OfBox2d from Bnd)
	---Purpose: Clears and initializes the selector.
	    is static;


	InitSelect (me    : in out;
	    	    x, y  : Real from Standard) 
	---Purpose: Searchs the items on this position.
	    is static;


	InitSelect (me    : in out;
	    	    rect  : Box2d from Bnd) 
	---Purpose: Searchs the items in this rectangle.
	    is static;



    	More(me)
	---Purpose: Returns true if there is something selected.
	    returns Boolean from Standard is static;

    	Next(me : in out) 
	---Purpose: Sets value on the next selected item.
	    is static;

    	Value(me)
	---Purpose: Returns the index of the selected rectangle.
	    returns Integer from Standard is static;


fields  clipRect   : Box2d            from Bnd;
	sizeArea   : Real             from Standard;
	sortedRect : BoundSortBox2d   from Bnd;
	myMap      : MapOfInteger     from TColStd;
	curResult  : MapIteratorOfMapOfInteger from TColStd;

end SortAlgo;



