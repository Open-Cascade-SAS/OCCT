-- Created on: 1992-04-03
-- Created by: Laurent BUCHARD
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class IntersectionPoint from IntRes2d

    ---Purpose: Definition of an intersection point between two
    --          2D curves.


inherits Storable from Standard

uses Pnt2d      from gp,
     Transition from IntRes2d
is

    Create

	---Purpose: Empty constructor.

    	returns IntersectionPoint from IntRes2d;


    Create(P: Pnt2d from gp; Uc1,Uc2:Real from Standard;
           Trans1,Trans2: Transition from IntRes2d;
           ReversedFlag: Boolean from Standard)
	   
	---Purpose: Creates an IntersectionPoint.
	--          if ReversedFlag is False, the parameter Uc1(resp. Uc2)
	--          and the Transition Trans1 (resp. Trans2) refer to 
	--          the first curve (resp. second curve) otherwise Uc1 
	--          and Trans1 (resp. Uc2 and Trans2) refer to the 
	--          second curve (resp. the first curve).

      	---C++: inline	   

	returns IntersectionPoint from IntRes2d;
	

    SetValues(me:in out; P: Pnt2d from gp; Uc1,Uc2:Real from Standard;
              Trans1,Trans2: Transition from IntRes2d;
              ReversedFlag: Boolean from Standard)

	---Purpose: Sets the values for an existing intersection 
	--          point. The meaning of the parameters are the same 
	--          as for the Create.

	---C++: inline

	is static;



    Value(me)
    
    	---Purpose: Returns the value of the coordinates of the
    	--          intersection point in the 2D space.

	---C++: inline
	---C++: return const &

    	returns Pnt2d from gp
    	is static;


    ParamOnFirst(me)

    	---Purpose: Returns the parameter on the first curve.

	---C++: inline

    	returns Real from Standard
	is static;


    ParamOnSecond(me)

    	---Purpose: Returns the parameter on the second curve.

       	---C++: inline

    	returns Real from Standard
	is static;


    TransitionOfFirst(me)
    
    	---Purpose: Returns the transition of the 1st curve compared to
    	--          the 2nd one.

	---C++: inline
        ---C++: return const &
    	returns Transition from IntRes2d
	is static;


    TransitionOfSecond(me)
    
    	---Purpose: returns the transition of the 2nd curve compared to
    	--          the 1st one.

	---C++: inline
        ---C++: return const &
    	returns Transition from IntRes2d
	is static;


fields

    pt       : Pnt2d      from gp;
    p1       : Real       from Standard;
    p2       : Real       from Standard;
    trans1   : Transition from IntRes2d;
    trans2   : Transition from IntRes2d;

end IntersectionPoint;
 

