-- Created on: 1997-08-07
-- Created by: Jean-Louis Frenkel
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Session from CDF inherits Transient from Standard


uses
    Directory from CDF,
    ExtendedString from TCollection,
    Application from CDF, 
    MetaDataDriver from CDF, 
    Writer from PCDM
raises

    NoSuchObject from Standard,MultiplyDefined from Standard

is
    Create  returns Session from CDF
    raises MultiplyDefined from Standard;

    Exists(myclass)
--- Purpose: returns true if a session has been created.
    returns Boolean from Standard;
    
    CurrentSession(myclass) returns Session from CDF;
    ---Purpose: returns the only one instance of Session 
    --          that has been created.

    
    Directory(me) returns Directory from CDF;
    ---Purpose: returns the directory of the session;
    ---Level: Public 

    
---Category: current application management
    HasCurrentApplication(me) returns Boolean from Standard;
    
    CurrentApplication(me) returns Application from CDF
    raises NoSuchObject from Standard;
    
    SetCurrentApplication(me: mutable; anApplication: Application from CDF);
    
    UnsetCurrentApplication(me: mutable);


---Category: database related methods

    MetaDataDriver(me) returns MetaDataDriver from CDF
    raises NoSuchObject from Standard;
    
    
    LoadDriver(me: mutable);

fields

    myDirectory            : Directory from CDF;
    myCurrentApplication   : Application from CDF;
    myHasCurrentApplication: Boolean from Standard;
    myMetaDataDriver       : MetaDataDriver from CDF;
friends
    class Application from CDF
end Session from CDF;
