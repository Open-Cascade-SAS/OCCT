-- Created on: 1997-02-06
-- Created by: Kernel
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class TypeData from Storage 

inherits TShared from MMgt

uses HSequenceOfAsciiString from TColStd,
     PType from Storage,
     AsciiString from TCollection,
     Error from Storage
     
raises NoSuchObject from Standard
is
    Create returns mutable TypeData from Storage;
    
    NumberOfTypes(me) returns Integer from Standard;
    
    IsType(me; aName : AsciiString from TCollection) returns Boolean from Standard;
    
    Types(me) returns HSequenceOfAsciiString from TColStd;

    ErrorStatus(me) returns Error from Storage;
    ErrorStatusExtension(me) returns AsciiString from TCollection;
   
    ClearErrorStatus(me : mutable);

    Clear(me : mutable); 
	
    -- PRIVATE

    AddType(me : mutable; aName : AsciiString from TCollection; aTypeNum : Integer from Standard) is private;
    ---Purpose: add a type to the list
    
    Type(me; aTypeNum : Integer from Standard) returns AsciiString from TCollection
      raises NoSuchObject is private;
    ---Purpose: returns the name of the type with number <aTypeNum>
    
    Type(me; aTypeName : AsciiString from TCollection) returns Integer from Standard
      raises NoSuchObject is private;
    ---Purpose: returns the name of the type with number <aTypeNum>

    SetErrorStatus(me : mutable; anError : Error from Storage) is private;
    SetErrorStatusExtension(me : mutable; anErrorExt : AsciiString from TCollection) is private;    
    
    fields
    
      myPt                 : PType from Storage;      
      myErrorStatus        : Error from Storage;
      myErrorStatusExt     : AsciiString      from TCollection;
     
    friends class Schema from Storage
    
end;
