-- Created on: 1999-06-16
-- Created by: Sergey RUIN
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class RealArray from TDataStd inherits Attribute from TDF

	---Purpose: A framework for an attribute composed of a real number array.

uses  
     HArray1OfReal            from TColStd, 
     GUID                     from Standard,     
     Attribute                from TDF,
     Label                    from TDF, 
     DeltaOnModification      from TDF,
     RelocationTable          from TDF

is 

    ---Purpose: class methods
    --          =============

    GetID (myclass)   
       	---C++: return const & 
    	---Purpose: Returns the GUID for arrays of reals.  
    returns GUID from Standard;

    Set (myclass; label : Label from TDF; lower, upper : Integer from Standard; 
    	    	  isDelta : Boolean from Standard = Standard_False)
    	---Purpose: Finds or creates on the <label> a real array attribute 
        -- with the specified <lower> and <upper> boundaries.  
    	-- If attribute is already set, all input parameters are refused and the found
    	-- attribute is returned.
    returns RealArray from TDataStd;

    
    ---Category: RealArray methods
    --          ===============

    Init(me : mutable; lower, upper : Integer from Standard);
    ---Purpose: Initialize the inner array with bounds from <lower> to <upper>  

    SetValue (me : mutable; Index :Integer from Standard; Value : Real from Standard);
    ---Purpose: Sets  the   <Index>th  element  of   the  array to <Value>
    -- OutOfRange exception is raised if <Index> doesn't respect Lower and Upper bounds of the internal  array.

    Value (me; Index : Integer from Standard)
    ---Purpose: Return the value of  the  <Index>th element of the array
    --
    ---C++: alias operator ()
    returns Real from Standard;

    Lower (me) returns Integer from Standard;      
    ---Purpose:  Returns the lower boundary of the array.

    Upper (me) returns Integer from Standard;
    ---Purpose: Returns the upper boundary of the array.
    
    Length (me) returns Integer from Standard;    
    ---Purpose: Returns the number of elements of the array of reals
    --    in terms of the number of elements it contains.
    
    ChangeArray(me : mutable; newArray : HArray1OfReal from TColStd; 
    	    	    	      isCheckItems : Boolean = Standard_True); 	    
    	---Purpose: Sets the inner array <myValue> of the RealArray attribute  
    	-- to <newArray>. If value of <newArray> differs from <myValue>, 
    	-- Backup performed and myValue refers to new instance of HArray1OfReal 
    	-- that holds <newArray> values 
	-- If <isCheckItems> equal True each item of <newArray> will be checked with each 
    	-- item of <myValue> for coincidence (to avoid backup).
    
    Array(me) returns HArray1OfReal from TColStd;
    ---Purpose: Returns the handle of this array of reals.
    ---C++: inline 
    ---C++: return const 
     
    GetDelta(me) returns Boolean from Standard;  
    ---C++: inline  
    
    SetDelta(me : mutable; isDelta : Boolean from Standard);     
    ---C++: inline  
    ---Purpose: for  internal  use  only!  
     
    RemoveArray(me  : mutable) is private;      
    ---C++: inline      
    
    ---Category: methodes of TDF_Attribute
    --           =========================
    Create    
    returns RealArray from TDataStd; 
    
    ID (me)
    	---C++: return const & 
    returns GUID from Standard;

    Restore (me: mutable; With : Attribute from TDF);

    NewEmpty (me)
    returns Attribute from TDF;

    Paste (me; Into : Attribute from TDF;
	       RT   : RelocationTable from TDF);    
    ---Purpose: Note. Uses inside ChangeArray() method 
    
    Dump(me; anOS : in out OStream from Standard)
    	returns OStream from Standard
    	is redefined;
	---C++: return &

    ---Category: methods to be added for using in DeltaOnModification  
    --           =====================================================
    DeltaOnModification(me; anOldAttribute : Attribute from TDF)
    	returns DeltaOnModification from TDF
    	---Purpose : Makes a DeltaOnModification between <me> and
    	--         <anOldAttribute>.  
    	is redefined virtual;  
fields

    myValue : HArray1OfReal from TColStd;
    myIsDelta : Boolean from Standard; 
     
friends   

    class DeltaOnModificationOfRealArray from TDataStd  
     
end RealArray;
