-- Created on: 1999-02-11
-- Created by: Xuan PHAM PHU
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class makeTransition from TopOpeBRepTool
uses
    Pnt2d from gp,
    Edge from TopoDS,
    Face from TopoDS,
    State from TopAbs	        	
is    
	   
    Create returns makeTransition from TopOpeBRepTool;
    
    Initialize(me : in out; 
    	       E : Edge from TopoDS; pbef,paft,parE : Real;
    	       FS : Face from TopoDS; uv : Pnt2d from gp;
    	       factor : Real)
    returns Boolean;
    -- <E> interfers with <FS> at point :
    -- Pt(parE,E) = Pt(uv,FS)
    --  <pbef>,<paft> greater and lower <parE>.    

    Setfactor(me : in out; factor : Real); -- 0 < factor < 1
    Getfactor(me) returns Real;

    IsT2d(me) returns Boolean;  
	   
    SetRest(me : in out; 
    	    ES : Edge from TopoDS; parES : Real)
    returns Boolean;
    -- Pt(parES,ES) = Pt(uv,FS)
    --  Transition is computed vs <ES>, restrition on <FS>
    HasRest(me) returns Boolean;

    MkT2donE(me; stb,sta : out State from TopAbs)
    returns Boolean;  
    -- returns false if (!isT2d)   
    -- computes transition on <myE>, using tangent vectors. 

    MkT3onE(me; stb,sta : out State from TopAbs)
    returns Boolean;  
    -- returns false if (isT2d)
    -- return states in/out/on
    
    MkT3dproj(me; stb,sta : out State from TopAbs)
    returns Boolean;
    -- using projections.
    -- return states in/out/on
    
    MkTonE(me : in out; stb,sta : out State from TopAbs)
    returns Boolean;  
    -- Compute for <T> = transition on <E> vs <FS>.
    -- return states in/out/on.
    -- modifies field myfactor.

fields
    myE : Edge from TopoDS; 
    mypb,mypa,mypE : Real;
    myFS : Face from TopoDS;
    myuv : Pnt2d from gp;
    
    hasES : Boolean;
    myES : Edge from TopoDS;
    mypES : Real;

    isT2d : Boolean;	
    myfactor : Real;
	
end makeTransition;
