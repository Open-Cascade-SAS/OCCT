-- File:	Vrml_Group.cdl
-- Created:	Thu Mar 27 11:19:40 1997
-- Author:	Alexander BRIVIN and Dmitry TARASOV
--		<brivin@meteox.nizhny.matra-dtv.fr>
---Copyright:	 Matra Datavision 1997


class Group from Vrml 

	---Purpose: defines a Group node of VRML specifying group properties.
    	--  This node defines the base class for all group nodes. Group is a node that  
    	--  contains an ordered list of child nodes. This node is simply a container for  
    	--  the child nodes and does not alter the traversal state in any way.
	--  During traversal, state accumulated for a child is passed on to each successive  
    	--  child and then to the parents of the group (Group does not push or pop traversal  
    	--  state as separator does). 

is
    Create  returns   Group from Vrml;

    Print  ( me : in out;  anOStream: in out OStream from Standard)  
    	    returns OStream from Standard;
    ---C++:  return  & 

fields
 
    myFlagPrint      :  Boolean                 from Standard; 

end Group;
