-- Created by: DAUTRY Philippe
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

--      	------------

---Version:	0.0
--Version	Date		Purpose
--		0.0	Feb 10 1997	Creation


class Data from DDF inherits Drawable3D from Draw

	---Purpose : Encapsulates a data framework from TDF in a drawable object

uses

    Data        from TDF,
    Interpretor from Draw,
    Display     from Draw

is


    Create  (aDF : Data from TDF)
    returns Data from DDF;
    
    
    DrawOn (me; dis : in out Display);
    
    
    Copy (me) 
    returns Drawable3D from Draw
    is redefined;

	
    Dump (me; S : in out OStream) 
    is redefined;


    DataFramework (me : mutable; aDF : Data from TDF);


    DataFramework (me)
    returns Data from TDF;
    

    Whatis (me; I : in out Interpretor from Draw)
    is redefined;

	
fields

    myDF : Data from TDF;

end Data;


