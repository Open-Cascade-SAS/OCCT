-- Created on: 1993-01-09
-- Created by: CKY / Contract Toubro-Larsen ( Kiran )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class BSplineSurface from IGESGeom  inherits IGESEntity

        ---Purpose: defines IGESBSplineSurface, Type <128> Form <0-9>
        --          in package IGESGeom
        --          A parametric equation obtained by dividing two summations
        --          involving weights (which are real numbers), the control
        --          points, and B-Spline basis functions

uses

        Pnt           from gp,
        HArray1OfReal from TColStd,
        HArray2OfReal from TColStd,
        HArray2OfXYZ  from TColgp

raises   DimensionMismatch, OutOfRange

is

        Create returns mutable BSplineSurface;

        -- Specific Methods pertaining to the class

        Init (me                           : mutable;
              anIndexU, anIndexV           : Integer;
              aDegU, aDegV                 : Integer;
              aCloseU, aCloseV             : Boolean;
              aPolynom, aPeriodU, aPeriodV : Boolean;
              allKnotsU, allKnotsV         : HArray1OfReal;
              allWeights                   : HArray2OfReal;
              allPoles                     : HArray2OfXYZ;
              aUmin, aUmax, aVmin, aVmax   : Real)
        raises DimensionMismatch;
        ---Purpose : This method is used to set the fields of the class
        --           BSplineSurface
        --       - anIndexU             : Upper index of first sum
        --       - anIndexV             : Upper index of second sum
        --       - aDegU, aDegV         : Degrees of first and second sets
        --                                of basis functions
        --       - aCloseU, aCloseV     : 1 = Closed in U, V directions
        --                                0 = open in U, V directions
        --       - aPolynom             : 0 = Rational, 1 = polynomial
        --       - aPeriodU, aPeriodV   : 0 = Non periodic in U or V direction
        --                                1 = Periodic in U or V direction
        --       - allKnotsU, allKnotsV : Knots in U and V directions
        --       - allWeights           : Array of weights
        --       - allPoles             : XYZ coordinates of all control points
        --       - aUmin                : Starting value of U direction
        --       - aUmax                : Ending value of U direction
        --       - aVmin                : Starting value of V direction
        --       - aVmax                : Ending value of V direction
        -- raises exception if allWeights & allPoles are not of same size.

    	SetFormNumber (me : mutable; form : Integer) raises OutOfRange;
	---Purpose : Changes FormNumber (indicates the Shape of the Surface)
	--           Error if not in range [0-9]


        UpperIndexU(me) returns Integer;
        ---Purpose : returns the upper index of the first sum (U)

        UpperIndexV(me) returns Integer;
        ---Purpose : returns the upper index of the second sum (V)

        DegreeU(me) returns Integer;
        ---Purpose : returns degree of first set of basis functions

        DegreeV(me) returns Integer;
        ---Purpose : returns degree of second set of basis functions

        IsClosedU(me) returns Boolean;
        ---Purpose : True if closed in U direction else False

        IsClosedV(me) returns Boolean;
        ---Purpose : True if closed in V direction else False

        IsPolynomial(me; flag : Boolean = Standard_False) returns Boolean;
        ---Purpose : True if polynomial, False if rational
        --           <flag> False (D) : computed from Weights
        --           <flag> True : recorded

        IsPeriodicU(me) returns Boolean;
        ---Purpose : True if periodic in U direction else False

        IsPeriodicV(me) returns Boolean;
        ---Purpose : True if periodic in V direction else False

        NbKnotsU(me) returns Integer;
        ---Purpose : returns number of knots in U direction
        -- KnotsU are numbered from -DegreeU

        NbKnotsV(me) returns Integer;
        ---Purpose : returns number of knots in V direction
        -- KnotsV are numbered from -DegreeV

        KnotU(me; anIndex : Integer) returns Real
        raises OutOfRange;
        ---Purpose : returns the value of knot referred to by anIndex in U direction
        -- raises exception if
        --      anIndex < -DegreeU() or anIndex > (NbKnotsU() - DegreeU())

        KnotV(me; anIndex : Integer) returns Real
        raises OutOfRange;
        ---Purpose : returns the value of knot referred to by anIndex in V direction
        -- raises exception if
        --      anIndex < -DegreeV() or anIndex > (NbKnotsV() - DegreeV())

        NbPolesU(me) returns Integer;
        ---Purpose : returns number of poles in U direction

        NbPolesV(me) returns Integer;
        ---Purpose : returns number of poles in V direction

        Weight(me; anIndex1, anIndex2 : Integer) returns Real
        raises OutOfRange;
        ---Purpose : returns the weight referred to by anIndex1, anIndex2
        -- raises exception if anIndex1 <= 0 or anIndex1 > NbPolesU()
        --               or if anIndex2 <= 0 or anIndex2 > NbPolesV()

        Pole(me; anIndex1, anIndex2 : Integer) returns Pnt
        raises OutOfRange;
        ---Purpose : returns the control point referenced by anIndex1, anIndex2
        -- raises exception if anIndex1 <= 0 or anIndex1 > NbPolesU()
        --               or if anIndex2 <= 0 or anIndex2 > NbPolesV()

        TransformedPole(me; anIndex1, anIndex2 : Integer) returns Pnt
        raises OutOfRange;
        ---Purpose : returns the control point referenced by anIndex1, anIndex2
        -- after applying the Transf.Matrix
        -- raises exception if anIndex1 <= 0 or anIndex1 > NbPolesU()
        --               or if anIndex2 <= 0 or anIndex2 > NbPolesV()

        UMin(me) returns Real;
        ---Purpose : returns starting value in the U direction

        UMax(me) returns Real;
        ---Purpose : returns ending value in the U direction

        VMin(me) returns Real;
        ---Purpose : returns starting value in the V direction

        VMax(me) returns Real;
        ---Purpose : returns ending value in the V direction

fields

--
-- Class    : IGESGeom_BSplineSurface
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class BSplineSurface.
--
-- Reminder : A BSplineSurface instance is defined by :
--            A parametric equation obtained by dividing two summations
--            involving weights (which are real numbers), the control
--            points, and B-Spline basis functions

        theIndexU     : Integer;
        theIndexV     : Integer;
        theDegreeU    : Integer;
        theDegreeV    : Integer;
        isClosedU     : Boolean;
        isClosedV     : Boolean;
        isPolynomial  : Boolean;
        isPeriodicU   : Boolean;
        isPeriodicV   : Boolean;
        theKnotsU     : HArray1OfReal;
        theKnotsV     : HArray1OfReal;
        theWeights    : HArray2OfReal;
        thePoles      : HArray2OfXYZ;
        theUmin       : Real;  -- Starting value for 1st parameter direction
        theUmax       : Real;  -- Ending   value for 1st parameter direction
        theVmin       : Real;  -- Starting value for 2nd parameter direction
        theVmax       : Real;  -- Ending   value for 2nd parameter direction

end BSplineSurface;
