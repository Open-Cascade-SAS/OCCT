-- Created on: 1994-08-24
-- Created by: Gilles DEBARBOUILLE
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class VariableGroup from Dynamic

inherits

    Variable from Dynamic
    
	---Purpose: This   inherited  class   from   variable is   for
	--          specifing  that the variable  does not accept only
	--          one   value    but a  collection   of  homogeneous
	--          values. This class is for describing the signature
	--          of the method definition. When an instance of this
	--          kind   of   method    is     done,    it   is    a
	--          CompositVariableInstance which is used.


is

    Create returns mutable VariableGroup from Dynamic;
    
    ---Level: Advanced 
    
    ---Purpose: Creates and Returns a new instance of this class.
    

end VariableGroup;
