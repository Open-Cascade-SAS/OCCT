-- Created on: 1991-10-23
-- Created by: Denis PASCAL
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


generic class SortedStrgCmptsIterator from GraphTools
             (Graph      as any;
    	      Vertex     as any;
	      GIterator  as any;
	      SSCIterator as any)

--generic class SortedStrgCmptsIterator from GraphTools
--            (Graph     as any;
--    	       Vertex    as any;
--	       GIterator as GraphIterator  (Graph,Vertex))
--	       SSCIterator as  SortedStrgCmptsFromIterator

    ---Purposes: This     generic    class        implements       the
    --           SortedStrgCptsFromIterator  with all  vertices of <G>
    --           reached by the Tool GIterator.
     
raises NoMoreObject from Standard,
       NoSuchObject from Standard
    
is


    Create 
    returns SortedStrgCmptsIterator from GraphTools;
	---Purpose: Create an empty algorithm.
    
    Create (G : Graph) 	
    	---Purpose: Create the   algorithm setting each vertex  of <G>
	--          reached by  GIterator tool, as initial conditions.
	--          Use Perform   method before visting  the result of
	--          the algorithm.
    returns SortedStrgCmptsIterator from GraphTools;
    
    FromGraph (me : in out; G : Graph);	
    	---Purpose: Add each vertex of <G>  reached by GIterator  tool
	--          as   initial  conditions.   Use  Perform  method
	--          before   visiting the  result  of   the algorithm.
        ---Level: Public 
    
    FromVertex (me : in out; V : Vertex);	
    	---Purpose: Add  <V>  as  initial  condition.  This method  is
	--          cumulative.  Use Perform method before visting the
	--          result of the algorithm.  
	---Level: Public

    Reset (me : in out);	
    	---Purpose: Reset the algorithm.  It may   be reused with  new
    	--          initial conditions.  
        ---Level: Public

    Perform (me : in out; G : Graph);
       ---Purpose: Peform the  algorithm  in  <G> from initial  setted
       --          conditions.  
       ---Level: Public
    
    More(me) returns Boolean from Standard;
        ---Purpose: returns  True   if  there are   others  strong
        --          components.
       ---Level: Public

    Next(me : in out) 
        ---Purpose: Set the iterator to the next strong component.
       ---Level: Public
    raises NoMoreObject from Standard;

    NbVertices (me) returns Integer from Standard
	---Purpose: Returns number  of vertices of  the current Strong
	--          Components.
       ---Level: Public
    raises NoSuchObject from Standard;

    Value(me; I : Integer from Standard) 
    returns any Vertex
	---Purpose: returns  the vertex of  index <I> of  the  current
	--          Strong Component.
	---C++: return const &
       ---Level: Public
    raises NoSuchObject from Standard;

fields

    myIterator : SSCIterator;
    
end SortedStrgCmptsIterator;
















    
