-- Created on: 1993-11-04
-- Created by: Christian CAILLET
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class BasicDumper  from IFSelect  inherits SessionDumper

    ---Purpose : BasicDumper takes into account, for SessionFile, all the
    --           classes defined in the package IFSelect : Selections,
    --           Dispatches (there is no Modifier)

uses Transient, AsciiString from TCollection, SessionFile

is

    Create returns mutable BasicDumper;
    ---Purpose : Creates a BasicDumper and puts it into the Library of Dumper

    WriteOwn (me; file : in out SessionFile; item : Transient) returns Boolean;
    ---Purpose : Write the Own Parameters of Types defined in package IFSelect
    --           Returns True if <item> has been processed, False else

    ReadOwn  (me; file : in out SessionFile;
    	    type : AsciiString from TCollection; item : out mutable Transient)
    	returns Boolean;
    ---Purpose : Recognizes and Read Own Parameters for Types of package
    --           IFSelect. Returns True if done and <item> created, False else

end BasicDumper;
