-- File:	RWStepFEA_RWFeaShellBendingStiffness.cdl
-- Created:	Thu Dec 12 17:51:06 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWFeaShellBendingStiffness from RWStepFEA

    ---Purpose: Read & Write tool for FeaShellBendingStiffness

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    FeaShellBendingStiffness from StepFEA

is
    Create returns RWFeaShellBendingStiffness from RWStepFEA;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : FeaShellBendingStiffness from StepFEA);
	---Purpose: Reads FeaShellBendingStiffness

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: FeaShellBendingStiffness from StepFEA);
	---Purpose: Writes FeaShellBendingStiffness

    Share (me; ent : FeaShellBendingStiffness from StepFEA;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWFeaShellBendingStiffness;
