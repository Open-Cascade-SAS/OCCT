-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class AutoDesignPersonAndOrganizationAssignment from StepAP214

inherits PersonAndOrganizationAssignment from StepBasic 

uses

	HArray1OfAutoDesignGeneralOrgItem from StepAP214, 
	AutoDesignGeneralOrgItem from StepAP214, 
	PersonAndOrganization from StepBasic, 
	PersonAndOrganizationRole from StepBasic
is

	Create returns mutable AutoDesignPersonAndOrganizationAssignment;
	---Purpose: Returns a AutoDesignPersonAndOrganizationAssignment


	Init (me : mutable;
	      aAssignedPersonAndOrganization : mutable PersonAndOrganization from StepBasic;
	      aRole : mutable PersonAndOrganizationRole from StepBasic) is redefined;

	Init (me : mutable;
	      aAssignedPersonAndOrganization : mutable PersonAndOrganization from StepBasic;
	      aRole : mutable PersonAndOrganizationRole from StepBasic;
	      aItems : mutable HArray1OfAutoDesignGeneralOrgItem from StepAP214) is virtual;

	-- Specific Methods for Field Data Access --

	SetItems(me : mutable; aItems : mutable HArray1OfAutoDesignGeneralOrgItem);
	Items (me) returns mutable HArray1OfAutoDesignGeneralOrgItem;
	ItemsValue (me; num : Integer) returns AutoDesignGeneralOrgItem;
	NbItems (me) returns Integer;

fields

	items : HArray1OfAutoDesignGeneralOrgItem from StepAP214; -- a SelectType

end AutoDesignPersonAndOrganizationAssignment;
