-- Created on: 2007-05-29
-- Created by: Vlad Romashko
-- Copyright (c) 2007-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ReferenceArray from TDataStd inherits Attribute from TDF

    ---Purpose: Contains an array of references to the labels.

uses 

    Attribute from TDF,
    GUID from Standard,
    Label from TDF,
    DataSet from TDF,
    RelocationTable from TDF,
    HLabelArray1 from TDataStd

is 

    ---Purpose: Static methods
    --          ==============

    GetID (myclass)   
    ---C++: return const & 
    ---Purpose: Returns the ID of the array of references (labels) attribute.
    returns GUID from Standard;

    Set (myclass; 
    	 label : Label from TDF; 
    	 lower, upper : Integer from Standard)
    ---Purpose: Finds or creates an array of reference values (labels) attribute.
    returns ReferenceArray from TDataStd;

    
    ---Category: ReferenceArray methods
    --           ======================
    
    Init (me : mutable; 
    	  lower, upper : Integer from Standard);
    ---Purpose: Initialize the inner array with bounds from <lower> to <upper>  

    SetValue (me : mutable; 
    	      index :Integer from Standard; 
    	      value : Label from TDF);
    ---Purpose: Sets the <Index>th element of the array to <Value>
    -- OutOfRange exception is raised if <Index> doesn't respect Lower and Upper bounds of the internal  array.

    Value (me; 
    	   Index : Integer from Standard)
    ---Purpose: Returns the value of the <Index>th element of the array.
    ---C++: alias operator ()
    returns Label from TDF;

    Lower (me) 
    ---Purpose: Returns the lower boundary of the array.
    returns Integer from Standard;      

    Upper (me) 
    ---Purpose: Returns the upper boundary of the array.
    returns Integer from Standard;
    
    Length (me) 
    ---Purpose: Returns the number of elements in the array.
    returns Integer from Standard;    

    
    ---Category: Advanced area
    --           =============

    InternalArray (me)
    ---C++: return const &
    returns HLabelArray1 from TDataStd;
    
    SetInternalArray (me : mutable;
    	    	      values : HLabelArray1 from TDataStd;
		      isCheckItems : Boolean = Standard_True);


    ---Category: Methodes of TDF_Attribute
    --           =========================
    
    Create
    returns mutable ReferenceArray from TDataStd; 

    ID (me)
    ---C++: return const & 
    returns GUID from Standard;

    Restore (me: mutable; With : Attribute from TDF);

    NewEmpty (me)
    returns mutable Attribute from TDF;

    Paste (me; Into : mutable Attribute from TDF;
	       RT   : mutable RelocationTable from TDF);    

    References (me; DS : DataSet from TDF) 
    is redefined;
    
    Dump(me; anOS : in out OStream from Standard)
    returns OStream from Standard
    is redefined;
    ---C++: return &


fields

    myArray : HLabelArray1 from TDataStd;


end ReferenceArray;
