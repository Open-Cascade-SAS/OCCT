-- Created on: 1992-11-18
-- Created by: Remi LEQUETTE
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package BRepClass 

	---Purpose: The  BRepClass packages provides    classification
	--          algorithms for the BRep topology.  It instantiates
	--          the algorithms from the package TopClass.

uses
    gp,
    TopAbs,
    TopoDS,
    TopExp,
    BRepTools,
    Geom2dInt,
    TopClass,
---    IntCurveSurface,
    Bnd




is
    class Edge;
	---Purpose: Stores the Edge and the Face.

    class Intersector;
	---Purpose: Intersect an Edge  with a segment.   This class is
	--          inherited   from   IntConicCurveOfGInter      from
	--          Geom2dInt.

    class FacePassiveClassifier instantiates Classifier2d from TopClass
    	(Edge         from BRepClass,
	 Intersector  from BRepClass);

    class FaceExplorer;
	---Purpose: Exploration of a Face to return UV edges.

    class FClassifier instantiates FaceClassifier from TopClass
    	(FaceExplorer from BRepClass,
	 Edge         from BRepClass,
	 Intersector  from BRepClass);
	 
    class FaceClassifier;
	---Purpose: Inherited    from   FClassifier   to   provide   a
	--          Constructor with a Face.

       
end BRepClass;
