-- Created on: 1998-08-04
-- Created by: Christian CAILLET
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class AutoDesignDocumentReference  from StepAP214    inherits DocumentReference

    -- introduced in STEP214 CC2

uses
     Document from StepBasic,
     HAsciiString from TCollection,
     AutoDesignReferencingItem from StepAP214,
     HArray1OfAutoDesignReferencingItem from StepAP214

is

    Create returns AutoDesignDocumentReference;

    Init (me : mutable;
           aAssignedDocument : Document;
           aSource : HAsciiString;
    	   aItems  : HArray1OfAutoDesignReferencingItem);

    Items (me) returns HArray1OfAutoDesignReferencingItem;
    SetItems (me : mutable; aItems : HArray1OfAutoDesignReferencingItem);
    ItemsValue (me; num : Integer) returns AutoDesignReferencingItem;
    NbItems (me) returns Integer;

fields

    items : HArray1OfAutoDesignReferencingItem;

end AutoDesignDocumentReference;
