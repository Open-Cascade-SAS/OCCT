-- Created on: 1993-07-06
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class CurveOnSurface from PBRep inherits GCurve from PBRep

	---Purpose: Representation  of a  curve   by a   curve  in the
	--          parametric space of a surface.

uses
    Curve    from PGeom2d,
    Surface  from PGeom,
    Pnt2d    from gp,
    Location from PTopLoc

is

    Create(PC : Curve    from PGeom2d;
    	   CF : Real     from Standard;
	   CL : Real     from Standard;
    	   S  : Surface  from PGeom; 
    	   L  : Location from PTopLoc)
    returns mutable CurveOnSurface from PBRep;
    	---Purpose: CF is curve first parameter
    	--          CL is curve last parameter
    	--          As far as they can't be computed from a Persistent Curve
    	--          they are given in the CurveOnSurface constructor

    Surface(me) returns  Surface from PGeom
    is static;
    	---Level: Internal 

    PCurve(me) returns  Curve from PGeom2d
    is static;
    	---Level: Internal 

    IsCurveOnSurface(me) returns Boolean
	---Purpose: Returns True.
    is redefined;
    
    SetUVPoints(me : mutable; Pnt1, Pnt2 : Pnt2d from gp);
    
    FirstUV(me) returns Pnt2d from gp;

    LastUV(me) returns Pnt2d from gp;
    
fields
    
    myPCurve      : Curve   from PGeom2d;
    mySurface     : Surface from PGeom;
    myUV1         : Pnt2d   from gp;
    myUV2         : Pnt2d   from gp;
    
end CurveOnSurface;
