-- Created on: 2002-12-10
-- Created by: data exchange team
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V2.0

class MeasureOrUnspecifiedValue from StepElement inherits SelectType from StepData

    ---Purpose: Representation of STEP SELECT type MeasureOrUnspecifiedValue

uses
    SelectMember from StepData,
    UnspecifiedValue from StepElement

is
    Create returns MeasureOrUnspecifiedValue from StepElement;
	---Purpose: Empty constructor

    CaseNum (me; ent: Transient) returns Integer;
	---Purpose: Recognizes a kind of MeasureOrUnspecifiedValue select type
	--          return 0 

    CaseMem (me; ent: SelectMember from StepData) returns Integer is redefined;
	---Purpose: Recognizes a items of select member MeasureOrUnspecifiedValueMember
	--          1 -> ContextDependentMeasure
	--          2 -> UnspecifiedValue
	--          0 else


     NewMember(me) returns SelectMember from StepData is redefined;
	---Purpose: Returns a new select member the type MeasureOrUnspecifiedValueMember

    SetContextDependentMeasure(me: in out; aVal :Real);
	---Purpose: Set Value for ContextDependentMeasure

    ContextDependentMeasure (me) returns Real;
	---Purpose: Returns Value as ContextDependentMeasure (or Null if another type)

    SetUnspecifiedValue(me: in out; aVal :UnspecifiedValue from StepElement);
	---Purpose: Set Value for UnspecifiedValue

    UnspecifiedValue (me) returns UnspecifiedValue from StepElement;
	---Purpose: Returns Value as UnspecifiedValue (or Null if another type)

end MeasureOrUnspecifiedValue;
