-- Created on: 1992-03-06
-- Created by: Isabelle GRIGNON
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

generic class Iterator from IntWalk (Point as any)
                       

	---Purpose: Template class to describe the exploration argument of the
	--          generic class IWalking 


raises OutOfRange from Standard

is

    Create
    
    	returns Iterator from IntWalk;


    Length(me)
    
    	---Purpose: returns the dimension of the exploration

    	returns Integer from Standard

    	is static;


    Value(me; Index : Integer)
    
    	---Purpose: returns the current point
    	--          an exception is raised if i>NbPoints

    	returns  Point

    	raises OutOfRange from Standard

    	is static;


    Append(me: in out; P: Point)
    
	---Purpose: Adds a point in the iterator.
    
    	is static;
	
	
end Iterator;
