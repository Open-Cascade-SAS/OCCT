-- Created on: 1993-06-03
-- Created by: Jean-Louis FRENKEL
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class LengthPresentation from DsgPrs
    	---Purpose: Framework for displaying lengths.
    	-- The length displayed is indicated by line segments
    	-- and text alone or by a combination of line segment,
    	-- text and   arrows at either or both of its ends.
uses
    Presentation from Prs3d,
    Pnt from gp,
    Dir from gp,
    Drawer from Prs3d,
    ExtendedString from TCollection,
    ArrowSide from DsgPrs,
    
    Pln from gp,
    Surface from Geom
is  
    Add( myclass; aPresentation: Presentation from Prs3d;
    	    	  aDrawer: Drawer from Prs3d;
		  aText: ExtendedString from TCollection;
                  AttachmentPoint1: Pnt from gp;
		  AttachmentPoint2: Pnt from gp;
		  aDirection: Dir from gp;
		  OffsetPoint: Pnt from gp);
	---Purpose: Draws a line segment representing a length in the
    	-- display aPresentation.
    	-- This segment joins the points AttachmentPoint1 and
    	-- AttachmentPoint2, along the direction aDirection.
    	-- The text aText will be displayed at the offset point OffsetPoint.
    	-- The line and text attributes are specified by the
    	-- attribute manager aDrawer.
        
    Add( myclass; aPresentation    : Presentation   from Prs3d;
    	    	  aDrawer          : Drawer         from Prs3d;
		  aText            : ExtendedString from TCollection;
                  AttachmentPoint1 : Pnt            from gp;
		  AttachmentPoint2 : Pnt            from gp;
		  aDirection       : Dir            from gp;
		  OffsetPoint      : Pnt            from gp;
	    	  ArrowSide        : ArrowSide      from DsgPrs );
	---Purpose: Draws a line segment representing a length in the
    	-- display aPresentation.
    	-- This segment joins the points AttachmentPoint1 and
    	-- AttachmentPoint2, along the direction aDirection.
    	-- The text aText will be displayed at the offset point
    	-- OffsetPoint. The value of the enumeration ArrowSide
    	-- controls whether arrows will be displayed at either or
    	-- both ends of the length.
    	-- The line, text and arrow attributes are specified by the
    	-- attribute manager aDrawer.
		   
    Add( myclass; aPresentation    : Presentation   from Prs3d;
    	    	  aDrawer          : Drawer         from Prs3d;
		  aText            : ExtendedString from TCollection;
                  AttachmentPoint1 : Pnt            from gp;
		  AttachmentPoint2 : Pnt            from gp;
		  PlaneOfFaces     : Pln            from gp;
		  aDirection       : Dir            from gp;
		  OffsetPoint      : Pnt            from gp;
	    	  ArrowSide        : ArrowSide      from DsgPrs );
	---Purpose: Draws a line segment representing a length in the
    	-- display aPresentation.
    	-- This segment joins the points AttachmentPoint1 and
    	-- AttachmentPoint2, along the direction aDirection.
    	-- The text aText will be displayed at the offset point
    	-- OffsetPoint. The value of the enumeration ArrowSide
    	-- controls whether arrows will be displayed at either or
    	-- both ends of the length.
    	-- The plane PlaneOfFaces is used if length is null.
    	-- The line, text and arrow attributes are specified by the
    	-- attribute manager aDrawer.
		   
    Add( myclass; aPresentation    : Presentation   from Prs3d;
    	    	  aDrawer          : Drawer         from Prs3d;
		  aText            : ExtendedString from TCollection;
		  SecondSurf       : Surface        from Geom;
                  AttachmentPoint1 : Pnt            from gp;
		  AttachmentPoint2 : Pnt            from gp;
		  aDirection       : Dir            from gp;
		  OffsetPoint      : Pnt            from gp;
	    	  ArrowSide        : ArrowSide      from DsgPrs );
	---Purpose: Draws a line segment representing a length in the
    	-- display aPresentation.
    	-- This segment joins the points AttachmentPoint1 and
    	-- AttachmentPoint2, along the direction
    	-- aDirection.   AttachmentPoint2 lies on the curvilinear
    	-- faces SecondSurf. The text aText will be displayed at
    	-- the offset point OffsetPoint. The value of the
    	-- enumeration ArrowSide controls whether arrows will
    	-- be displayed at either or both ends of the length.
    	-- The line, text and arrow attributes are specified by the
    	-- attribute manager aDrawer.


    Add(myclass;
    	aPresentation: Presentation from Prs3d;
    	aDrawer      : Drawer from Prs3d;
	Pt1          : Pnt from gp;
	Pt2          : Pnt from gp;
	ArrowSide    : ArrowSide from DsgPrs);
	---Purpose: Draws a line segment representing a length in the
    	-- display aPresentation.
    	-- This segment joins the points AttachmentPoint1 and
    	-- AttachmentPoint2, along the direction aDirection.
    	-- The value of the enumeration ArrowSide controls
    	-- whether arrows will be displayed at either or both ends of the length.
    	-- The line and arrow attributes are specified by the attribute manager aDrawer.

end LengthPresentation;
