-- Created on: 1992-10-01
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class InteriorPointTool from IntSurf 

	---Purpose: This class provides a tool on the "interior point"
	--          that can be used to instantiates the Walking
	--          algorithmes (see package IntWalk).

uses Pnt           from gp,
     Vec           from gp,
     Dir2d         from gp,
     InteriorPoint from IntSurf


is


    Value3d(myclass; PStart: InteriorPoint from IntSurf)
    
      	---Purpose: Returns the 3d coordinates of the starting point.

    	returns Pnt from gp;

	---C++: inline


    Value2d(myclass; PStart: InteriorPoint from IntSurf;
                         U, V: out Real from Standard);
    
	---Purpose: Returns the <U,V> parameters which are associated 
	--          with <P>
	--          it's the parameters which start the marching algorithm

	---C++: inline


    Direction3d(myclass; PStart: InteriorPoint from IntSurf)
    
        ---Purpose: returns the tangent at the intersectin in 3d space
        --          associated to <P>

    	returns Vec from gp;

	---C++: inline


    Direction2d(myclass; PStart: InteriorPoint from IntSurf)
    
        ---Purpose: returns the tangent at the intersectin in the
        --          parametric space of the parametrized surface.This tangent
        --          is associated to the value2d

    	returns Dir2d from gp;

	---C++: inline


end InteriorPointTool;
