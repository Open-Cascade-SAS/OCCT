-- Created on: 1998-10-20
-- Created by: DCB
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


private class BMPAlienData from AlienImage inherits AlienImageData from AlienImage

uses
  File                    from OSD,
  GenericColorMap         from Aspect,
  PseudoColorImage        from Image,
  ColorImage              from Image,
  Image                   from Image

raises
  OutOfRange      from Standard,
  TypeMismatch    from Standard

is
  Create returns mutable BMPAlienData from AlienImage ;

  Clear( me : in out mutable );
  ---Level: Public
  ---Purpose: Frees memory allocated by BMPAlienData
  ---C++: alias ~

  Read ( me : in out mutable ; afile : in out File from OSD )
  returns Boolean from Standard;
  ---Level: Public
  ---Purpose: Read content of a  BMPAlienData object from a file
  --          Returns True if file is a BMP file .

  Write( me : in immutable; afile : in out File from OSD )
  returns Boolean from Standard;
  ---Level: Public
  ---Purpose: Write content of a  BMPAlienData object to a file

  ToImage( me : in  immutable) 
  returns mutable Image from Image 
  raises TypeMismatch from Standard ;
  ---Level: Public
  ---Purpose : convert a BMPAlienData object to a Image object.

  FromImage( me : in out mutable ; anImage : in Image from Image )
  raises TypeMismatch from Standard ;
  ---Level: Public
  ---Purpose : convert a Image object to a BMPAlienData object.

  ------------------------------------------------------
  --- Private methods
  ------------------------------------------------------
  FromPseudoColorImage (me      : in out mutable; 
                        anImage : in PseudoColorImage from Image )
  is private;
  ---Level: Internal
  ---Purpose : convert a Image object to a GIFAlienData object.

  FromColorImage (me      : in out mutable;
                  anImage : in ColorImage from Image)
  is private;
  ---Level: Internal
  ---Purpose : convert a Image object to a GIFAlienData object.

fields
  myColorMap           : GenericColorMap from Aspect;
  myData               : Address         from Standard; --BYTE* or DWORD*
  myWidth              : Integer         from Standard;
  myHeight             : Integer         from Standard;

end;
 
