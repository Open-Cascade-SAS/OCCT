-- Created on: 1994-09-02
-- Created by: Yves FRICAUD
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class AnalyticCurInf from LProp 

	---Purpose: Computes the locals extremas of curvature of a gp curve
	--          Remark : a gp curve has not inflection.

uses
    CurveType from GeomAbs,
    CurAndInf from LProp
is
    Create;
    
    Perform (me     : in out; 
    	     T      :        CurveType from GeomAbs ;
             UFirst :        Real      from Standard ;
	     ULast  :        Real      from Standard ;
             Result : in out CurAndInf from LProp) 
    is static;
    
end AnalyticCurInf;
