-- Created on: 1992-06-04
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class CurveTool from Geom2dGcc

	---Purpose: 

uses Curve from Geom2dAdaptor,
     Pnt2d from gp,
     Vec2d from gp

is

    FirstParameter(myclass; C: Curve from Geom2dAdaptor)
    	returns Real;

    LastParameter(myclass; C: Curve from Geom2dAdaptor)
    	returns Real;

    EpsX (myclass                           ; 
    	  C       : Curve from Geom2dAdaptor;
    	  Tol     : Real  from Standard     )
    	returns Real;

    NbSamples(myclass                    ;
    	      C       : Curve from Geom2dAdaptor)
    	returns Integer;

    Value (myclass; C: Curve from Geom2dAdaptor; X: Real)
    	returns Pnt2d from gp;

    D1 (myclass; C: Curve from Geom2dAdaptor; U: Real ; 
                 P: out Pnt2d; T: out Vec2d);

    D2 (myclass; C: Curve from Geom2dAdaptor; U: Real ; 
                 P: out Pnt2d; T,N: out Vec2d);

    D3 (myclass; C: Curve from Geom2dAdaptor; U: Real ; 
                 P: out Pnt2d; T,N,dN: out Vec2d);

end CurveTool;

