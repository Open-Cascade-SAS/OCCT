-- File:        CompositeTextWithExtent.cdl
-- Created:     Mon Dec  4 12:02:24 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWCompositeTextWithExtent from RWStepVisual

	---Purpose : Read & Write Module for CompositeTextWithExtent

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     CompositeTextWithExtent from StepVisual,
     EntityIterator from Interface

is

	Create returns RWCompositeTextWithExtent;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable CompositeTextWithExtent from StepVisual);

	WriteStep (me; SW : in out StepWriter; ent : CompositeTextWithExtent from StepVisual);

	Share(me; ent : CompositeTextWithExtent from StepVisual; iter : in out EntityIterator);

end RWCompositeTextWithExtent;
