-- Created on: 1992-01-15
-- Created by: GG
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Modified:    FMN - 24/12/97 -> Suppression GEOMLITE
--              CQO - 24/12/97 -> BUC50037
--              stt:25-02-98; S3558: ajout IfManageStandardEvent
--              stt:08-04-98; suppr IfManageStandardEvent
--              CAL - 18/08/98 -> S3892. Ajout grilles 3d.
--              BGN - 16-09-98; Points d'entree du Triedre (S3819, Phase 1)
--              22-09-98 ; BGN : S3989 (anciennement S3819)
--                               TypeOfTriedron* from Aspect(et pas V3d)
--              CAL - 21/10/98 -> Speciale. Ajout methode Tumble.
--              29-OCT-98 : DCB : Adding ScreenCopy () method.
--      GG - 10/11/99 : PRO19603 Adding Redraw( area ) method
--      GG - 15/12/99 : GER61351 Adding SetBackgroundColor()
--                   and    BackgroundColor() methods
--      GG - 24/01/00 : -> Remove internal PixToRef() method, use Convert()
--                method instead.
--              -> Rename internal RefToPix() to Convert() method.
--              -> Add ConvertToGrid() methods,
--                 the Compute() internal method become private.
--              -> Add SetProjModel() method.
--      VKH - 15/11/99 : G004
--              -> Add method Dump()
--      THA  - 17/08/00 Thomas HARTL <t-hartl@muenchen.matra-dtv.fr>
--              -> Add Print method (works only under Windows).
--      GG  - IMP231100
--              -> Add IsActiveLight() & IsActivePlane() methods
--      SZV - IMP100701
--              -> Add ToPixMap() method
--              GG - RIC120302 Add NEW SetWindow method.
--              SAV - 22/10/01
--                              -> Add EnableDepthTest() & IsDepthTestEnabled().
--              VSV - 28/05/02: ZBUFFER mode of Trihedron
--              SAV - 23/12/02  -> Added methods to set background image
--              NKV - 23/07/07  -> Define custom projection and model view matrixes
--              NKV - 08/02/07  -> Add ConvertWithProj() method

class View from V3d inherits TShared from MMgt

        ---Purpose: Defines the application object VIEW for the
        --          VIEWER application.
        --          The methods of this class allow the editing
        --          and inquiring the parameters linked to the view.
        --          (Projection,Mapping,Zclipping,DepthCueing,AntiAliasing
        --           et Conversions) .
        --          Provides a set of services common to all types of view.
        --  Warning: The default parameters are defined by the class
        --          Viewer (Example : SetDefaultViewSize()).
        --          Certain methods are mouse oriented, and it is
        --          necessary to know the difference between the start and
        --          the continuation of this gesture in putting the method
        --          into operation.
        --          Example : Shifting the eye-view along the screen axes.
        --
        --              View->Move(10.,20.,0.,True)     (Starting motion)
        --              View->Move(15.,-5.,0.,False)    (Next motion)

uses

        -- S3892
        Pnt                     from gp,
        Dir                     from gp,
        Ax3                     from gp,
        LayerMgr                from V3d,
        ColorScale              from V3d,
        ColorScale              from Aspect,
        Array2OfReal            from TColStd,
        Grid                    from Aspect,
        Handle                  from Aspect,
        Structure               from Graphic3d,
        Group                   from Graphic3d,

        ListOfTransient                   from V3d,
        ListIteratorOfListOfTransient     from TColStd,
        TypeOfView                        from V3d,
        TypeOfAxe                         from V3d,
        TypeOfOrientation                 from V3d,
        TypeOfShadingModel                from V3d,
        TypeOfSurfaceDetail               from V3d,
        TextureEnv                        from Graphic3d,
        TypeOfVisualization               from V3d,
        TypeOfZclipping                   from V3d,
        TypeOfBackfacingModel             from V3d,
        StereoDumpOptions                 from V3d,
        Viewer                            from V3d,
        Light                             from V3d,
        View                              from Visual3d,
        ContextView                       from Visual3d,
        Vector                            from Graphic3d,
        Vertex                            from Graphic3d,
        Camera_Handle                     from Graphic3d,
        Window                            from Aspect,
        PixMap                            from Image,
        BufferType                        from Graphic3d,
        Background                        from Aspect,
        GradientBackground                from Aspect,
        TypeOfColor                       from Quantity,
        NameOfColor                       from Quantity,
        Color                             from Quantity,
        Length                            from Quantity,
        PlaneAngle                        from Quantity,
        Parameter                         from Quantity,
        Factor                            from Quantity,
        Ratio                             from Quantity,
        Coefficient                       from Quantity,
        Coordinate                        from V3d,
        Array2OfReal                      from TColStd,
        ViewerPointer                     from V3d,
        TypeOfTriedronEcho                from Aspect,
        TypeOfTriedronPosition            from Aspect,
        RenderingContext                  from Aspect,
        GraphicCallbackProc               from Aspect,
        FillMethod                        from Aspect,
        GradientFillMethod                from Aspect,
        FontAspect                        from Font,
        AsciiString                       from TCollection,
        ExtendedString                    from TCollection,
        PrintAlgo                         from Aspect,
        ClipPlane_Handle                  from Graphic3d,
        SequenceOfHClipPlane              from Graphic3d,
        RenderingMode                     from Graphic3d,
        RenderingParams                   from Graphic3d,
        XYZ                               from gp,
        Box                               from Bnd
raises

        BadValue from V3d, TypeMismatch from Standard,
        MultiplyDefined from Standard,UnMapped from V3d

is

        Create ( VM : Viewer; Type : TypeOfView from V3d = V3d_ORTHOGRAPHIC );
        ---Purpose: Initializes the view.

        Create (theVM : Viewer; theView : View from V3d);
        ---Purpose: Initializes the view by copying.

        --------------------------------------------------------
        ---Category: Methods to modify the Status of the view
        --------------------------------------------------------

        SetWindow ( me : mutable ; IdWin : Window )
        ---Purpose: Activates the view in the window specified and Map the
        --          Window to the screen.
        raises MultiplyDefined from Standard;
        ---Level: Public
        ---Purpose:  Warning! raises MultiplyDefined from Standard
        --      if the view is already activated in a window.
        --  Warning: The view is centered and resized to preserve
        --          the height/width ratio of the window.

        SetWindow ( me            : mutable ;
                    aWindow       : Window from Aspect;
                    aContext      : RenderingContext from Aspect;
                    aDisplayCB    : GraphicCallbackProc from Aspect;
                    aClientData   : Address from Standard
          )
        ---Purpose: Activates the view in the specified Window
        --      If <aContext> is not NULL the graphic context is used
        --          to draw something in this view.
        --      Otherwise an internal graphic context is created.
        --      If <aDisplayCB> is not NULL then a user display CB is
        --      call at the end of the OCC graphic traversal and just
        --      before the swap of buffers. The <aClientData> is pass
        --      to this call back.
        raises MultiplyDefined from Standard;
        ---Level: Public
        ---Purpose:  Warning! raises MultiplyDefined from Standard
        --      if the view is already activated in a window.
        --  Warning: The view is centered and resized to preserve
        --          the height/width ratio of the window.

        SetMagnify (me: mutable; IdWin            : Window;
                                 aPreviousView    : View from V3d;
                                 x1 , y1 , x2 , y2: Integer from Standard)
        is static;

        Remove ( me );
        ---Level: Public
        ---Purpose: Destroys the view.

        Update ( me ) is static;
        ---Level: Public
        ---Purpose: Deprecated, Redraw() should be used instead.

        Redraw ( me );
        ---Level: Public
        ---Purpose: Redisplays the view even if there has not
        --          been any modification.
        --          Must be called if the view is shown.
        --          (Ex: DeIconification ) .

        RedrawImmediate ( me );
        ---Level: Public
        ---Purpose: Updates layer of immediate presentations.

        Invalidate ( me );
        ---Level: Public
        ---Purpose: Invalidates view content but does not redraw it.

        Redraw ( me ;x,y,width,height: Integer from Standard);
        ---Level: Public
        ---Purpose: Redisplays the view area after esxposure.
    -- [x,y] define the min xy area position
    -- [width,height] the size of the area in pixel unit.

        MustBeResized ( me : mutable )
        ---Level: Public
        ---Purpose: Must be called when the window supporting the
        --          view changes size.
        raises UnMapped from V3d;
        ---Purpose:      if the view is not mapped on a window.
        --  Warning: The view is centered and resized to preserve
        --          the height/width ratio of the window.

        DoMapping ( me : mutable );
        ---Level: Advanced
        ---Purpose: Must be called when the window supporting the
        --          view is mapped or unmapped.

        IsEmpty ( me ) returns Boolean;
        ---Level: Public
        ---Purpose: Returns the status of the view regarding
        --          the displayed structures inside
        --          Returns True is The View is empty

        UpdateLights (me);
        ---Level: Public
        ---Purpose: Updates the lights of the view. The view is redrawn.

        AutoZFit (me : mutable);
        ---Level: Public
        ---Purpose: If automatic z-range fitting is turned on, adjusts Z-min and Z-max
        --          projection volume planes with call to ZFitAll.

        ZFitAll (me : mutable; theScaleFactor : Real from Standard = 1.0);
        ---Level: Public
        ---Purpose: Change Z-min and Z-max planes of projection volume to match the
        --          displayed objects. 

        --------------------------------------------------------
        ---Category: Methods to modify the Attributes of the view
        --------------------------------------------------------

        SetBackgroundColor ( me : mutable ;
                        Type : TypeOfColor; V1, V2, V3 : Parameter );
        ---Level: Public
        ---Purpose: Defines the background colour of the view
        --          by supplying :
        --          the colour definition type,
        --          and the three corresponding values.

        SetBackgroundColor ( me : mutable ; Color : Color from Quantity );
        ---Level: Public
        ---Purpose: Defines the background colour of the view
        --          by supplying :
        --          the colour object.

        SetBackgroundColor ( me : mutable ; Name : NameOfColor );
        ---Level: Public
        ---Purpose: Defines the background colour of the view
        --          by supplying :
        --          the colour name in the form Quantity_NOC_xxxx .

        SetBgGradientColors ( me : mutable ;
                              Color1 : Color from Quantity;
                              Color2 : Color from Quantity;
                              FillStyle : GradientFillMethod from Aspect = Aspect_GFM_HOR;
                              update    : Boolean from Standard = Standard_False );
        ---Level: Public
        ---Purpose: Defines the gradient background colours of the view
        --          by supplying :
        --          two colour objects,
        --          and fill method (horizontal by default)

        SetBgGradientColors ( me : mutable ;
                              Color1 : NameOfColor;
                              Color2 : NameOfColor;
                              FillStyle : GradientFillMethod from Aspect = Aspect_GFM_HOR;
                              update    : Boolean from Standard = Standard_False );
        ---Level: Public
        ---Purpose: Defines the gradient background colours of the view
        --          by supplying :
        --          two colour names in the form Quantity_NOC_xxxx,
        --          and fill method (horizontal by default)

        SetBgGradientStyle( me : mutable ;
                            AMethod : GradientFillMethod from Aspect = Aspect_GFM_HOR;
                            update  : Boolean from Standard = Standard_False);
        ---Level: Public
        ---Purpose: Defines the gradient background fill method of the view

        SetBackgroundImage( me : mutable; FileName  : CString from Standard;
              FillStyle : FillMethod from Aspect = Aspect_FM_CENTERED;
                  update    : Boolean from Standard = Standard_False );
        ---Level: Public
        ---Purpose: Defines the background texture of the view
        ---         by supplying :
        ---         texture image file name,
        ---         and fill method (centered by default)

        SetBgImageStyle( me : mutable; FillStyle : FillMethod from Aspect;
                                   update    : Boolean from Standard = Standard_False );
        ---Level: Public
        ---Purpose: Defines the textured background fill method of the view

        SetAxis ( me : mutable; X,Y,Z : Coordinate ;
                                Vx,Vy,Vz : Parameter )
        ---Level: Public
        ---Purpose: Definition of an axis from its origin and
        --          its orientation .
        --          This will be the current axis for rotations and movements.
        raises BadValue from V3d;
        ---Purpose:  Warning! raises BadValue from V3d if the vector normal is NULL. .

        SetShadingModel ( me : mutable; Model : TypeOfShadingModel );
        ---Level: Public
        ---Purpose: Defines the shading model for the
        --          visualisation ZBUFFER mode.
        --          Various models are available.

        SetSurfaceDetail(me  : mutable; SurfaceDetail : TypeOfSurfaceDetail);
        ---Level: Public
        ---Purpose: select the kind of rendering for texture mapping
        --          no texture mapping by default

        SetTextureEnv(me  : mutable; ATexture  :  TextureEnv  from  Graphic3d);
        ---Level: Public
        ---Purpose: set the environment texture to use
        --          no environment texture by default

        SetVisualization ( me : mutable;
                                Mode : TypeOfVisualization from V3d );
        ---Level: Public
        ---Purpose: Defines the visualisation mode in the view.

        SetAntialiasingOn ( me : mutable );
        ---Level: Public
        ---Purpose: Activates antialiasing in the view.

        SetAntialiasingOff ( me : mutable );
        ---Level: Public
        ---Purpose: Desactivates antialiasing in the view.

        SetZClippingDepth ( me : mutable; Depth : Length );
        ---Level: Public
        ---Purpose: Defines the depth of the medium clipping plane.

        SetZClippingWidth ( me : mutable; Width : Length )
        ---Level: Public
        ---Purpose: Defines the thicknes around the medium clippling plane.   .
                raises BadValue from V3d;
        --      If the thickness is <= 0

        SetZClippingType ( me : mutable; Type : TypeOfZclipping );
        ---Level: Public
        ---Purpose: Defines the type of ZClipping.

        SetZCueingDepth ( me : mutable; Depth : Length );
        ---Level: Public
        ---Purpose: Defines the depth of the medium plane.

        SetZCueingWidth ( me : mutable; Width : Length )
        ---Level: Public
        ---Purpose: Defines the thickness around the medium plane.
                raises BadValue from V3d;
        --      If thickness is <= 0

        SetZCueingOn ( me : mutable );
        ---Level: Public
        ---Purpose: Activates ZCueing in the view.

        SetZCueingOff ( me : mutable );
        ---Level: Public
        ---Purpose: Desactivates ZCueing in the view.

        SetLightOn( me : mutable ; MyLight : Light from V3d )
        ---Level: Public
        ---Purpose: Activates MyLight in the view.
                raises BadValue from V3d;
        --      If No More Light can be activated in MyView .

        SetLightOn( me : mutable )
        ---Level: Public
        ---Purpose: Activates all the lights defined in this view.
                raises BadValue from V3d;
        --      If No More Light can be activated in MyView .

        SetLightOff( me : mutable ; MyLight : Light  from V3d );
        ---Level: Public
        ---Purpose: Desactivate MyLight in this view.

        SetLightOff( me : mutable );
        ---Level: Public
        ---Purpose: Deactivate all the Lights defined in this view.

        IsActiveLight( me ; aLight: Light  from V3d )
        returns Boolean from Standard;
        ---Level: Public
        ---Purpose: Returns TRUE when the light is active in this view.

        SetImmediateUpdate(me: mutable; theImmediateUpdate: Boolean from Standard)
        returns Boolean from Standard;
    	  ---Purpose: sets the immediate update mode and returns the previous one.

        ---------------------------------------------------
        --           Triedron methods
        ---------------------------------------------------

        ZBufferTriedronSetup ( me      : mutable;
                           XColor  : NameOfColor from Quantity = Quantity_NOC_RED;
                           YColor  : NameOfColor from Quantity = Quantity_NOC_GREEN;
                           ZColor  : NameOfColor from Quantity = Quantity_NOC_BLUE1;
                   SizeRatio : Real from Standard = 0.8;
                   AxisDiametr : Real from Standard = 0.05;
                   NbFacettes  : Integer from Standard = 12)
         is static;
        ---Level: Advanced
        ---Purpose: Customization of the ZBUFFER Triedron.
        ---         XColor,YColor,ZColor - colors of axis
        ---         SizeRatio - ratio of decreasing of the trihedron size when its phisical
        ---                     position comes out of the view
        ---         AxisDiametr - diameter relatively to axis length
        ---         NbFacettes - number of facettes of cylinders and cones

        TriedronDisplay ( me            : mutable;
                          APosition     : TypeOfTriedronPosition from Aspect  = Aspect_TOTP_CENTER;
                          AColor        : NameOfColor from Quantity = Quantity_NOC_WHITE ;
                          AScale        : Real from Standard  =  0.02;
                          AMode         : TypeOfVisualization from V3d = V3d_WIREFRAME )
                is static;
        ---Level: Advanced
        ---Purpose: Display of the Triedron.
        ---         Initialize position, color and length of Triedron axes.
        ---         The scale is a percent of the window width.
        ---Category:

        TriedronErase ( me : mutable )
                is static;
        ---Level: Advanced
        ---Purpose: Erases the Triedron.
        ---Category:

        TriedronEcho ( me       : mutable;
                       AType    : TypeOfTriedronEcho from Aspect  = Aspect_TOTE_NONE )
                is static;
        ---Level: Advanced
        ---Purpose: Highlights the echo zone of the Triedron.
        ---Category:

        ---------------------------------
        ---Category: Graduated trihedron
        ---------------------------------

        GetGraduatedTrihedron(me;
                              -- Names of axes --
                              xname, yname, zname : out ExtendedString from TCollection;
                              -- Draw names --
                              xdrawname, ydrawname, zdrawname : out Boolean from Standard;
                              -- Draw values --
                              xdrawvalues, ydrawvalues, zdrawvalues : out Boolean from Standard;
                              -- Draw grid --
                              drawgrid : out Boolean from Standard;
                              -- Draw axes --
                              drawaxes : out Boolean from Standard;
                              -- Number of splits along axes --
                              nbx, nby, nbz : out Integer from Standard;
                              -- Offset for drawing values --
                              xoffset, yoffset, zoffset : out Integer from Standard;
                              -- Offset for drawing names of axes --
                              xaxisoffset, yaxisoffset, zaxisoffset : out Integer from Standard;
                              -- Draw tickmarks --
                              xdrawtickmarks, ydrawtickmarks, zdrawtickmarks : out Boolean from Standard;
                              -- Length of tickmarks --
                              xtickmarklength, ytickmarklength, ztickmarklength : out Integer from Standard;
                              -- Grid color --
                              gridcolor : out Color from Quantity;
                              -- Colors of axis names --
                              xnamecolor, ynamecolor, znamecolor : out Color from Quantity;
                              -- Colors of axis and values --
                              xcolor, ycolor, zcolor : out Color from Quantity;
                              -- Name of font for names of axes --
                              fontOfNames : out AsciiString from TCollection;
                              -- Style of names of axes --
                              styleOfNames : out FontAspect from Font;
                              -- Size of names of axes --
                              sizeOfNames : out Integer from Standard;
                              -- Name of font for values --
                              fontOfValues : out AsciiString from TCollection;
                              -- Style of values --
                              styleOfValues : out FontAspect from Font;
                              -- Size of values --
                              sizeOfValues : out Integer from Standard)
        ---Purpose: Returns data of a graduated trihedron.
        is static;

        GraduatedTrihedronDisplay(me : mutable;
                                  -- Names of axes --
                                  xname : ExtendedString from TCollection = "X";
                                  yname : ExtendedString from TCollection = "Y";
                                  zname : ExtendedString from TCollection = "Z";
                                  -- Draw names --
                                  xdrawname : Boolean from Standard = Standard_True;
                                  ydrawname : Boolean from Standard = Standard_True;
                                  zdrawname : Boolean from Standard = Standard_True;
                                  -- Draw values --
                                  xdrawvalues : Boolean from Standard = Standard_True;
                                  ydrawvalues : Boolean from Standard = Standard_True;
                                  zdrawvalues : Boolean from Standard = Standard_True;
                                  -- Draw grid --
                                  drawgrid : Boolean from Standard = Standard_True;
                                  -- Draw axes --
                                  drawaxes : Boolean from Standard = Standard_True;
                                  -- Number of splits along axes --
                                  nbx : Integer from Standard = 3;
                                  nby : Integer from Standard = 3;
                                  nbz : Integer from Standard = 3;
                                  -- Offset for drawing values --
                                  xoffset : Integer from Standard = 10;
                                  yoffset : Integer from Standard = 10;
                                  zoffset : Integer from Standard = 10;
                                  -- Offset for drawing names of axes --
                                  xaxisoffset : Integer from Standard = 30;
                                  yaxisoffset : Integer from Standard = 30;
                                  zaxisoffset : Integer from Standard = 30;
                                  -- Draw tickmarks --
                                  xdrawtickmarks : Boolean from Standard = Standard_True;
                                  ydrawtickmarks : Boolean from Standard = Standard_True;
                                  zdrawtickmarks : Boolean from Standard = Standard_True;
                                  -- Length of tickmarks --
                                  xtickmarklength : Integer from Standard = 10;
                                  ytickmarklength : Integer from Standard = 10;
                                  ztickmarklength : Integer from Standard = 10;
                                  -- Grid color --
                                  gridcolor : Color from Quantity = Quantity_NOC_WHITE;
                                  -- X name color --
                                  xnamecolor : Color from Quantity = Quantity_NOC_RED;
                                  -- Y name color --
                                  ynamecolor : Color from Quantity = Quantity_NOC_GREEN;
                                  -- Z name color --
                                  znamecolor : Color from Quantity = Quantity_NOC_BLUE1;
                                  -- X color of axis and values --
                                  xcolor : Color from Quantity = Quantity_NOC_RED;
                                  -- Y color of axis and values --
                                  ycolor : Color from Quantity = Quantity_NOC_GREEN;
                                  -- Z color of axis and values --
                                  zcolor : Color from Quantity = Quantity_NOC_BLUE1;
                                  -- Name of font for names of axes --
                                  fontOfNames : AsciiString from TCollection = "Arial";
                                  -- Style of names of axes --
                                  styleOfNames : FontAspect from Font = Font_FA_Bold;
                                  -- Size of names of axes --
                                  sizeOfNames : Integer from Standard = 12;
                                  -- Name of font for values --
                                  fontOfValues : AsciiString from TCollection = "Arial";
                                  -- Style of values --
                                  styleOfValues : FontAspect from Font = Font_FA_Regular;
                                  -- Size of values --
                                  sizeOfValues : Integer from Standard = 12)
        ---Purpose: Displays a graduated trihedron.
        is static;

        GraduatedTrihedronErase(me : mutable)
        ---Purpose: Erases a graduated trihedron from the view.
        is static;

        ---------------------------------------------------
        --           Color Scale methods
        ---------------------------------------------------

        SetLayerMgr(me : mutable; aMgr : LayerMgr from V3d);

        ColorScaleDisplay(me : mutable);

        ColorScaleErase(me : mutable);

        ColorScaleIsDisplayed(me)
        returns Boolean from Standard;

        ColorScale(me)
        returns ColorScale from Aspect;

        --------------------------------------------------------
        ---Category: Methods to modify the Projection of the view
        --------------------------------------------------------

        SetFront(me: mutable);
        ---Level: Public
        ---Purpose: modify the Projection of the view perpendicularly to
        --          the privileged plane of the viewer.

        Rotate ( me : mutable ; Ax,Ay,Az : PlaneAngle ;
                                Start    : Boolean = Standard_True )
        ---Level: Public
        ---Purpose: Rotates the eye about the coordinate system of
        --          reference of the screen
        --          for which the origin is the view point of the projection,
        --          with a relative angular value in RADIANS with respect to
        --          the initial position expressed by Start = Standard_True
        raises BadValue from V3d;
        ---Purpose:  Warning! raises BadValue from V3d
        --      If the eye, the view point, or the high point are
        --          aligned or confused.

        Rotate ( me : mutable ; Ax,Ay,Az : PlaneAngle ;
                                X,Y,Z    : Coordinate ;
                                Start    : Boolean = Standard_True )
        ---Level: Public
        ---Purpose: Rotates the eye about the coordinate system of
        --          reference of the screen
        --          for which the origin is Gravity point {X,Y,Z},
        --          with a relative angular value in RADIANS with respect to
        --          the initial position expressed by Start = Standard_True
                raises BadValue from V3d;
        ---Purpose:      If the eye, the view point, or the high point are
        --          aligned or confused.

        Rotate ( me : mutable ; Axe      : TypeOfAxe ; Angle : PlaneAngle ;
                                X,Y,Z    : Coordinate ;
                                Start    : Boolean = Standard_True );
        ---Level: Public
        ---Purpose: Rotates the eye about one of the coordinate axes of
        --          of the view for which the origin is the Gravity point{X,Y,Z}
        --          with an relative angular value in RADIANS with
        --          respect to the initial position expressed by
        --          Start = Standard_True

        Rotate ( me : mutable ; Axe    : TypeOfAxe ; Angle : PlaneAngle ;
                                Start : Boolean = Standard_True ) ;
        ---Level: Public
        ---Purpose: Rotates the eye about one of the coordinate axes of
        --          of the view for which the origin is the view point of the
        --          projection with an relative angular value in RADIANS with
        --          respect to the initial position expressed by
        --          Start = Standard_True

        Rotate ( me : mutable ; Angle : PlaneAngle ;
                                Start : Boolean = Standard_True );
        ---Level: Public
        ---Purpose: Rotates the eye around the current axis a relative
        --          angular value in RADIANS with respect to the initial
        --          position expressed by Start = Standard_True

        Move ( me : mutable ; Dx,Dy,Dz : Length ;
                              Start    : Boolean = Standard_True )
        ---Level: Public
        ---Purpose: Movement of the eye parallel to the coordinate system
        --          of reference of the screen a distance relative to the
        --          initial position expressed by Start = Standard_True.
                raises BadValue from V3d;
        --      If the eye, the view point, or the high point are
        --      aligned or confused.

        Move ( me : mutable ; Axe   : TypeOfAxe ; Length : Length ;
                              Start : Boolean = Standard_True )
        ---Level: Public
        ---Purpose: Movement of the eye parallel to one of the axes of the
        --          coordinate system of reference of the view a distance
        --          relative to the initial position expressed by
        --          Start = Standard_True.
                raises BadValue from V3d;
        --      If the eye, view point, or high point are aligned or confused.

        Move ( me : mutable ; Length : Length ;
                              Start  : Boolean = Standard_True )
        ---Level: Public
        ---Purpose: Movement of the eye parllel to the current axis
        --          a distance relative to the initial position
        --          expressed by Start = Standard_True
                raises BadValue from V3d;
        --      If the eye, view point, or high point are aligned or confused.

        Translate ( me : mutable ; Dx,Dy,Dz : Length ;
                                   Start    : Boolean = Standard_True )
        ---Level: Public
        ---Purpose: Movement of the ye and the view point parallel to the
        --          frame of reference of the screen a distance relative
        --          to the initial position expressed by
        --          Start = Standard_True
                raises BadValue from V3d;
        --      If the eye, view point, or high point are aligned or confused.

        Translate ( me : mutable ; Axe   : TypeOfAxe ; Length : Length ;
                                   Start : Boolean = Standard_True );
        ---Level: Public
        ---Purpose: Movement of the eye and the view point parallel to one
        --          of the axes of the fame of reference of the view a
        --          distance relative to the initial position
        --          expressed by Start = Standard_True

        Translate ( me : mutable ; Length : Length ;
                                   Start  : Boolean = Standard_True );
        ---Level: Public
        ---Purpose: Movement of the eye and view point parallel to
        --          the current axis a distance relative to the initial
        --          position expressed by Start = Standard_True

        Place (me            : mutable;
               theXp         : Integer from Standard;
               theYp         : Integer from Standard;
               theZoomFactor : Factor from Quantity = 1)
        ---Level: Public
        ---Purpose: places the point of the view corresponding
        --          at the pixel position x,y at the center of the window
        --          and updates the view.
        is static;

        Turn ( me : mutable ; Ax,Ay,Az : PlaneAngle ;
                              Start    : Boolean = Standard_True )
        ---Level: Public
        ---Purpose: Rotation of the view point around the frame of reference
        --          of the screen for which the origin is the eye of the
        --          projection with a relative angular value in RADIANS
        --          with respect to the initial position expressed by
        --          Start = Standard_True
                raises BadValue from V3d;
        --      If the eye, view point, or high point are aligned or confused.

        Turn ( me : mutable ; Axe : TypeOfAxe ; Angle : PlaneAngle ;
                              Start : Boolean = Standard_True )
       ;
        ---Level: Public
        ---Purpose: Rotation of the view point around one of the axes of the
        --          frame of reference of the view for which the origin is
        --          the eye of the projection with an angular value in
        --          RADIANS relative to the initial position expressed by
        --          Start = Standard_True

        Turn ( me : mutable ; Angle : PlaneAngle ;
                              Start : Boolean = Standard_True );
        ---Level: Public
        ---Purpose: Rotation of the view point around the current axis an
        --          angular value in RADIANS relative to the initial
        --          position expressed by Start = Standard_True

        SetTwist ( me : mutable ; Angle : PlaneAngle )
        ---Level: Public
        ---Purpose: Defines the angular position of the high point of
        --          the reference frame of the view with respect to the
        --          Y screen axis with an absolute angular value in
        --          RADIANS.
                raises BadValue from V3d;
        --      If the eye, view point, or high point are aligned or confused.

        SetEye( me : mutable ; X,Y,Z : Coordinate )
        ---Level: Public
        ---Purpose: Defines the position of the eye..
                raises BadValue from V3d ;
        --      If the eye, view point, or high point are aligned or confused.

        SetDepth( me : mutable ; Depth : Length )
        ---Level: Public
        ---Purpose: Defines the Depth of the eye from the view point
        --          without update the projection .
                raises BadValue from V3d ;
        --      If the Depth is <= 0.

        SetProj( me : mutable ; Vx,Vy,Vz : Parameter )
        ---Level: Public
        ---Purpose: Defines the orientation of the projection.
                raises BadValue from V3d ;
        --      If the eye, view point, or high point are aligned or confused.

        SetProj( me : mutable ; Orientation : TypeOfOrientation )
        ---Level: Public
        ---Purpose: Defines the orientation of the projection .
                raises BadValue from V3d ;
        --      If the eye, view point, or high point are aligned or confused.
        --          Updates the view

        SetAt( me : mutable ; X,Y,Z : Coordinate )
        ---Level: Public
        ---Purpose: Defines the position of the view point.
                raises BadValue from V3d ;
        --      If the eye, view point, or high point are aligned or confused.

        SetUp( me : mutable ; Vx,Vy,Vz : Parameter )
        ---Level: Public
        ---Purpose: Defines the orientation of the high point.
                raises BadValue from V3d ;
        --      If the eye, view point, or high point are aligned or confused.

        SetUp( me : mutable ; Orientation : TypeOfOrientation )
        ---Level: Public
        ---Purpose: Defines the orientation(SO) of the high point.
                raises BadValue from V3d ;
        --      If the eye, view point, or high point are aligned or confused.

        SetViewOrientationDefault( me : mutable );
        ---Level: Public
        ---Purpose: Saves the current state of the orientation of the view
        --          which will be the return state at ResetViewOrientation.

        ResetViewOrientation ( me : mutable );
        ---Level: Public
        ---Purpose: Resets the orientation of the view.
        --          Updates the view

        --------------------------------------------------------
        ---Category: Methods to modify the Mapping of the view
        --------------------------------------------------------

        Panning (me            : mutable;
                 theDXv        : Real from Standard;
                 theDYv        : Real from Standard;
                 theZoomFactor : Factor from Quantity = 1;
                 theToStart    : Boolean = Standard_True);
        ---Level: Public
        ---Purpose: Translates the center of the view along "x" and "y" axes of
        -- view projection. Can be used to perform interactive panning operation.
        -- In that case the DXv, DXy parameters specify panning relative to the
        -- point where the operation is started.
        -- @param theDXv [in] the relative panning on "x" axis of view projection, in view space coordinates.
        -- @param theDYv [in] the relative panning on "y" axis of view projection, in view space coordinates.
        -- @param theZoomFactor [in] the zooming factor.
        -- @param theToStart [in] pass TRUE when starting panning to remember view
        -- state prior to panning for relative arguments. If panning is started,
        -- passing {0, 0} for {theDXv, theDYv} will return view to initial state.
        -- Performs update of view.

        SetCenter (me : mutable; theXp, theYp : Integer from Standard)
        ---Level: Public
        ---Purpose: Relocates center of screen to the point, determined by
        -- {Xp, Yp} pixel coordinates relative to the bottom-left corner of
        -- screen. To calculate pixel coordinates for any point from world
        -- coordinate space, it can be projected using "Project".
        -- @param theXp [in] the x coordinate.
        -- @param theYp [in] the y coordinate.
        raises BadValue from V3d;
        -- If one of the dimensions of the projection is NULL.

        SetSize ( me : mutable; theSize : Length )
        ---Level: Public
        ---Purpose: Defines the view projection size in its maximum dimension,
        --          keeping the inital height/width ratio unchanged.
                raises BadValue from V3d;
        --      If <theSize> is <= 0.0

        SetZSize ( me : mutable ; Size : Length )
        ---Level: Public
        ---Purpose: Defines the Depth size of the view
        --          Front Plane will be set to Size/2.
        --          Back  Plane will be set to -Size/2.
        --          Any Object located Above the Front Plane or
        --                             behind the Back Plane will be Clipped .
        --          NOTE than the XY Size of the View is NOT modified .
                raises BadValue from V3d ;
        --      If the size of the view is <= 0

        SetZoom ( me : mutable ; Coef : Factor ; Start : Boolean = Standard_True )
        ---Level: Public
        ---Purpose: Zooms the view by a factor relative to the initial
        --          value expressed by Start = Standard_True
        --          Updates the view.
                raises BadValue from V3d ;
        --      If the zoom coefficient is <= 0

        SetScale ( me : mutable ; Coef : Factor )
        ---Level: Public
        ---Purpose: Zooms the view by a factor relative to the value
        --          initialised by SetViewMappingDefault().
        --          Updates the view.
                raises BadValue from V3d ;
        --      If the zoom coefficient is <= 0

    SetAxialScale ( me : mutable ; Sx, Sy, Sz : Real from Standard )
        ---Level: Public
        ---Purpose: Sets  anisotropic (axial)  scale  factors  <Sx>, <Sy>, <Sz>  for  view <me>.
    -- Anisotropic  scaling  operation  is  performed  through  multiplying
    -- the current view  orientation  matrix  by  a  scaling  matrix:
    -- || Sx  0   0   0 ||
    -- || 0   Sy  0   0 ||
    -- || 0   0   Sz  0 ||
    -- || 0   0   0   1 ||
        -- Updates the view.
                raises BadValue from V3d ;
        --      If the one of factors <= 0

        FitAll (me : mutable;
                theMargin : Coefficient = 0.01;
                theToUpdate : Boolean from Standard = Standard_True);
        ---Level: Public
        ---Purpose: Adjust view parameters to fit the displayed scene, respecting height / width ratio.
        --          The Z clipping range (depth range) is fitted if AutoZFit flag is TRUE.
        --          Throws program error exception if margin coefficient is < 0 or >= 1.
        --          Updates the view.
        --          @param theMargin [in] the margin coefficient for view borders.
        --          @param theToUpdate [in] flag to perform view update.

        DepthFitAll( me : mutable ;   Aspect : Coefficient = 0.01;
                                      Margin : Coefficient = 0.01 );
        ---Level: Public
        ---Purpose: Adjusts the viewing volume so as not to clip the displayed objects by front and back
        --          and back clipping planes. Also sets depth value automatically depending on the
        --          calculated Z size and Aspect parameter.
        --          NOTE than the original XY size of the view is NOT modified .

        FitAll (me : mutable;
                theMinXv : Real from Standard;
                theMinYv : Real from Standard;
                theMaxXv : Real from Standard;
                theMaxYv : Real from Standard)
        ---Level: Public
        ---Purpose: Centers the defined projection window so that it occupies
        --          the maximum space while respecting the initial
        --          height/width ratio.
        --          NOTE than the original Z size of the view is NOT modified .
                raises BadValue from V3d;
        --              If the defined projection window has zero size.

        WindowFit (me : mutable; theMinXp, theMinYp, theMaxXp, theMaxYp : Integer)
        ---Level: Public
        ---Purpose: Centers the defined PIXEL window so that it occupies
        -- the maximum space while respecting the initial height/width ratio.
        -- NOTE than the original Z size of the view is NOT modified.
        -- @param theMinXp [in] pixel coordinates of minimal corner on x screen axis.
        -- @param theMinYp [in] pixel coordinates of minimal corner on y screen axis.
        -- @param theMaxXp [in] pixel coordinates of maximal corner on x screen axis.
        -- @param theMaxYp [in] pixel coordinates of maximal corner on y screen axis.
        is static;
        SetViewMappingDefault( me : mutable );
        ---Level: Public
        ---Purpose: Saves the current view mapping. This will be the
        --          state returned from ResetViewmapping.

        ResetViewMapping ( me : mutable );
        ---Level: Public
        ---Purpose: Resets the centering of the view.
        --          Updates the view

        Reset ( me : mutable; update : Boolean from Standard = Standard_True );
        ---Level: Public
        ---Purpose: Resets the centering and the orientation of the view
        --          Updates the view
        ---------------------------------------------------
        ---Category: Inquire methods
        ---------------------------------------------------

        Convert( me ; Vp : Integer ) returns Length
        ---Level: Public
        ---Purpose : Converts the PIXEL value
        --           to a value in the projection plane.
        raises UnMapped from V3d;
        --      If the view is not mapped on the window.

        Convert( me ; Xp,Yp : Integer ; Xv,Yv : out Coordinate )
        ---Level: Public
        ---Purpose : Converts the point PIXEL into a point projected
        --           in the reference frame of the projection plane.
        raises UnMapped from V3d;
        --      If the view is not mapped on the window.

        Convert( me ; Vv : Length ) returns Integer
        ---Level: Public
        ---Purpose : Converts tha value of the projection plane into
        --           a PIXEL value.
        raises UnMapped from V3d;
        --      If the view is not mapped on the window.

        Convert( me ; Xv,Yv : Coordinate ; Xp,Yp : out Integer )
        ---Level: Public
        ---Purpose : Converts the point defined in the reference frame
        --           of the projection plane into a point PIXEL.
        raises UnMapped from V3d;
        --      If the view is not mapped on the window.

        Convert( me ; Xp,Yp : Integer ; X,Y,Z : out Coordinate)
        ---Level: Public
        ---Purpose : Converts the projected point into a point
        --           in the reference frame of the view corresponding
        --           to the intersection with the projection plane
        --           of the eye/view point vector.
        raises UnMapped from V3d;
        --      If the view is not mapped on the window.

        ConvertWithProj( me ; Xp,Yp : Integer ; X,Y,Z : out Coordinate ; Vx,Vy,Vz : out Parameter)
        ---Level: Public
        ---Purpose : Converts the projected point into a point
        --           in the reference frame of the view corresponding
        --           to the intersection with the projection plane
        --           of the eye/view point vector and returns the
        --           projection ray for further computations.
        raises UnMapped from V3d;
        --      If the view is not mapped on the window.

        ConvertToGrid( me ; Xp,Yp : Integer ; Xg,Yg,Zg : out Coordinate)
        ---Level: Public
        ---Purpose : Converts the projected point into the nearest grid point
        --           in the reference frame of the view corresponding
        --           to the intersection with the projection plane
        --           of the eye/view point vector and display the grid marker.
    --  Warning: When the grid is not active the result is identical to the above Convert() method.
    -- How to use:
    -- 1) Enable the grid echo display
    --    myViewer->SetGridEcho(Standard_True);
    -- 2) When application receive a move event:
    --   2.1) Check if any object is detected
    --     if( myInteractiveContext->MoveTo(x,y) == AIS_SOD_Nothing ) {
    --   2.2) Check if the grid is active
        --     if( myViewer->Grid()->IsActive() ) {
    --   2.3) Display the grid echo and gets the grid point
        --       myView->ConvertToGrid(x,y,X,Y,Z);
        --       myView->Viewer()->ShowGridEcho (myView, Graphic3d_Vertex (X,Y,Z));
        --       myView->RedrawImmediate();
    --   2.4) Else this is the standard case
        --     } else myView->Convert(x,y,X,Y,Z);
        raises UnMapped from V3d;
        --      If the view is not mapped on the window.

        ConvertToGrid( me ; X,Y,Z : Coordinate ; Xg,Yg,Zg : out Coordinate)
        ---Level: Public
        ---Purpose : Converts the point into the nearest grid point
        --           and display the grid marker.
    ---Warning: When the grid is not active the result is identical
    --     to the previous point.
        raises UnMapped from V3d;
        --      If the view is not mapped on the window.

        Convert( me ; X,Y,Z : Coordinate; Xp,Yp : out Integer) ;
        ---Level: Public
        ---Purpose : Projects the point defined in the reference frame of
        --           the view into the projected point in the associated window.

--        RefToPix( me ; X,Y,Z : Coordinate; Xp,Yp : out Integer) ;
--        ---Purpose : Projects the point defined in the reference frame of
--        --           the view into the projected point in the associated window.
--  Obsolete : Use Convert(X,Y,Z,Xp,Yp);

--        PixToRef( me ; Xp,Yp : Integer; X,Y,Z : out Coordinate) ;
--        ---Purpose : Converts the projected point in the associated window of
--        --           the view into the point defined in the reference frame.
--  Obsolete : Use Convert(Xp,Yp,X,Y,Z);

        Project( me ; X,Y,Z : Coordinate; Xp,Yp : out Coordinate) ;
        ---Level: Public
        ---Purpose : Converts the point defined in the user space of
        --           the view to the projected view plane point at z 0.

        BackgroundColor( me; Type : TypeOfColor ; V1, V2, V3 : out Parameter) ;
        ---Level: Public
        ---Purpose: Returns the Background color values of the view
        --          depending of the color Type.

        BackgroundColor( me ) returns Color from Quantity;
        ---Level: Public
        ---Purpose: Returns the Background color object of the view.

        GradientBackgroundColors( me;
                                  Color1 : out Color from Quantity;
                                  Color2 : out Color from Quantity) ;
        ---Level: Public
        ---Purpose: Returns the gradient background colour objects of the view.

	GradientBackground ( me ) returns GradientBackground from Aspect;
	---Level: Public
	---Purpose: Returns the gradient background of the view.

        Scale ( me ) returns Factor ;
        ---Level: Public
        ---Purpose: Returns the current value of the zoom expressed with
        --          respect to SetViewMappingDefault().

    AxialScale ( me ; Sx, Sy, Sz : out Real from Standard ) ;
        ---Level: Public
        ---Purpose: Returns the current values of the anisotropic (axial) scale factors.

        Size ( me; Width, Height : out Length );
        ---Level: Public
        ---Purpose: Returns the height and width of the view.

        ZSize ( me ) returns Real ;
        ---Level: Public
        ---Purpose: Returns the Depth of the view .

        Eye( me ; X,Y,Z : out Coordinate );
        ---Level: Public
        ---Purpose: Returns the position of the eye.

        FocalReferencePoint (me ; X,Y,Z : out Coordinate );
        ---Level: Public
        ---Purpose: Returns the position of point which emanating the
        --          projections.

        ProjReferenceAxe( me ; Xpix,Ypix           : Integer ;
                               XP,YP,ZP,VX,VY,VZ   : out Coordinate );
        ---Level: Public
        ---Purpose: Returns the coordinate of the point (Xpix,Ypix)
        --          in the view (XP,YP,ZP), and the projection vector of the
        --          view passing by the point (for PerspectiveView).

        Depth( me ) returns Length ;
        ---Level: Public
        ---Purpose: Returns the Distance between the Eye and View Point.

        Proj( me ; Vx,Vy,Vz : out Parameter );
        ---Level: Public
        ---Purpose: Returns the projection vector.

        At( me ; X,Y,Z : out Coordinate );
        ---Level: Public
        ---Purpose: Returns the position of the view point.

        Up( me ; Vx,Vy,Vz : out Parameter );
        ---Level: Public
        ---Purpose: Returns the vector giving the position of the high point.

        Twist( me ) returns PlaneAngle ;
        ---Level: Public
        ---Purpose: Returns in RADIANS the orientation of the view around
        --          the visual axis measured from the Y axis of the screen.

        ShadingModel ( me ) returns TypeOfShadingModel ;
        ---Level: Public
        ---Purpose: Returns the current shading model.

        SurfaceDetail(me) returns  TypeOfSurfaceDetail;
        ---Level: Public
        -- purpose: returns the current SurfaceDetail mode

        TextureEnv(me)  returns  TextureEnv  from  Graphic3d;
        ---Level: Public
        -- purpose: return the current environment texture used

        Visualization ( me ) returns TypeOfVisualization from V3d;
        ---Level: Public
        ---Purpose: Returns the current visualisation mode.

        Antialiasing ( me ) returns Boolean;
        ---Level: Public
        ---Purpose: Indicates if the antialiasing is active (True) or
        --          inactive (False).

        ZCueing ( me; Depth, Width : out Length ) returns Boolean ;
        ---Level: Public
        ---Purpose: Returns activity and information on the Zcueing.
        --          <Depth> : Depth of plane.
        --          <Width> : Thickness around the plane.

        ZClipping ( me; Depth, Width : out Length ) returns TypeOfZclipping;
        ---Level: Public
        ---Purpose: Returns current information on the ZClipping.
        --          <Depth> : Depth of plane.
        --          <Width> : Thickness around the plane.
        --          <TypeOfZclipping>  :        "BACK"
        --                                      "FRONT"
        --                                      "SLICE"
        --                                      "OFF"

        IfMoreLights( me ) returns Boolean;
        ---Level: Advanced
        ---Purpose: Returns True if One light more can be
        --          activated in this View.

        InitActiveLights(me: mutable);
        ---Level: Advanced
        ---Purpose: initializes an iteration on the active Lights.

        MoreActiveLights (me) returns Boolean from Standard;
        ---Level: Advanced
        ---Purpose: returns true if there are more active Light(s) to return.

        NextActiveLights (me: mutable);
        ---Level: Advanced
        ---Purpose : Go to the next active Light
        --           (if there is not, ActiveLight will raise an exception)

        ActiveLight(me) returns Light from V3d;
        ---Level: Advanced

        Viewer ( me ) returns Viewer from V3d;
        ---Level: Advanced
        ---Purpose: Returns the viewer in which the view has been created.

        IfWindow ( me ) returns Boolean;
        ---Level: Public
        ---Purpose: Returns True if MyView is associated with a window .

        Window ( me ) returns Window from Aspect
        ---Level: Public
        ---Purpose: Returns the Aspect Window associated with the view.
                raises BadValue from V3d;
        --      If MyView is not associated with a window

        Type( me ) returns TypeOfView from V3d;
        ---Level: Public
        ---Purpose: Returns the Type of the View

        Pan (me            : mutable;
             theDXp        : Integer from Standard;
             theDYp        : Integer from Standard;
             theZoomFactor : Factor from Quantity = 1;
             theToStart    : Boolean = Standard_True);
        ---Level: Public
        ---Purpose: Translates the center of the view along "x" and "y" axes of
        -- view projection. Can be used to perform interactive panning operation.
        -- In that case the DXp, DXp parameters specify panning relative to the
        -- point where the operation is started.
        -- @param theDXp [in] the relative panning on "x" axis of view projection, in pixels.
        -- @param theDYp [in] the relative panning on "y" axis of view projection, in pixels.
        -- @param theZoomFactor [in] the zooming factor.
        -- @param theToStart [in] pass TRUE when starting panning to remember view
        -- state prior to panning for relative arguments. Passing 0 for relative
        -- panning parameter should return view panning to initial state.
        -- Performs update of view.

        Zoom (me     : mutable;
              theXp1 : Integer from Standard;
              theYp1 : Integer from Standard;
              theXp2 : Integer from Standard;
              theYp2 : Integer from Standard)
        is static;
        ---Level: Public
        ---Purpose: Zoom the view according to a zoom factor computed
        -- from the distance between the 2 mouse position.
        -- @param theXp1 [in] the x coordinate of first mouse position, in pixels.
        -- @param theYp1 [in] the y coordinate of first mouse position, in pixels.
        -- @param theXp2 [in] the x coordinate of second mouse position, in pixels.
        -- @param theYp2 [in] the y coordinate of second mouse position, in pixels.

        StartZoomAtPoint (me    : mutable;
                          theXp : Integer from Standard;
                          theYp : Integer from Standard);
        ---Level: Public
        ---Purpose: Defines starting point for ZoomAtPoint view operation.
        -- @param theXp [in] the x mouse coordinate, in pixels.
        -- @param theYp [in] the y mouse coordinate, in pixels.

        ZoomAtPoint(me : mutable;
                    theMouseStartX : Integer from Standard;
                    theMouseStartY : Integer from Standard;
                    theMouseEndX   : Integer from Standard;
                    theMouseEndY   : Integer from Standard);
        ---Level: Public
        ---Purpose: Zooms the model at a pixel defined by the method StartZoomAtPoint().

        AxialScale  ( me: mutable; Dx, Dy: Integer from Standard;  Axis:  TypeOfAxe  from  V3d );
        ---Level: Public
        ---Purpose: Performs  anisotropic scaling  of  <me>  view  along  the  given  <Axis>.
            -- The  scale  factor  is  calculated on a basis of
            -- the mouse pointer displacement <Dx,Dy>.
        -- The  calculated  scale  factor  is  then  passed  to  SetAxialScale(Sx,  Sy,  Sz)  method.

        StartRotation(me : mutable ; X,Y :Integer from Standard;
               zRotationThreshold: Ratio from Quantity = 0.0);
        ---Level: Public
    ---Purpose: Begin the rotation of the view around the screen axis
    -- according to the mouse position <X,Y>.
    --  Warning: Enable rotation around the Z screen axis when <zRotationThreshold>
    -- factor is > 0 soon the distance from the start point and the center
    -- of the view is > (medium viewSize * <zRotationThreshold> ).
    -- Generally a value of 0.4 is usable to rotate around XY screen axis
    -- inside the circular threshold area and to rotate around Z screen axis
    -- outside this area.

        Rotation(me:mutable;  X,Y :Integer from Standard);
        ---Level: Public
    ---Purpose: Continues the rotation of the view
    -- with an angle computed from the last and new mouse position <X,Y>.

        FitAll ( me : mutable ; aWindow: Window from Aspect;
                      Umin, Vmin, Umax, Vmax : Coordinate )
        is static private;
        ---Level: Public
    ---Purpose: Change the scale factor and position of the view
    -- such as the bounding box <Umin, Vmin, Umax, Vmax> is contains
    -- in the view.


        -----------------------------------------
        ---Category: Private or Protected methods
        -----------------------------------------

        SetFocale( me : mutable ; Focale : Length )
        ---Purpose: Change View Plane Distance for Perspective Views
        raises TypeMismatch from Standard
        ---Purpose:  Warning! raises TypeMismatch from Standard if the view
        --          is not a perspective view.
        is static ;

        Focale( me ) returns Length;
        ---Purpose: Returns the View Plane Distance for Perspective Views

        View ( me) returns View from Visual3d is static ;
        ---Level: Advanced
        ---Purpose: Returns the associated Visual3d view.

        ScreenAxis( myclass ; Vpn,Vup        : Dir from gp ;
                              Xaxe,Yaxe,Zaxe : out Vector from Graphic3d )
                                        returns Boolean is private ;
        ---Purpose: Determines the screen axes in the reference
        --          framework of the view.


        TrsPoint( myclass ; V : Vertex from Graphic3d ;
                                Matrix : Array2OfReal from TColStd )
                                returns Vertex from Graphic3d is private ;
        ---Purpose: Transforms the Vertex V according to the matrice Matrix .
        
        ImmediateUpdate (me) is static protected;
    	  ---Purpose: 

        SetComputedMode ( me : mutable; aMode : Boolean from Standard )
        is static;
        ---Level: Advanced
        ---Purpose: Switches computed HLR mode in the view
        ---Category: Methods to modify the class definition

        ComputedMode ( me )
        returns Boolean from Standard
        is static;
        ---Level: Advanced
        ---Purpose: Returns the computed HLR mode state
        ---Category: Inquire methods

        MinMax ( me; Umin,Vmin, Umax,Vmax : out Coordinate ) returns Integer
        ---Purpose: Returns the objects number and the projection window
        --          of the objects contained in the view.
        is static private;

        MinMax ( me; Xmin,Ymin,Zmin, Xmax,Ymax,Zmax : out Coordinate )
        returns Integer
        ---Purpose: Returns the objects number and the box encompassing
        --          the objects contained in the view
        is static private;

        Gravity ( me; X,Y,Z : out Coordinate ) returns Integer
        ---Purpose: Returns the Objects number and the gravity center
        --          of ALL viewable points in the view
        is static private;

        Init(me: mutable) is private;

        ---Category: for compatibility.

        WindowFitAll ( me : mutable ; Xmin, Ymin, Xmax, Ymax : Integer);
        ---Purpose: idem than WindowFit

        Compute ( me; AVertex   : Vertex from Graphic3d )
                returns Vertex from Graphic3d
                is static private;
        ---Level: Internal
        ---Purpose: Returns a new vertex when the grid is activated.

        SetGrid ( me    : mutable;
                  aPlane: Ax3 from gp;
                  aGrid : Grid from Aspect )
                is static;
        ---Level: Internal
        ---Purpose: Defines or Updates the definition of the
        --          grid in <me>
        ---Category: Methods to modify the class definition

        SetGridGraphicValues ( me       : mutable;
                               aGrid    : Grid from Aspect )
                is static;
        ---Level: Internal
        ---Purpose: Defines or Updates the graphic definition of the
        --          grid in <me>
        ---Category: Methods to modify the class definition

        SetGridActivity ( me    : mutable;
                          aFlag : Boolean from Standard )
                is static;
        ---Level: Internal
        ---Purpose: Defines or Updates the activity of the
        --          grid in <me>
        ---Category: Methods to modify the class definition

        Dump ( me: mutable;
               theFile       : CString from Standard;
               theBufferType : BufferType from Graphic3d = Graphic3d_BT_RGB )
    returns Boolean from Standard;
        ---Level: Public
        ---Purpose: dump the full contents of the view at the same
        --          scale in the file <theFile>. The file name
        --          extension must be one of ".png",".bmp",".jpg",".gif".
        --          Returns FALSE when the dump has failed

      Print (me; hPrnDC: Handle from Aspect = 0;
             showDialog: Boolean = Standard_True;
             showBackground : Boolean = Standard_True;
             filename: CString = NULL;
             printAlgorithm : PrintAlgo from Aspect = Aspect_PA_STRETCH)
      returns Boolean from Standard is static;

        ---Level: Public
        ---Purpose: print the contents of the view to printer with preview.
    -- <hPrnDC> : If you have already an PrinterDeviceContext (HDC),
    -- then you can pass it to the print routines.
        -- If you don't have an PrinterDeviceContext, then this parameter should
    -- be NULL.
    -- <showDialog> : If hPrnDC == NULL, then you can force the print routines to
    -- open a Print Dialog box.
        -- If you want to do this, then set showDialog to TRUE
        -- If you don't want to see a dialog (only possible, if you have a hPrnDC
    -- or the dialog box was opened once before) then set <showDialog> to FALSE.
    -- <showBackground> : When set to FALSE then print the view without background color
    -- (background is white)
        -- else set to TRUE for printing with current background color.
    -- <filename>: If != NULL, then the view will be printed to a file.
    -- <printAlgorithm>: If you want to select the print algorithm, then you can
        -- specify one of existing algorithms: Aspect_PA_STRETCH, Aspect_PA_TILE.
    -- Returns Standard_True if the data is passed to the printer, otherwise
    -- Standard_False if the print operation failed. This might be related to
    -- insufficient memory or some internal errors. All this errors are
    -- indicated by the message boxes (on level of OpenGl_GraphicDriver).
    --  Warning: This function can reuse FBO assigned to the 
    --  view on level of OpenGl_GraphicDriver; Please take it into account if
    --  you use it for your purposes;
    --  Warning: Works only under Windows.

        ToPixMap (me : mutable;
                  theImage  : in out PixMap from Image;
                  theWidth  : Integer from Standard;
                  theHeight : Integer from Standard;
                  theBufferType : BufferType from Graphic3d = Graphic3d_BT_RGB;
                  theToKeepAspect : Boolean from Standard = Standard_True;
                  theStereoOptions : StereoDumpOptions from V3d = V3d_SDO_MONO)
        returns Boolean from Standard;
        ---Level   : Public
        ---Purpose : Dumps the full contents of the view
        --           to a pixmap of pixel size <theWidth> * <theHeight> and
        --           buffer type <theBufferType>. If <theToKeepAspect> is true
        --           the aspect ratio of view will be kept if <theWidth> and <theHeight>
        --           define another ratio.
        --           Pixmap will be automatically (re)allocated when needed.
        --           When dumping stereographic camera - the corresponding
        --           middle-point monographic projection will be used for dumping by default.
        --           <theStereoOptions> flags are to be used for dumping then left or
        --           right eye projections.

        SetBackFacingModel ( me     : mutable;
            aModel : TypeOfBackfacingModel from V3d = V3d_TOBM_AUTOMATIC)
            is static;
         ---Level   : Public
         ---Purpose : Manages display of the back faces
     -- When <aModel> is TOBM_AUTOMATIC the object backfaces
     -- are displayed only for surface objects and
     -- never displayed for solid objects.
     -- this was the previous mode.
     --      <aModel> is TOBM_ALWAYS_DISPLAYED the object backfaces
     --       are always displayed both for surfaces or solids.
     --      <aModel> is TOBM_NEVER_DISPLAYED the object backfaces
     --       are never displayed.

        BackFacingModel ( me )
            returns TypeOfBackfacingModel from V3d
        is static;
         ---Level   : Public
         ---Purpose : Returns current state of the back faces display

        EnableDepthTest( me; enable : Boolean from Standard = Standard_True )
        is static;
     ---Level: Public
     ---Purpose: turns on/off opengl depth testing

        IsDepthTestEnabled( me ) returns Boolean from Standard
        is static;
     ---Level: Public
     ---Purpose: returns the current state of the depth testing

        EnableGLLight( me; enable : Boolean from Standard = Standard_True )
        is static;
     ---Level: Public
     ---Purpose: turns on/off opengl lighting, currently used in triedron displaying

        IsGLLightEnabled( me ) returns Boolean from Standard
        is static;
     ---Level: Public
     ---Purpose: returns the current state of the gl lighting
     --          currently used in triedron displaying

     AddClipPlane (me : mutable; thePlane : ClipPlane_Handle from Graphic3d) is virtual;
     ---Purpose: Adds clip plane to the view. The composition of clip planes truncates the
     -- rendering space to convex volume. Number of supported clip planes can be consulted
     -- by PlaneLimit method of associated Visual3d_View. Please be aware that the planes
     -- which exceed the limit are ignored during rendering. 
     -- @param thePlane [in] the clip plane to be added to view.

     RemoveClipPlane (me : mutable; thePlane : ClipPlane_Handle from Graphic3d) is virtual;
     ---Purpose: Removes clip plane from the view.
     -- @param thePlane [in] the clip plane to be removed from view.

     SetClipPlanes (me : mutable; thePlanes : SequenceOfHClipPlane from Graphic3d);
     ---Purpose: Sets sequence of clip planes to the view. The planes that have been set
     -- before are removed from the view. The composition of clip planes
     -- truncates the rendering space to convex volume. Number of supported
     -- clip planes can be consulted by PlaneLimit method of associated
     -- Visual3d_View. Please be aware that the planes which exceed the limit
     -- are ignored during rendering. 
     -- @param thePlanes [in] the clip planes to set.

     GetClipPlanes (me) returns SequenceOfHClipPlane from Graphic3d;
     ---C++: return const&
     ---Purpose: Get clip planes.
     -- @return sequence clip planes that have been set for the view

    SetCamera (me : mutable; theCamera : Camera_Handle from Graphic3d) is static;
    ---Level: Public
    ---Purpose: Change camera used by view.

    Camera (me) returns Camera_Handle from Graphic3d is static;
    ---Level: Public
    ---C++: return const&
    ---Purpose: Returns camera object of the view.
    -- @return: handle to camera object, or NULL if 3D view does not use
    -- the camera approach.

    FitMinMax (me;
               theCamera          : Camera_Handle from Graphic3d;
               theBox             : Box from Bnd;
               theMargin          : Real from Standard;
               theResolution      : Real from Standard = 0.0;
               theToEnlargeIfLine : Boolean from Standard = Standard_True)
               returns Boolean from Standard is protected;
    ---Level: Protected
    ---Purpose: Transform camera eye, center and scale to fit in the
    -- passed bounding box specified in WCS.
    -- @param theCamera [in] the camera.
    -- @param theBox [in] the bounding box.
    -- @param theMargin [in] the margin coefficient for view borders.
    -- @param theResolution [in] the minimum size of projection of
    --        bounding box in Xv or Yv direction when it considered to
    --        be a thin plane or point (without a volume).
    --        In this case only the center of camera is adjusted.
    -- @param theToEnlargeIfLine [in] if passed TRUE - in cases when the
    -- whole bounding box projected into thin line going along
    -- Z-axis of screen, the view plane is enlarged such that
    -- we see the whole line on rotation, otherwise only the
    -- center of camera is adjusted.
    -- @return TRUE if the fit all operation can be done.

    Scale (me;
           theCamera : Camera_Handle from Graphic3d;
           theSizeXv : Real from Standard;
           theSizeYv : Real from Standard) is protected;
    ---Level: Protected
    ---Purpose: Scales camera to fit the view frame of defined width and height
    -- keeping the aspect. For orthogonal camera the method changes scale,
    -- for perspective adjusts Eye location about the Center point.
    -- @param theSizeXv [in] size of viewport frame on "x" axis.
    -- @param theSizeYv [in] size of viewport frame on "y" axis.

    Translate (me;
         theCamera : Camera_Handle from Graphic3d;
         theDXv    : Real from Standard;
         theDYv    : Real from Standard) is protected;
    ---Level: Protected
    -- Purpose: Translates camera eye and center along the view plane.
    -- @param theCamera [in] the camera to translate.
    -- @param theDXv [in] the translation in "x" direction.
    -- @param theDYv [in] the translation in "y" direction.

    RenderingParams (me) returns RenderingParams from Graphic3d is static;
    ---C++: return const &
    ---Level: Public
    ---Purpose: Returns current rendering parameters and effect settings.
    
    ChangeRenderingParams (me : mutable) returns RenderingParams from Graphic3d is static;
    ---C++: return &
    ---Level: Public
    ---Purpose: Returns reference to current rendering parameters and effect settings.

        IsCullingEnabled (me) returns Boolean from Standard is static;
     ---Level: Public
     ---Purpose: @return flag value of objects culling mechanism

        SetFrustumCulling (me : mutable; theMode : Boolean from Standard) is static;
     ---Level: Public
     ---Purpose: Turn on/off automatic culling of objects outside frustrum (ON by default)

fields

        myOldMouseX : Real is protected;
        myOldMouseY : Real is protected;
        myCamStartOpUp : Dir from gp is protected;
        myCamStartOpEye : Pnt from gp is protected;
        myCamStartOpBnd : Real[6] is protected;
        myCamStartOpCenter : Pnt from gp is protected;
        myCamera : Camera_Handle from Graphic3d is protected;

        MyViewer :              ViewerPointer from V3d ;
        MyActiveLights:         ListOfTransient from V3d;

        MyView :                View from Visual3d is protected ;
        MyViewContext :         ContextView from Visual3d ;
        MyBackground:           Background from Aspect ;
        MyGradientBackground:   GradientBackground from Aspect ;
        MyDefaultViewAxis:      Vector from Graphic3d ;
        MyDefaultViewPoint:     Vertex from Graphic3d ;

        MyWindow:               Window from Aspect;

        myActiveLightsIterator: ListIteratorOfListOfTransient from TColStd;

        sx,sy: Integer from Standard;
        rx,ry: Real from Standard;
        gx,gy,gz: Real from Standard;
        myComputedMode: Boolean from Standard;
        SwitchSetFront: Boolean from Standard;
        MyZoomAtPointX, MyZoomAtPointY : Integer from Standard;

        -- the 3d grid
        MyGrid                  :       Grid from Aspect;
        MyPlane                 :       Ax3 from gp;

        --MyColorScale            :       ColorScale from V3d;
        MyLayerMgr              :       LayerMgr from V3d;

        -- the transformation between XoY and the grid plane
        MyTrsf                  :       Array2OfReal from TColStd;

        -- echo
        MyGridEchoStructure             :       Structure from Graphic3d;
        MyGridEchoGroup                 :       Group from Graphic3d;

        myImmediateUpdate: Boolean from Standard is protected;

        myXscreenAxis           : Vector from Graphic3d;
        myYscreenAxis           : Vector from Graphic3d;
        myZscreenAxis           : Vector from Graphic3d;
        myViewAxis              : Vector from Graphic3d;
        myGravityReferencePoint : Vertex from Graphic3d;
        myCamProjectionShift    : Pnt from gp;

friends

        SetViewOn from class Viewer from V3d ( me : mutable ),
        SetViewOn from class Viewer from V3d ( me : mutable ; View : View from V3d ),
        SetViewOff from class Viewer from V3d ( me : mutable ),
        SetViewOff from class Viewer from V3d ( me : mutable ; View : View from V3d )

end View;
