-- Created on: 1997-05-09
-- Created by: Christian CAILLET
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ESDescr  from StepData    inherits EDescr

    ---Purpose : This class is intended to describe the authorized form for a
    --           Simple (not Plex) Entity, as a list of fields

uses CString, AsciiString from TCollection,
     HArray1OfTransient from TColStd, DictionaryOfInteger from Dico,
     PDescr from StepData, Described from StepData

is

    Create (name : CString) returns ESDescr;
    ---Purpose : Creates an ESDescr with a type name

    SetNbFields (me : mutable; nb : Integer);
    ---Purpose : Sets a new count of fields
    --           Each one is described by a PDescr

    SetField (me : mutable; num : Integer; name : CString; descr : PDescr);
    ---Purpose : Sets a PDescr to describe a field
    --           A Field is designated by its rank and name

    SetBase  (me : mutable; base : ESDescr);
    ---Purpose : Sets an ESDescr as based on another one
    --           Hence, if there are inherited fields, the derived ESDescr
    --           cumulates all them, while the base just records its own ones

    SetSuper (me : mutable; super : ESDescr);
    ---Purpose : Sets an ESDescr as "super-type". Applies an a base (non
    --           derived) ESDescr

    TypeName (me) returns CString;
    ---Purpose : Returns the type name given at creation time

    StepType (me) returns AsciiString from TCollection;
    ---Purpose : Returns the type name as an AsciiString
    ---C++ : return const &

    Base (me) returns ESDescr;
    ---Purpose : Returns the basic ESDescr, null if <me> is not derived

    Super (me) returns ESDescr;
    ---Purpose : Returns the super-type ESDescr, null if <me> is root

    IsSub (me; other : ESDescr) returns Boolean;
    ---Purpose : Tells if <me> is sub-type of (or equal to) another one

    NbFields (me) returns Integer;
    ---Purpose : Returns the count of fields

    Rank  (me; name : CString) returns Integer;
    ---Purpose : Returns the rank of a field from its name. 0 if unknown

    Name  (me; num  : Integer) returns CString;
    ---Purpose : Returns the name of a field from its rank. empty if outofrange

    Field (me; num : Integer) returns PDescr;
    ---Purpose : Returns the PDescr for the field <num> (or Null)

    NamedField (me; name : CString) returns PDescr;
    ---Purpose : Returns the PDescr for the field named <name> (or Null)

    	--  inherited

    Matches    (me; steptype : CString) returns Boolean;
    ---Purpose : Tells if a ESDescr matches a step type : exact or super type

    IsComplex  (me) returns Boolean;
    ---Purpose : Returns False

    NewEntity  (me) returns Described;
    ---Purpose : Creates a described entity (i.e. a simple one)

fields

    thenom   : AsciiString;
    thedescr : HArray1OfTransient;
    thenames : DictionaryOfInteger;
    thebase  : ESDescr;
    thesuper : ESDescr;

end ESDescr;
