-- Created by: Peter KURNEV
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Set from BOPTools 

	---Purpose: 

uses  
    ShapeEnum from TopAbs,
    Shape from TopoDS,
    ListOfShape from BOPCol,
    BaseAllocator from BOPCol 
    
--raises

is 
    Create 
    	returns Set from BOPTools;  
    ---C++: alias "virtual ~BOPTools_Set();"  
    ---C++: inline 
    
    Create (theAllocator: BaseAllocator from BOPCol)
    	returns Set from BOPTools; 
    ---C++: inline
     
    Assign(me:out;  
    	    Other : Set from BOPTools) 
    	returns Set from BOPTools; 
    ---C++: alias operator =
    ---C++: return &   
    ---C++: inline 
    
    Clear(me:out) 
    	is protected; 
    ---C++: inline
     
    Shape(me) 
    	 returns Shape from TopoDS; 
    ---C++: return const & 
    ---C++: inline 
     
    Add(me:out; 
    	    theS:Shape from TopoDS; 
    	    theType: ShapeEnum from TopAbs);  
    ---C++: inline 
     
    AddEdges(me:out; 
    	    theS:Shape from TopoDS);  
    ---C++: inline 
     
    NbShapes(me) 
    	    returns Integer from Standard; 
    ---C++: inline 
     
    IsEqual(me; 
    	    aOther:Set from BOPTools) 
	returns Boolean from Standard;   
    ---C++: inline 
     
    HashCode(me; 
	    Upper : Integer  from Standard)  
    	returns Integer from Standard;   	 
    ---C++: inline 
    
fields   
    myAllocator : BaseAllocator from BOPCol is protected; 
    myShapes    : ListOfShape from BOPCol is protected;   
    myShape     : Shape from TopoDS is protected; 
    myNbShapes  : Integer from Standard is protected;
    mySum       : Integer from Standard is protected; 
    myUpper     : Integer from Standard is protected; 
    
end Set;
