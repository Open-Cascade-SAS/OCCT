-- Created on: 2003-01-28
-- Created by: data exchange team
-- Copyright (c) 2003-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class ProductOrFormationOrDefinition from StepBasic
inherits SelectType from StepData

    ---Purpose: Representation of STEP SELECT type ProductOrFormationOrDefinition

uses
    Product from StepBasic,
    ProductDefinitionFormation from StepBasic,
    ProductDefinition from StepBasic

is
    Create returns ProductOrFormationOrDefinition from StepBasic;
	---Purpose: Empty constructor

    CaseNum (me; ent: Transient) returns Integer;
	---Purpose: Recognizes a kind of ProductOrFormationOrDefinition select type
	--          1 -> Product from StepBasic
	--          2 -> ProductDefinitionFormation from StepBasic
	--          3 -> ProductDefinition from StepBasic
	--          0 else

    Product (me) returns Product from StepBasic;
	---Purpose: Returns Value as Product (or Null if another type)

    ProductDefinitionFormation (me) returns ProductDefinitionFormation from StepBasic;
	---Purpose: Returns Value as ProductDefinitionFormation (or Null if another type)

    ProductDefinition (me) returns ProductDefinition from StepBasic;
	---Purpose: Returns Value as ProductDefinition (or Null if another type)

end ProductOrFormationOrDefinition;
