-- Created on: 1997-07-28
-- Created by: Pierre CHALAMET
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Texture2Dplane from Graphic3d

inherits Texture2D from Graphic3d

  ---Purpose: This class allows the management of a 2D texture defined from a plane equation
  -- Use the SetXXX() methods for positioning the texture as you want.

uses

  NameOfTexture2D    from Graphic3d,
  NameOfTexturePlane from Graphic3d,
  AsciiString        from TCollection,
  PixMap_Handle      from Image

is

  Create (theFileName : AsciiString from TCollection) returns mutable Texture2Dplane from Graphic3d;
  ---Purpose: Creates a texture from a file

  Create (theNOT : NameOfTexture2D from Graphic3d) returns mutable Texture2Dplane from Graphic3d;
  ---Purpose: Creates a texture from a predefined texture name set.

  Create (thePixMap : PixMap_Handle from Image) returns mutable Texture2Dplane from Graphic3d;
  ---Purpose: Creates a texture from the pixmap.

  SetPlaneS (me : mutable; A, B, C, D : ShortReal from Standard);
  ---Purpose:  Defines the texture projection plane for texture coordinate S
  -- default is <1.0, 0.0, 0.0, 0.0>

  SetPlaneT (me : mutable; A, B, C, D : ShortReal from Standard);
  ---Purpose: Defines the texture projection plane for texture coordinate T
  -- default is <0.0, 1.0, 0.0, 0.0>

  SetPlane (me : mutable; thePlane : NameOfTexturePlane from Graphic3d);
  ---Purpose:  Defines the texture projection plane for both S and T texture coordinate
  -- default is NOTP_XY meaning:
  --      <1.0, 0.0, 0.0, 0.0> for S
  -- and  <0.0, 1.0, 0.0, 0.0> for T

  SetScaleS (me : mutable; theVal : ShortReal from Standard);
  ---Purpose: Defines the texture scale for the S texture coordinate
  -- much easier than recomputing the S plane equation
  -- but the result is the same
  -- default to 1.0

  SetScaleT (me : mutable; theVal : ShortReal from Standard);
  ---Purpose: Defines the texture scale for the T texture coordinate
  -- much easier than recompution the T plane equation
  -- but the result is the same
  -- default to 1.0

  SetTranslateS (me : mutable; theVal : ShortReal from Standard);
  ---Purpose: Defines the texture translation for the S texture coordinate
  -- you can obtain the same effect by modifying the S plane
  -- equation but its not easier.
  -- default to 0.0

  SetTranslateT (me : mutable; theVal : ShortReal from Standard);
  ---Purpose:  Defines the texture translation for the T texture coordinate
  -- you can obtain the same effect by modifying the T plane
  -- equation but its not easier.
  -- default to 0.0

  SetRotation (me : mutable; theVal : ShortReal from Standard);
  ---Purpose: Sets the rotation angle of the whole texture.
  -- the same result might be achieved by recomputing the
  -- S and T plane equation but it's not the easiest way...
  -- the angle is expressed in degrees
  -- default is 0.0

  --
  -- inquire methods
  --

  Plane (me) returns NameOfTexturePlane from Graphic3d;
  ---Purpose: Returns the current texture plane name or NOTP_UNKNOWN
  -- when the plane is user defined.

  PlaneS (me; A, B, C, D : out ShortReal from Standard);
  ---Purpose: Returns the current texture plane S equation

  PlaneT (me; A, B, C, D : out ShortReal from Standard);
 ---Purpose: Returns   the current texture plane T equation

  TranslateS (me; theVal : out ShortReal from Standard);
  ---Purpose: Returns  the current texture S translation value

  TranslateT (me; theVal : out ShortReal from Standard);
  ---Purpose: Returns the current texture T translation value

  ScaleS (me; theVal : out ShortReal from Standard);
  ---Purpose: Returns the current texture S scale value

  ScaleT (me; theVal : out ShortReal from Standard);
  ---Purpose: Returns the current texture T scale value

  Rotation (me; theVal : out ShortReal from Standard);
  ---Purpose: Returns the current texture rotation angle

fields

  myPlaneName : NameOfTexturePlane from Graphic3d;

end Texture2Dplane;
