-- Created on: 2004-02-11
-- Created by: Sergey KUUL
-- Copyright (c) 2004-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MassMeasureWithUnit from StepBasic 

inherits MeasureWithUnit from StepBasic 

uses

	Real from Standard, 
	NamedUnit from StepBasic
is

	Create returns mutable MassMeasureWithUnit;
	---Purpose: Returns a MassMeasureWithUnit


end MassMeasureWithUnit;
