-- Created on: 1996-01-29
-- Created by: Christian CAILLET
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SignType  from IFSelect  inherits Signature

    ---Purpose : This Signature returns the cdl Type of an entity, under two
    --           forms :
    --           - complete dynamic type (package and class)
    --           - class type, without package name

uses CString, Transient, InterfaceModel

is

    Create (nopk : Boolean = Standard_False) returns mutable SignType;
    ---Purpose : Returns a SignType
    --           <nopk> false (D) : complete dynamic type (name = Dynamic Type)
    --           <nopk> true : class type without pk (name = Class Type)

    Value (me; ent : any Transient; model : InterfaceModel) returns CString;
    ---Purpose : Returns the Signature for a Transient object, as its Dynamic
    --           Type, with or without package name, according starting option

fields

    thenopk : Boolean;

end SignType;
