---Copyright:   Matra Datavision 1991

class Ax22d   from gp  inherits Storable
        --- Purpose :
        --  Describes a coordinate system in a plane (2D space).
        -- A coordinate system is defined by:
        -- -   its origin (also referred to as its "Location point"), and
        -- -   two orthogonal unit vectors, respectively, called the "X
        --   Direction" and the "Y Direction".
        --   A gp_Ax22d may be right-handed ("direct sense") or
        -- left-handed ("inverse" or "indirect sense").
        -- You use a gp_Ax22d to:
        -- - describe 2D geometric entities, in particular to position
        --   them. The local coordinate system of a geometric
        --   entity serves for the same purpose as the STEP
        --   function "axis placement two axes", or
        -- -   define geometric transformations.
        -- Note: we refer to the "X Axis" and "Y Axis" as the axes having:
        -- -   the origin of the coordinate system as their origin, and
        -- -   the unit vectors "X Direction" and "Y Direction",
        --   respectively, as their unit vectors. 

uses Ax2d  from gp,
     Dir2d  from gp,
     Pnt2d  from gp,
     Trsf2d from gp,
     Vec2d  from gp

raises ConstructionError from Standard

is

 
  Create  returns Ax22d;
        ---C++:inline
        --- Purpose : Creates an object representing the reference 
        --            co-ordinate system (OXY).
     
  Create (P : Pnt2d; Vx, Vy : Dir2d)   returns Ax22d
        ---C++:inline
        --- Purpose : 
        --  Creates a coordinate system with origin P and where:
        --   -   Vx is the "X Direction", and
        --   -   the "Y Direction" is orthogonal to Vx and
        --    oriented so that the cross products Vx^"Y
        --    Direction" and Vx^Vy have the same sign.
        -- Raises ConstructionError if Vx and Vy are parallel (same or opposite orientation).
    raises ConstructionError;
  
                            
  Create (P     : Pnt2d; 
    	  V     : Dir2d;
    	  Sense : Boolean from Standard = Standard_True)  returns Ax22d;
        ---C++:inline
	--- Purpose :
	--  Creates -   a coordinate system with origin P and "X Direction"
        --   V, which is:
        --   -   right-handed if Sense is true (default value), or
        --   -   left-handed if Sense is false

  Create (A : Ax2d; 
    	  Sense : Boolean from Standard = Standard_True)  returns Ax22d;
        ---C++:inline
	--- Purpose :
	--  Creates -   a coordinate system where its origin is the origin of
        --   A and its "X Direction" is the unit vector of A, which   is:
        --   -   right-handed if Sense is true (default value), or
        --   -   left-handed if Sense is false.

  SetAxis (me : in out; A1 : Ax22d)
        ---C++:inline
        --- Purpose :
        --  Assigns the origin and the two unit vectors of the
        -- coordinate system A1 to this coordinate system.
     is static;


  SetXAxis (me : in out; A1 : Ax2d)
        ---C++:inline
        --- Purpose :
        --  Changes the XAxis and YAxis ("Location" point and "Direction") 
        --  of <me>.
        --  The "YDirection" is recomputed in the same sense as before.
     is static;


  SetYAxis (me : in out; A1 : Ax2d) 
        ---C++:inline
        --- Purpose : Changes the XAxis and YAxis ("Location" point and "Direction") of <me>.
        --  The "XDirection" is recomputed in the same sense as before.
     is static;

  SetLocation (me : in out; P : Pnt2d)   is static;
        ---C++:inline
        --- Purpose :
        --  Changes the "Location" point (origin) of <me>.


  SetXDirection (me : in out; Vx : Dir2d)
        ---C++:inline
        --- Purpose :
        -- Assigns Vx to the "X Direction"  of
        -- this coordinate system. The other unit vector of this
        -- coordinate system is recomputed, normal to Vx ,
        -- without modifying the orientation (right-handed or
        -- left-handed) of this coordinate system.
     is static;


  SetYDirection(me : in out; Vy : Dir2d)
        ---C++:inline
        --- Purpose : Assignsr Vy to the  "Y Direction" of
        -- this coordinate system. The other unit vector of this
        -- coordinate system is recomputed, normal to Vy,
        -- without modifying the orientation (right-handed or
        -- left-handed) of this coordinate system.
     is static;


  XAxis (me)  returns Ax2d         is static;
        ---C++:inline
        --- Purpose : Returns an axis, for which
        -- -   the origin is that of this coordinate system, and
        -- -   the unit vector is either the "X Direction"  of this coordinate system.
        -- Note: the result is the "X Axis" of this coordinate system.

  YAxis (me)  returns Ax2d         is static;
        ---C++:inline
        --- Purpose : Returns an axis, for which
        --    -   the origin is that of this coordinate system, and
        -- - the unit vector is either the  "Y Direction" of this coordinate system.
        -- Note: the result is the "Y Axis" of this coordinate system.

  Location (me)  returns Pnt2d is static;
        ---C++:inline
        --- Purpose :
        --  Returns the "Location" point (origin) of <me>.
    	---C++: return const&


  XDirection (me)  returns Dir2d   is static;
        ---C++:inline
        --- Purpose :
        --  Returns the "XDirection" of <me>.
    	---C++: return const&

  YDirection(me)  returns Dir2d  is static;
        ---C++:inline
        --- Purpose :
        --  Returns the "YDirection" of <me>.
    	---C++: return const&


  Mirror (me : in out; P : Pnt2d)          is static;

  Mirrored (me; P : Pnt2d)  returns Ax22d    is static;

        --- Purpose :
        --  Performs the symmetrical transformation of an axis
        --  placement with respect to the point P which is the
        --  center of the symmetry.
        --- Warnings :
        --  The main direction of the axis placement is not changed.
        --  The "XDirection" and the "YDirection" are reversed. 
        --  So the axis placement stay right handed.


  Mirror (me : in out; A : Ax2d)         is static;

  Mirrored (me; A : Ax2d)  returns Ax22d   is static;

        --- Purpose :
        --  Performs the symmetrical transformation of an axis
        --  placement with respect to an axis placement which
        --  is the axis of the symmetry.
        --  The transformation is performed on the "Location"
        --  point, on the "XDirection" and "YDirection". 
        --  The resulting main "Direction" is the cross product between 
        --  the "XDirection" and the "YDirection" after transformation.



  Rotate (me : in out; P : Pnt2d; Ang : Real)         is static;
        ---C++:inline

  Rotated (me; P : Pnt2d; Ang : Real)  returns Ax22d    is static;
        ---C++:inline
        --- Purpose :
        --  Rotates an axis placement. <A1> is the axis of the
        --  rotation . Ang is the angular value of the rotation
        --  in radians.




  Scale (me : in out; P : Pnt2d; S : Real)             is static;
        ---C++:inline

  Scaled (me; P : Pnt2d; S : Real)  returns Ax22d       is static;
        ---C++:inline
        --- Purpose :
        --  Applies a scaling transformation on the axis placement.
        --  The "Location" point of the axisplacement is modified.
        --- Warnings :
        --  If the scale <S> is negative :
        --   . the main direction of the axis placement is not changed.
        --   . The "XDirection" and the "YDirection" are reversed. 
        --  So the axis placement stay right handed.
              

 

  Transform (me : in out; T : Trsf2d)                  is static;
        ---C++:inline

  Transformed (me; T : Trsf2d)   returns Ax22d           is static;
        ---C++:inline
        --- Purpose :  
        --  Transforms an axis placement with a Trsf.
        --  The "Location" point, the "XDirection" and the
        --  "YDirection" are transformed with T.  The resulting
        --  main "Direction" of <me> is the cross product between 
        --  the "XDirection" and the "YDirection" after transformation.


  Translate (me : in out; V : Vec2d)            
        ---C++:inline
      is static;

  Translated (me; V : Vec2d)  returns Ax22d  is static;
        ---C++:inline
        --- Purpose : 
        --  Translates an axis plaxement in the direction of the vector
        --  <V>. The magnitude of the translation is the vector's magnitude.



      
  Translate (me : in out; P1, P2 : Pnt2d)      
        ---C++:inline
        is static;

  Translated (me; P1, P2 : Pnt2d)   returns Ax22d        is static;
        ---C++:inline
        --- Purpose :
        --  Translates an axis placement from the point <P1> to the 
        --  point <P2>.




fields

   point  : Pnt2d;
   vydir : Dir2d;
   vxdir : Dir2d;

end;
