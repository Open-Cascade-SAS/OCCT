-- Created on: 1994-10-24
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class DrawableP3D from TestTopOpeDraw inherits Marker3D from Draw

    ---Purpose: 

uses  

    Color           from Draw,
    Display         from Draw,
    Text3D          from Draw,
    MarkerShape     from Draw,
    CString         from Standard,
    Pnt             from gp,
    Pnt2d           from gp,
    Circ            from gp
    
is

    Create (P : Pnt from gp; PColor : Color from Draw;
    	    moveX : Real = 0.0; moveY : Real = 0.0)
    returns mutable DrawableP3D from TestTopOpeDraw;

    Create (P : Pnt from gp; PColor : Color from Draw;
    	    Text : CString; TextColor : Color from Draw;
    	    moveX : Real = 0.0; moveY : Real = 0.0)
    returns mutable DrawableP3D from TestTopOpeDraw;

    Create (P : Pnt from gp; T : MarkerShape from Draw; PColor : Color from Draw;
    	    Text : CString from Standard; TextColor : Color from Draw;
	    Size : Integer from Standard = 2;
    	    moveX : Real = 0.0; moveY : Real = 0.0)
    returns mutable DrawableP3D from TestTopOpeDraw;

    Create (P : Pnt from gp; T : MarkerShape from Draw; 
    	    PColor : Color from Draw;
    	    Text : CString from Standard; TextColor : Color from Draw;
    	    Tol : Real from Standard;
    	    moveX : Real = 0.0; moveY : Real = 0.0)
    returns mutable DrawableP3D from TestTopOpeDraw;

    ChangePnt(me : mutable; P : Pnt);
    
    DrawOn(me; dis : in out Display from Draw)
    is redefined;
    
fields

    myPnt    : Pnt from gp;
    myText   : CString from Standard;
    myTextColor : Color from Draw;
    myMoveX  : Real from Standard;
    myMoveY  : Real from Standard;

    myText3D : Text3D from Draw;

end DrawableP3D;
