-- File:	GeomToStep_MakeCircle.cdl
-- Created:	Mon Jun 14 15:18:28 1993
-- Author:	Martine LANGLOIS
--		<mla@mastox>
---Copyright:	 Matra Datavision 1993

class MakeCircle from GeomToStep inherits Root from GeomToStep

    ---Purpose: This class implements the mapping between classes 
    --          Circle from Geom, and Circ from gp, and the class
    --          Circle from StepGeom which describes a circle from
    --          Prostep. 
  
uses Circ from gp,
     Circ2d from gp,
     Circle from Geom,
     Circle from Geom2d,
     Circle from StepGeom
     
raises NotDone from StdFail
     
is 

Create ( C : Circ from gp ) returns MakeCircle;

Create ( C : Circle from Geom ) returns MakeCircle;

Create ( C : Circle from Geom2d ) returns MakeCircle;

Value (me) returns Circle from StepGeom
    raises NotDone
    is static;
    ---C++: return const&
    
fields

    theCircle : Circle from StepGeom;
    	-- The solution from StepGeom
    	
end MakeCircle;


