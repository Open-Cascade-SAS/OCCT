-- Created on: 1993-06-24
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class InterferenceTool from TopOpeBRepDS
     
uses

    Curve        from Geom2d,
    Orientation  from TopAbs,
    Transition   from TopOpeBRepDS,
    Interference from TopOpeBRepDS,
    Config       from TopOpeBRepDS,
    Kind         from TopOpeBRepDS
    
is

    MakeEdgeInterference(myclass;
			 T : Transition from TopOpeBRepDS;
	      	    	 SK : Kind; SI : Integer;
   	    	    	 GK : Kind; GI : Integer;
	      	    	 P : Real from Standard) 
    returns any Interference from TopOpeBRepDS;

    MakeCurveInterference(myclass;
    	     		  T : Transition from TopOpeBRepDS;
	      	    	  SK : Kind; SI : Integer;
    	    	    	  GK : Kind; GI : Integer;
	      	    	  P : Real from Standard) 
    returns any Interference from TopOpeBRepDS;

    DuplicateCurvePointInterference(myclass; I : Interference from TopOpeBRepDS)
    ---Purpose :  duplicate I in a new interference with Complement() transition.
    returns any Interference from TopOpeBRepDS;

    MakeFaceCurveInterference(myclass;
		    	      Transition : Transition from TopOpeBRepDS;
	      	    	      FaceI, CurveI : Integer from Standard;
	      	    	      PC : Curve from Geom2d) 
    returns any Interference from TopOpeBRepDS;

    MakeSolidSurfaceInterference(myclass;
    	      	    	    	 Transition : Transition from TopOpeBRepDS;
	      	    	    	 SolidI, SurfaceI : Integer from Standard)
    returns any Interference from TopOpeBRepDS;

    MakeEdgeVertexInterference(myclass;
    	      	    	       Transition : Transition from TopOpeBRepDS;
	      	    	       EdgeI, VertexI : Integer from Standard;
    	      	    	       VertexIsBound : Boolean from Standard;
    	      	    	       Config : Config from TopOpeBRepDS;
    	      	    	       param : Real from Standard)
    returns any Interference from TopOpeBRepDS;

    MakeFaceEdgeInterference(myclass;
    	      	    	       Transition : Transition from TopOpeBRepDS;
	      	    	       FaceI, EdgeI : Integer from Standard;
    	      	    	       EdgeIsBound : Boolean from Standard;
    	      	    	       Config : Config from TopOpeBRepDS)
    returns any Interference from TopOpeBRepDS;

    Parameter(myclass; CPI : Interference from TopOpeBRepDS)
    returns Real from Standard;

    Parameter(myclass; CPI : Interference from TopOpeBRepDS; 
                       Par : Real from Standard);
    
end InterferenceTool from TopOpeBRepDS;
