-- Created on: 1991-12-02
-- Created by: Laurent PAINNOT
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MultiPoint from AppParCurves
    	---Purpose: This class describes Points composing a MultiPoint.
    	--          These points can be 2D or 3D. The user must first give the 
    	--          3D Points and then the 2D Points.
   	--          They are Poles of a Bezier Curve.
    	-- This class is used either to define data input or
    	-- results when performing the approximation of several lines in parallel.


uses Pnt                from gp,
     Pnt2d              from gp,
     Vec                from gp,
     Vec2d              from gp,
     Array1OfPnt        from TColgp,
     Array1OfPnt2d      from TColgp,
     HArray1OfPnt       from TColgp,
     HArray1OfPnt2d     from TColgp,
     OStream            from Standard,
     TShared            from MMgt
     
raises OutOfRange     from Standard,
       DimensionError from Standard

is

    Create returns MultiPoint;
    	---Purpose: creates an indefinite MultiPoint.


    Create(NbPoints, NbPoints2d: Integer)
    	---Purpose: constructs a set of Points used to approximate a 
    	--          Multiline.
    	--          These Points can be of 2 or 3 dimensions.
    	--          Points will be initialized with SetPoint and SetPoint2d.
    	--          NbPoints is the number of 3D Points.
    	--          NbPoints2d is the number of 2D Points.

    returns MultiPoint from AppParCurves;


    Create(tabP: Array1OfPnt)
    	---Purpose: creates a MultiPoint only composed of 3D points.

    returns MultiPoint from AppParCurves;


    Create(tabP2d: Array1OfPnt2d)
    	---Purpose: creates a MultiPoint only composed of 2D points.

    returns MultiPoint from AppParCurves;
    
		
    Create(tabP: Array1OfPnt; tabP2d: Array1OfPnt2d)
    	---Purpose: constructs a set of Points used to approximate a 
    	--          Multiline.
    	--          These Points can be of 2 or 3 dimensions.
    	--          Points will be initialized with SetPoint and SetPoint2d.
    	--          NbPoints is the total number of Points.
   
    returns MultiPoint from AppParCurves;   

    ---C++: alias "  Standard_EXPORT virtual ~AppParCurves_MultiPoint();"
    
    SetPoint(me: in out; Index: Integer; Point: Pnt)
    	---Purpose: the 3d Point of range Index of this MultiPoint is 
    	--          set to <Point>.
    	--          An exception is raised if Index < 0 or 
    	--          Index > number of 3d Points.

    raises OutOfRange from Standard
    is static;
    


    Point(me; Index: Integer)
    	---Purpose: returns the 3d Point of range Index.
    	--          An exception is raised if Index < 0 or
    	--          Index < number of 3d Points.
    	---C++: return const&
    
    returns Pnt from gp
    raises OutOfRange from Standard
    is static;
    
    
    SetPoint2d(me: in out; Index: Integer; Point: Pnt2d)
    	---Purpose: The 2d Point of range Index is set to <Point>.
    	--          An exception is raised if Index > 3d Points or 
    	--          Index > total number of Points.
    
    raises OutOfRange from Standard,
    	   DimensionError from Standard
    is static;
    

    Point2d(me; Index: Integer)
    	---Purpose: returns the 2d Point of range Index.
    	--          An exception is raised if index <= number of 
    	--          3d Points or Index > total number of Points.
    	---C++: return const&

    returns Pnt2d from gp
    raises OutOfRange from Standard
    is static;



    Dimension(me; Index: Integer)
    	---Purpose: returns the dimension of the point of range Index.
    	--          An exception is raised if Index <0 or Index > NbCurves.
    	---C++: inline

    returns Integer
    raises OutOfRange from Standard
    is static;
    

    NbPoints(me)
    	---Purpose: returns the number of points of dimension 3D.
    	---C++: inline

    returns Integer
    is static;
	
			    
    NbPoints2d(me)
    	---Purpose: returns the number of points of dimension 2D.
    	---C++: inline

    returns Integer
    is static;


    Transform(me: in out; CuIndex: Integer; x, dx, y, dy, z, dz: Real)
        ---Purpose: Applies a transformation to the curve of range 
        --          <CuIndex>.
        --          newx = x + dx*oldx
        --          newy = y + dy*oldy    for all points of the curve.
        --          newz = z + dz*oldz

    raises OutOfRange from Standard
    is static;


    Transform2d(me: in out; CuIndex: Integer; x, dx, y, dy: Real)
        ---Purpose: Applies a transformation to the Curve of range 
        --          <CuIndex>.
        --          newx = x + dx*oldx
        --          newy = y + dy*oldy    for all points of the curve.

    raises OutOfRange from Standard
    is static;


    Dump(me; o: in out OStream)
    	---Purpose: Prints on the stream o information on the current 
    	--          state of the object.
    	--          Is used to redefine the operator <<.
    is virtual;

fields

ttabPoint  : TShared from MMgt is protected;
ttabPoint2d: TShared from MMgt is protected;
nbP        : Integer is protected;
nbP2d      : Integer is protected;

end MultiPoint;

