-- Created on: 2001-09-26
-- Created by: Julia DOROVSKIKH
-- Copyright (c) 2001-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ADriverTable from XmlMDF inherits TShared from MMgt

        ---Purpose: A driver table is an object building links between
        --          object types and object drivers. In the
        --          translation process, a driver table is asked to
        --          give a translation driver for each current object
        --          to be translated.

uses
    Type               from Standard,
    MapTransientHasher from TColStd,
    ADriver            from XmlMDF,    
    TypeADriverMap     from XmlMDF

is
    Create returns ADriverTable from XmlMDF;
        ---Purpose: Creates a mutable ADriverTable from XmlMDF.

    AddDriver(me : mutable; anHDriver : ADriver from XmlMDF);
        ---Purpose: Sets a translation driver: <aDriver>.

    GetDrivers(me)
        returns TypeADriverMap from XmlMDF;
        ---Purpose: Gets a map of drivers. 
        ---C++: return const &

    GetDriver(me; aType     : Type from Standard;
                  anHDriver : in out ADriver from XmlMDF)
        returns Boolean from Standard;
        ---Purpose: Gets a driver <aDriver> according to <aType>
        --          
        --          Returns True if a driver is found; false otherwise.

fields
    myMap : TypeADriverMap from XmlMDF;

end ADriverTable;
