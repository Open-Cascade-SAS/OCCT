-- Created on: 2003-06-04
-- Created by: Galina KULIKOVA
-- Copyright (c) 2003-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class CommonDatum from StepDimTol
inherits CompositeShapeAspect from StepRepr

    ---Purpose: Representation of STEP entity CommonDatum

uses
    HAsciiString from TCollection,
    ProductDefinitionShape from StepRepr,
    Logical from StepData,
    Datum from StepDimTol

is
    Create returns CommonDatum from StepDimTol;
	---Purpose: Empty constructor

    Init (me: mutable; aShapeAspect_Name: HAsciiString from TCollection;
                       aShapeAspect_Description: HAsciiString from TCollection;
                       aShapeAspect_OfShape: ProductDefinitionShape from StepRepr;
                       aShapeAspect_ProductDefinitional: Logical from StepData;
                       aDatum_Name: HAsciiString from TCollection;
                       aDatum_Description: HAsciiString from TCollection;
                       aDatum_OfShape: ProductDefinitionShape from StepRepr;
                       aDatum_ProductDefinitional: Logical from StepData;
                       aDatum_Identification: HAsciiString from TCollection);
	---Purpose: Initialize all fields (own and inherited)

    Datum (me) returns Datum from StepDimTol;
	---Purpose: Returns data for supertype Datum
    SetDatum (me: mutable; Datum: Datum from StepDimTol);
	---Purpose: Set data for supertype Datum

fields
    theDatum: Datum from StepDimTol; -- supertype

end CommonDatum;
