-- Created on: 1999-02-12
-- Created by: Andrey BETENEV
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class TranslateCurveBoundedSurface from StepToTopoDS 
    inherits Root from StepToTopoDS
    ---Purpose: Translate curve_bounded_surface into TopoDS_Face

uses
    TransientProcess from Transfer,
    CurveBoundedSurface from StepGeom,
    Face                from TopoDS

is
    Create returns TranslateCurveBoundedSurface;
        ---Purpose: Create empty tool

    Create (CBS: CurveBoundedSurface from StepGeom;
    	    TP: TransientProcess from Transfer)
    	returns TranslateCurveBoundedSurface;
        ---Purpose: Translate surface
	
    Init (me: in out;
          CBS: CurveBoundedSurface from StepGeom;
    	  TP: TransientProcess from Transfer)
    	returns Boolean;
        ---Purpose: Translate surface
	
    Value (me) returns Face from TopoDS;
        ---Purpose: Returns result of last translation or null wire if failed.
	---C++: return const &

fields

    myFace: Face from TopoDS;

end TranslateCurveBoundedSurface;
