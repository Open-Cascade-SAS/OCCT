-- Created on: 1999-06-17
-- Created by: data exchange team
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



private class ConvertToBSpline from ShapeCustom inherits Modification from BRepTools

    	---Purpose: implement a modification for BRepTools
	--          Modifier algortihm. Converts Surface of
	--          Linear Exctrusion, Revolution and Offset
	--          surfaces into BSpline Surface according to
	--          flags.
	
uses

    Face     from TopoDS,
    Edge     from TopoDS,
    Vertex   from TopoDS,
    Shape    from GeomAbs,
    Surface  from Geom,
    Curve    from Geom,
    Curve    from Geom2d,
    Pnt      from gp,
    Location from TopLoc
is

    Create returns mutable ConvertToBSpline from ShapeCustom;
    
    SetExtrusionMode(me: mutable; extrMode: Boolean);
    	---Purpose: Sets mode for convertion of Surfaces of Linear
	--          extrusion.
    
    SetRevolutionMode(me: mutable; revolMode: Boolean);
    	---Purpose: Sets mode for convertion of Surfaces of Revolution.

    SetOffsetMode(me: mutable; offsetMode: Boolean);
    	---Purpose: Sets mode for convertion of Offset surfaces.
    
    SetPlaneMode(me: mutable; planeMode: Boolean);
    	---Purpose: Sets mode for convertion of Plane surfaces.
    
    NewSurface(me: mutable; F  :     Face     from TopoDS;
                            S  : out Surface  from Geom;
		            L  : out Location from TopLoc;
		            Tol: out Real     from Standard;
                            RevWires : out Boolean from Standard;
                            RevFace  : out Boolean from Standard)
    returns Boolean from Standard;
      	---Purpose: Returns Standard_True if the face <F> has  been
	--          modified. In this case, <S> is the new geometric
	--          support of the face, <L> the new location,  <Tol>
	--          the new tolerance.  Otherwise, returns
	--          Standard_False, and <S>, <L>, <Tol> are  not
	--          significant.
    
    NewCurve(me: mutable; E  :     Edge     from TopoDS;
                          C  : out Curve    from Geom;
		          L  : out Location from TopLoc;
		          Tol: out Real     from Standard)
    returns Boolean from Standard;
	---Purpose: Returns Standard_True  if  the edge  <E> has  been
	--          modified.  In this case,  <C> is the new geometric
	--          support of the  edge, <L> the  new location, <Tol>
	--          the         new    tolerance.   Otherwise, returns
	--          Standard_False,    and  <C>,  <L>,   <Tol> are not
	--          significant.

    NewPoint(me: mutable; V  :     Vertex   from TopoDS;
                          P  : out Pnt      from gp;
		          Tol: out Real     from Standard)
    returns Boolean from Standard;
	---Purpose: Returns  Standard_True if the  vertex <V> has been
	--          modified.  In this  case, <P> is the new geometric
	--          support of the vertex,   <Tol> the new  tolerance.
	--          Otherwise, returns Standard_False, and <P>,  <Tol>
	--          are not significant.

    NewCurve2d(me: mutable; E    :     Edge     from TopoDS;
                            F    :     Face     from TopoDS;
                            NewE :     Edge     from TopoDS;
                            NewF :     Face     from TopoDS;
                            C    : out Curve    from Geom2d;
		            Tol  : out Real     from Standard)
    returns Boolean from Standard;
    	---Purpose: Returns Standard_True if  the edge  <E> has a  new
	--          curve on surface on the face <F>.In this case, <C>
	--          is the new geometric support of  the edge, <L> the
	--          new location, <Tol> the new tolerance.
	--          
	--          Otherwise, returns  Standard_False, and <C>,  <L>,
	--          <Tol> are not significant.
	--          
	--          <NewE> is the new  edge created from  <E>.  <NewF>
	--          is the new face created from <F>. They may be usefull.

    NewParameter(me: mutable; V  :     Vertex from TopoDS;
                              E  :     Edge   from TopoDS;
                              P  : out Real   from Standard;
  		              Tol: out Real   from Standard)
    returns Boolean from Standard;
	---Purpose: Returns Standard_True if the Vertex  <V> has a new
	--          parameter on the  edge <E>. In  this case,  <P> is
	--          the parameter,    <Tol>  the     new    tolerance.
	--          Otherwise, returns Standard_False, and <P>,  <Tol>
	--          are not significant.

    Continuity(me: mutable; E          : Edge from TopoDS;
    	                    F1,F2      : Face from TopoDS;
			    NewE       : Edge from TopoDS;
			    NewF1,NewF2: Face from TopoDS)
    returns Shape from GeomAbs;
	---Purpose: Returns the  continuity of  <NewE> between <NewF1>
	--          and <NewF2>.
	--          
	--          <NewE> is the new  edge created from <E>.  <NewF1>
	--          (resp. <NewF2>) is the new  face created from <F1>
	--          (resp. <F2>).
    
    IsToConvert(me; S :    Surface from Geom;
    	    	    SS:out Surface from Geom)
    returns Boolean is private;

fields

    myExtrMode  : Boolean;
    myRevolMode : Boolean;
    myOffsetMode: Boolean;
    myPlaneMode : Boolean;
    
end ConvertToBSpline;
