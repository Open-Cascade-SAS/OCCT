-- Created on: 2001-04-13
-- Created by: Peter KURNEV
-- Copyright (c) 2001-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class ConnexityBlock from BOP 

	---Purpose: 
    	---  Auxiliary class to store data about set  
    	---  of connex shapes 
	--- 
	
uses
    ListOfShape               from TopTools,
    IndexedMapOfOrientedShape from TopTools

is 
    Create
    	returns ConnexityBlock from BOP; 
    	---Purpose:  
    	--- Empty constructor; 
    	---
    SetShapes    (me:out; 
        anEdges: ListOfShape from TopTools); 
    	---Purpose:  
    	--- Modifier
    	---
    SetShapes    (me:out; 
    	nEdges: IndexedMapOfOrientedShape from TopTools); 
    	---Purpose:  
    	--- Modifier
    	---
    SetRegularity(me:out;  
    		   aFlag:Boolean from Standard);    	    	    
    	---Purpose:  
    	--- Modifier
    	---
    Shapes  (me) 
    	returns ListOfShape from TopTools; 
    	---C++:  return const &  
    	---Purpose:  
    	--- Selector
    	---
    IsRegular(me) 
        returns Boolean from Standard;  
    	---Purpose:  
    	--- Selector 
    	--- Returns TRUE if all elements in the block are 
    	--- biconnexity     	
    	---
    
fields
    
    myRegularity  :  Boolean from Standard;  
    myShapes      :  ListOfShape from TopTools; 

end ConnexityBlock;
