-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Person from StepBasic 

inherits TShared from MMgt

uses

	HAsciiString from TCollection, 
	HArray1OfHAsciiString from Interface, 
	Boolean from Standard
is

	Create returns mutable Person;
	---Purpose: Returns a Person

	Init (me : mutable;
	      aId : mutable HAsciiString from TCollection;
	      hasAlastName : Boolean from Standard;
	      aLastName : mutable HAsciiString from TCollection;
	      hasAfirstName : Boolean from Standard;
	      aFirstName : mutable HAsciiString from TCollection;
	      hasAmiddleNames : Boolean from Standard;
	      aMiddleNames : mutable HArray1OfHAsciiString from Interface;
	      hasAprefixTitles : Boolean from Standard;
	      aPrefixTitles : mutable HArray1OfHAsciiString from Interface;
	      hasAsuffixTitles : Boolean from Standard;
	      aSuffixTitles : mutable HArray1OfHAsciiString from Interface) is virtual;

	-- Specific Methods for Field Data Access --

	SetId(me : mutable; aId : mutable HAsciiString);
	Id (me) returns mutable HAsciiString;
	SetLastName(me : mutable; aLastName : mutable HAsciiString);
	UnSetLastName (me:mutable);
	LastName (me) returns mutable HAsciiString;
	HasLastName (me) returns Boolean;
	SetFirstName(me : mutable; aFirstName : mutable HAsciiString);
	UnSetFirstName (me:mutable);
	FirstName (me) returns mutable HAsciiString;
	HasFirstName (me) returns Boolean;
	SetMiddleNames(me : mutable; aMiddleNames : mutable HArray1OfHAsciiString);
	UnSetMiddleNames (me:mutable);
	MiddleNames (me) returns mutable HArray1OfHAsciiString;
	HasMiddleNames (me) returns Boolean;
	MiddleNamesValue (me; num : Integer) returns mutable HAsciiString;
	NbMiddleNames (me) returns Integer;
	SetPrefixTitles(me : mutable; aPrefixTitles : mutable HArray1OfHAsciiString);
	UnSetPrefixTitles (me:mutable);
	PrefixTitles (me) returns mutable HArray1OfHAsciiString;
	HasPrefixTitles (me) returns Boolean;
	PrefixTitlesValue (me; num : Integer) returns mutable HAsciiString;
	NbPrefixTitles (me) returns Integer;
	SetSuffixTitles(me : mutable; aSuffixTitles : mutable HArray1OfHAsciiString);
	UnSetSuffixTitles (me:mutable);
	SuffixTitles (me) returns mutable HArray1OfHAsciiString;
	HasSuffixTitles (me) returns Boolean;
	SuffixTitlesValue (me; num : Integer) returns mutable HAsciiString;
	NbSuffixTitles (me) returns Integer;

fields

	id : HAsciiString from TCollection;
	lastName : HAsciiString from TCollection;   -- OPTIONAL can be NULL
	firstName : HAsciiString from TCollection;   -- OPTIONAL can be NULL
	middleNames : HArray1OfHAsciiString from Interface;   -- OPTIONAL can be NULL
	prefixTitles : HArray1OfHAsciiString from Interface;   -- OPTIONAL can be NULL
	suffixTitles : HArray1OfHAsciiString from Interface;   -- OPTIONAL can be NULL
	hasLastName : Boolean from Standard;
	hasFirstName : Boolean from Standard;
	hasMiddleNames : Boolean from Standard;
	hasPrefixTitles : Boolean from Standard;
	hasSuffixTitles : Boolean from Standard;

end Person;
