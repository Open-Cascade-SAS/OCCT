-- Created on: 1993-01-26
-- Created by: Isabelle GRIGNON
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred generic class CurveTool from IntImp (Curve as any)

	---Purpose: Template class for the methods on a curve.
	--          It is possible to implement this class with
	--          an instantiation of the CurveTool from Adaptor3d.

uses Pnt from gp,
     Vec from gp


is

    FirstParameter(myclass;C : Curve ) returns Real;
    
    LastParameter(myclass;C : Curve ) returns Real;

    Resolution(myclass; C : Curve; Tol3d: Real from Standard)
    
        ---Purpose :  Returns the parametric  resolution corresponding
        --         to the space resolution Tol3d.

    	returns Real from Standard;

end CurveTool;
