-- Created on: 1993-02-10
-- Created by: Mireille MERCIEN
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class HExtendedString from PCollection 
	inherits Persistent    
	   
        ---Purpose: Describes a persistent Unicode character string
    	-- of a variable length.


uses       VArrayOfExtCharacter from DBC,
           ExtendedString from TCollection,
           HAsciiString from PCollection 
	    

    raises OutOfRange from Standard, 
           NegativeValue from Standard,
    	   NumericError from Standard
is
		

	Create(S : ExtendedString from TCollection) 
            returns mutable HExtendedString from PCollection;
		---Purpose: Creation and initialization with the string S from
		-- TCollection.

	Create(C : ExtCharacter from Standard)
            returns mutable HExtendedString from PCollection;
		---Purpose: Creation and initialisation with the character C

	Create(S : HExtendedString from PCollection;
    	       FromIndex, ToIndex : Integer from Standard) 
	    returns mutable HExtendedString from PCollection
	    raises NegativeValue from Standard;
                ---Purpose: Creation of a sub-string of the string S
                -- the sub-string starts at the index Fromindex and ends
                -- at the index ToIndex.
                -- Raises an exception if ToIndex is less than FromIndex 

        Create( astring : CString)
            returns mutable HExtendedString from PCollection;
        ---Purpose: Creation by converting a CString to an extended string. 
	
        Create(S : HAsciiString from PCollection)
            returns mutable HExtendedString from PCollection;
	---Purpose: Creation by converting a normal Ascii string to an extended string. 
	
	Append(me : mutable; S : HExtendedString from PCollection);
        ---Level: Public
	---Purpose: Pushing a string at the end of the string me.

	Center(me : mutable; Width : Integer from Standard;
      	       Filler : ExtCharacter from Standard) 
	raises NegativeValue from Standard;
        ---Level: Public
	---Purpose: Center.
        -- Length becomes equal to Width and the new characters are
        -- equal to Filler.
        -- Raises an exception if Width is less than zero.
	-- If Width < Length nothing happens.

	ChangeAll(me : mutable; C, NewC : ExtCharacter from Standard);
        ---Level: Public
        ---Purpose: Substitutes all the characters equal to C by NewC in the
        -- string <me>.

	Clear(me : mutable);
        ---Level: Public
	---Purpose: Removes all characters in the string <me>.
        -- Length is equal to zero now.

        Convert(me) returns ExtendedString from TCollection;
        ---Level: Public
        ---Purpose: Converts a persistent HExtendedString to a non
        -- persistent ExtendedString.

	FirstLocationInSet(me; Set : HExtendedString from PCollection;
                                 FromIndex : Integer from Standard; 
                                 ToIndex   : Integer from Standard)
        returns Integer
	raises OutOfRange from Standard;
        ---Level: Public
        ---Purpose: Returns the index of the first character of <Set> founded in <me>.
        -- The search begins to the index FromIndex and ends to the index ToIndex.
        -- Returns zero if failure.
        -- Raises an exception if FromIndex or ToIndex is out of range.

	FirstLocationNotInSet(me; Set : HExtendedString from PCollection;
                              FromIndex : Integer; 
                              ToIndex   : Integer) 
        returns Integer
	raises OutOfRange from Standard;
                ---Level: Public
                ---Purpose: Returns the index of the first character of <me> 
                -- that is not present in the set <Set>.
                -- The search begins to the index FromIndex and ends to the
                -- the index ToIndex in <me>. Returns zero if failure.
                -- Raises an exception if FromIndex or ToIndex is out of range.

	InsertAfter(me : mutable; 
                    Index : Integer; 
                    S : HExtendedString from PCollection)
	raises OutOfRange from Standard;
                ---Level: Public
		---Purpose: Pushing a string after a specific index in the string <me>.
                -- Raises an exception if Index is out of bounds.

	InsertBefore(me : mutable; Index : Integer; 
                     S : HExtendedString from PCollection)
        raises OutOfRange from Standard;
                ---Level: Public
		---Purpose: Pushing a string before a specific index in the string <me>.
                -- Raises an exception if Index is out of bounds.

        IsAscii(me) returns Boolean;
        ---Level: Public
	---Purpose: Returns True if the string <me> is in the "Ascii range".
     
        IsDifferent (me ; other : HExtendedString) returns Boolean;
        ---Level: Public
        ---Purpose: Test if characters are different between <me> and <other>.
   
	IsEmpty(me) returns Boolean from Standard;
        ---Level: Public
	---Purpose: Returns True if the string <me> contains zero character.

        IsGreater (me ; other : HExtendedString from PCollection) 
        returns Boolean;
        ---Level: Public
        ---Purpose: Returns TRUE if <me> is greater than <other>.

        IsLess (me ; other : HExtendedString from PCollection) 
        returns Boolean;
        ---Level: Public
        ---Purpose: Returns TRUE if <me> is less than <other>.

	IsSameString(me; S : HExtendedString from PCollection)
	returns Boolean from Standard;
                ---Level: Advanced
                ---Purpose: Returns True if two strings are equal.
                -- The comparison is case sensitive if the flag is set.
  
	LeftAdjust(me : mutable)
        raises OutOfRange from Standard;
        ---Level: Public
        ---Purpose: Removes all space characters in the begining of the string.
        -- Raises an exception if the string <me> is not in the "Ascii range".

	LeftJustify(me : mutable; Width : Integer; 
                    Filler : ExtCharacter from Standard) 
	raises NegativeValue from Standard;
                ---Level: Public
		---Purpose: Left justify.
                -- Length becomes equal to Width and the new characters are
                -- equal to Filler.
                -- If Width < Length nothing happens.
                -- Raises an exception if Width is less than zero.

	Length(me) returns Integer;
        ---Level: Public
	---Purpose: Number of characters of the String

	Location(me; N : Integer; C : ExtCharacter from Standard; 
                    FromIndex : Integer; 
                    ToIndex   : Integer) 
        returns Integer
	raises OutOfRange from Standard;
                ---Level: Public
                ---Purpose: Returns the index of the nth occurence of the character C
                -- in the string <me> from the starting index FromIndex to the
                -- ending index ToIndex. Returns zero if failure.
                -- Raises an exception if FromIndex or ToIndex is out of range

	Location(me; S : HExtendedString from PCollection;
                    FromIndex : Integer; 
                    ToIndex   : Integer) 
        returns Integer
	raises OutOfRange from Standard;
                ---Level: Public
                ---Purpose: Returns an index in the string <me> of the first occurence
                -- of the string S in the string <me> from the starting index.
                -- FromIndex to the ending index ToIndex.
                -- Returns zero if failure.
                -- Raises an exception if FromIndex or ToIndex is out of range.

	Prepend(me : mutable; S : HExtendedString from PCollection);
                ---Level: Public
		---Purpose: Pushing a string at the begining of the string <me>.

	Print(me ; S : in out OStream);
        ---Level: Public
	---Purpose: Prints the content of <me> on the stream S.

	Remove(me : mutable; Index : Integer) 
        ---Level: Public
	---Purpose: Removes the character located at the index Index in the string.
        -- Raises an exception if Index is out of bounds.
	raises OutOfRange from Standard;

	Remove(me : mutable; FromIndex, ToIndex : Integer) 
	---Level: Public
	---Purpose: Removes all the characters from the index FromIndex to the
        -- index ToIndex.
        -- Raises an exception if FromIndex or ToIndex is out of bounds.
        raises OutOfRange from Standard;

	RemoveAll(me : mutable; C : ExtCharacter from Standard);
	---Level: Public
        ---Purpose: Removes all the occurences of the character C in the string.

	RightAdjust(me : mutable)
	raises OutOfRange from Standard;
	---Level: Public
        ---Purpose: Removes all space characters at the end of the string.
        -- Raises an exception if the string <me> is not in the Unicod "Ascii range".

	RightJustify(me : mutable; Width : Integer;
    	    	    	    	    	 Filler : ExtCharacter from Standard) 
		raises NegativeValue from Standard;
	        ---Level: Public
		---Purpose: Right justify.
                -- Length becomes equal to Width and the new characters are
                -- equal to Filler.
                -- If Width < Length nothing happens.
                -- Raises an exception if Width is less than zero.

	SetValue(me : mutable; Index : Integer; 
                 C : ExtCharacter from Standard) 
	raises OutOfRange from Standard;
	        ---Level: Public
                ---Purpose: Substitutes the character located to the position Index
                -- by the character C.
                -- Raises an exception if the Index is out of bounds

	SetValue(me : mutable; Index : Integer;
                 S : HExtendedString from PCollection) 
		raises OutOfRange from Standard;
	        ---Level: Public
                ---Purpose: Substitutes from the index Index to the end by the string S.
                -- Raises an exception if Index is out of bounds.

	Split(me : mutable; Index  : Integer) 
	---Level: Public
        ---Purpose: Splits a string of characters into two sub-strings.
	returns mutable HExtendedString from PCollection
	raises OutOfRange from Standard;

	SubString(me; FromIndex, ToIndex : Integer) 
	---Level: Public
        ---Purpose: Creation of a sub-string of the string <me>.
        -- The sub-string starts to the index FromIndex and ends
        -- to the index ToIndex.
        -- Raises an exception if ToIndex or FromIndex is out of bounds.
	returns mutable HExtendedString from PCollection
	raises OutOfRange from Standard;

	UsefullLength(me) returns Integer
        raises OutOfRange from Standard;
	---Level: Public
        ---Purpose: Length of the string ignoring all spaces (' ') and the 
        -- control character at the end.
        -- Raises an exception if the string <me> is not in the "Ascii range".

	Value(me; Index : Integer) returns ExtCharacter from Standard 
	raises OutOfRange from Standard;
         	---Level: Public
		---Purpose: Returns the character of index Index of the string.
                ---Example: me = "abcd", Index = 2, Value returns 'b'

     	ShallowDump (me; s: in out OStream) 
            	is redefined;
 		---Level: Advanced
   	    	---C++: function call


	Assign(me : mutable ;TheData : VArrayOfExtCharacter) is private;
	        ---Level: Internal
	    	---Purpose : Assigns the field of the current structure with
	    	--  the given value.

fields
   Data : VArrayOfExtCharacter from DBC;
end HExtendedString;
