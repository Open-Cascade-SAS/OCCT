-- Created on: 2007-08-22
-- Created by: Sergey ZARITCHNY
-- Copyright (c) 2007-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class AsciiString from PDataStd inherits Attribute from PDF

	---Purpose: Persistance attribute of  TDataStd_AsciiString

uses  HAsciiString from PCollection

is
    Create returns mutable  AsciiString from  PDataStd;
    
    
    Create (V : HAsciiString from PCollection) 
    returns mutable  AsciiString from PDataStd;
    
    
    Get (me) returns HAsciiString from PCollection;
    
    
    Set (me : mutable; V : HAsciiString from PCollection);
    
fields

    myValue : HAsciiString from PCollection;


end AsciiString;
