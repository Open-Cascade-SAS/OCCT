-- Created by: Peter KURNEV
-- Copyright (c) 2010-2012 OPEN CASCADE SAS
-- Copyright (c) 2007-2010 CEA/DEN, EDF R&D, OPEN CASCADE
-- Copyright (c) 2003-2007 OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN, CEDRAT,
--                         EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class WireEdgeSet from BOPAlgo 

	---Purpose: 

uses
    Face   from TopoDS, 
    Shape  from TopoDS, 
    ListOfShape from BOPCol,
    BaseAllocator from BOPCol 
    
--raises

is 
    Create   
    	returns WireEdgeSet from BOPAlgo;  
    ---C++: inline  
    ---C++: alias " virtual ~BOPAlgo_WireEdgeSet();"  
     
    Create (theAllocator: BaseAllocator from BOPCol)   
    	returns WireEdgeSet from BOPAlgo;   
    ---C++: inline  
     
    Clear(me:out);
    ---C++: inline   
 
    SetFace(me:out; 
    	    aF:Face from TopoDS); 
    ---C++: inline        
    
    Face(me) 
	 returns Face from TopoDS; 
    ---C++: return const &  
    ---C++: inline    
    
    AddStartElement(me:out; 
    	    sS: Shape from TopoDS);  
    ---C++: inline       
    
    StartElements(me)  
    	returns ListOfShape from BOPCol;
    ---C++: return const & 
    ---C++: inline   
    
    AddShape(me:out; 
    	    sS:Shape from TopoDS); 
    ---C++: inline        
    
    Shapes(me)  
    	returns ListOfShape from BOPCol;
    ---C++: return const & 
    ---C++: inline   
    
fields
    myFace         : Face from TopoDS is protected; 
    myStartShapes  : ListOfShape from BOPCol is protected;
    myShapes       : ListOfShape from BOPCol is protected;  

end WireEdgeSet;
