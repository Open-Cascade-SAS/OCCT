-- Created on: 1993-01-07
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

generic class MapHasher from TCollection (Key as any)

	---Purpose: A hasher on the keys of a map instantiated from the
    	-- Collections component.
    	-- A hasher provides two functions:
    	-- -   The hashing function (HashCode) transforms a key
    	--   into a bucket index in the map. The number of values
    	--   that can be computed by the hashing function is equal
    	--   to the number of buckets in the map.
    	-- -   IsEqual is the equality test between two keys.
    	--   Hashers are used as parameters in generic maps
    	-- provided by the Collections component.
    	-- MapHasher is a generic class which depends on the type
    	-- of keys, provided that Key is a type from the Standard
    	-- package. In such cases MapHasher may be directly
    	-- instantiated with Key. Note that the package TColStd
    	-- provides some of these instantiations.
    	-- But if Key is not a type from the Standard package you
    	-- must consider MapHasher as a template and build a class
    	-- which includes its functions, in order to use it as a hasher
    	-- in a map instantiated from the Collections component.
    	-- Note that TCollection_AsciiString and
    	-- TCollection_ExtendedString classes correspond to
    	-- these specifications, in consequence they may be used as
    	-- hashers: when Key is one of these two types you may just
    	-- define the hasher as the same type at the time of
    	-- instantiation of your map.

is
    HashCode(myclass; K : Key; Upper : Integer) returns Integer;
	---Level: Public
	---Purpose: Returns a HasCode value  for  the  Key <K>  in the
	-- range 0..Upper.
	-- Default ::HashCode(K,Upper)
	
    IsEqual(myclass; K1, K2 : Key) returns Boolean;
	---Level: Public
	---Purpose: Returns True  when the two  keys are the same. Two
	-- same  keys  must   have  the  same  hashcode,  the
	-- contrary is not necessary.
	-- Default K1 == K2
	
end MapHasher;
