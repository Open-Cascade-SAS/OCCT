-- File:        ClosedShell.cdl
-- Created:     Mon Dec  4 12:02:24 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWClosedShell from RWStepShape

	---Purpose : Read & Write Module for ClosedShell

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     ClosedShell from StepShape,
     EntityIterator from Interface

is

	Create returns RWClosedShell;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable ClosedShell from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : ClosedShell from StepShape);

	Share(me; ent : ClosedShell from StepShape; iter : in out EntityIterator);

end RWClosedShell;
