-- Created on: 1999-03-10
-- Created by: data exchange team
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class AppliedDocumentReference from StepAP214 inherits DocumentReference from StepBasic
 

	
uses
     Document from StepBasic,
     HAsciiString from TCollection,
     DocumentReferenceItem from StepAP214,
     HArray1OfDocumentReferenceItem from StepAP214
	
is
    
    Create returns AppliedDocumentReference;

    Init (me : mutable;
           aAssignedDocument : Document;
           aSource : HAsciiString;
    	   aItems  : HArray1OfDocumentReferenceItem);

    Items (me) returns HArray1OfDocumentReferenceItem ;
    SetItems (me : mutable; aItems : HArray1OfDocumentReferenceItem);
    ItemsValue (me; num : Integer) returns DocumentReferenceItem;
    NbItems (me) returns Integer;

    	
fields
    
    items : HArray1OfDocumentReferenceItem;

end AppliedDocumentReference;
