-- Created on: 1993-03-09
-- Created by: Jean-Louis Frenkel
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


generic class HLRShapeTool from Prs3d ( Shape as any ; Curve as any)
uses
    Projector from HLRAlgo
is
    Create (TheShape: Shape; TheProjector: Projector from HLRAlgo) 
    	    returns HLRShapeTool from Prs3d;
    NbEdges(me) returns Integer from Standard;
    InitVisible(me; EdgeNumber: Integer from Standard);
    MoreVisible(me) returns Boolean from Standard;
    NextVisible(me);
    Visible(me; TheCurve: out Curve; U1,U2: out Real from Standard);
    InitHidden(me; EdgeNumber: Integer from Standard);
    MoreHidden(me) returns Boolean from Standard;
    NextHidden(me);
    Hidden(me; TheCurve: out Curve; U1,U2: out Real from Standard);
    
end HLRShapeTool from Prs3d;
