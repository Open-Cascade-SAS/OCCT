-- Created on: 2001-11-26
-- Created by: Sergey ZARITCHNY
-- Copyright (c) 2001-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

class Gluing from QANewBRepNaming inherits TopNaming from QANewBRepNaming

	---Purpose: Loads a result of Gluing operation in  Data Framework

uses

     Glue      from QANewModTopOpe,
     Shape     from TopoDS, 
     ShapeEnum from  TopAbs,
     Label     from TDF,
     LabelMap  from TDF,
     IndexedDataMapOfShapeListOfShape from TopTools,
     DataMapOfShapeInteger from TopTools

     
raises  NullObject from Standard 

is

    Create returns Gluing from QANewBRepNaming; 
 
    Create(theResultLabel : Label from TDF) 
    returns Gluing from QANewBRepNaming;

    Init(me : in out; theResultLabel : Label from TDF);


    Load (me : in out; theMkGluing : in out Glue from QANewModTopOpe);
      ---Purpose: Loads a Gluing in a data framework  
     
    ---Category: Protected methods
    --           ====================
 
    ShapeType(me; theShape : Shape from TopoDS) 
    ---Purpose: If the shape is a compound the method  
    --          returns the underlying shape type.
    returns ShapeEnum from TopAbs 
    is private; 
     
    GetShape(me; theShape : Shape from TopoDS) 
    ---Purpose: If the shape is a compound the method  
    --          returns the underlying shape.
    returns Shape from TopoDS
    is  private;  
     
    LoadModifiedShapes(me; theMakeShape : in out Glue from QANewModTopOpe)
    ---Purpose: A default implementation for naming of modified shapes of the operation
    is  private; 

    LoadDeletedShapes(me; theMakeShape : in out Glue from QANewModTopOpe)
    ---Purpose: A default implementation for naming of modified shapes of the operation
    is  private; 
     
    Content (me)
    	---Purpose : 
    returns Label from TDF; 
        
    LoadContent(me; theMakeShape : in out Glue from QANewModTopOpe)
    ---Purpose: Loads the content of the result.
    is private;  
     
    LoadResult(me; theMakeShape : in out Glue from QANewModTopOpe) 
    ---Purpose: Loads the result.
    is private; 
    
    IsResultChanged(me; theMakeShape : in out Glue from QANewModTopOpe)  
     ---Purpose: Returns true if the result is not the same as the object shape.
    returns Boolean from Standard is private ;  
     
    SetContext(me :in out; theObject, theTool : Shape from TopoDS);
    
    SetLog(me: in out; theLog : LabelMap from TDF);
     
    LoadSectionEdges(me; theMakeShape : in out Glue from QANewModTopOpe)
    ---Purpose: Loads the deletion of the degenerated edges.
    is private; 
         
    AddToTheUnique(me: in out; theUnique, theIdentifier : Shape from TopoDS) is private;

    RecomputeUnique(me : in out; theMakeShape : in out Glue from QANewModTopOpe)
    ---Purpose: Reset myShared map - shapes, which are modified by both object and tool.
    is private; 

    LoadSourceShapes(me; theSources : in out DataMapOfShapeInteger from TopTools)
    is private;

    LoadUniqueShapes(me: in out; theMakeShape : in out Glue from QANewModTopOpe;
                                 theSources : DataMapOfShapeInteger from TopTools)
    ---Purpose: A default implementation for naming of generated  shapes of the operation
    is  private; 
     
    
fields

    myUnique  : IndexedDataMapOfShapeListOfShape from TopTools;

    myContext : Shape from TopoDS;
    myLog : LabelMap from TDF;

end Gluing;
