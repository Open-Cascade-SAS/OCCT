-- Created on: 1993-01-26
-- Created by: Jean-Louis FRENKEL
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ToolRFace from StdPrs 

	---Purpose: 
uses 
    Curve        from Geom2dAdaptor,
    Face         from TopoDS,
    HSurface     from BRepAdaptor,
    Curve2dPtr   from Adaptor2d,
    Orientation  from TopAbs,
    Explorer     from TopExp

is
    Create returns ToolRFace from StdPrs;    

    Create ( aSurface :HSurface from BRepAdaptor ) 
    returns ToolRFace from StdPrs;

    IsOriented (me) returns Boolean from Standard;

    Init(me: in out); 


    More(me) returns Boolean from Standard;

    Next(me: in out);

    Value(me) returns Curve2dPtr from Adaptor2d;

    Orientation(me) returns Orientation from TopAbs;    

fields
    myFace      : Face       from TopoDS;
    myExplorer  : Explorer   from TopExp;
    DummyCurve  : Curve      from Geom2dAdaptor;
    
end ToolRFace;


