-- Created on: 1994-06-01
-- Created by: Christian CAILLET
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class UpdateLastChange  from IGESSelect  inherits ModelModifier from IGESSelect

    ---Purpose : Allows to Change the Last Change Date indication in the Header
    --           (Global Section) of IGES File. It is taken from the operating
    --           system (time of application of the Modifier).
    --           The Selection of the Modifier is not used : it simply acts as
    --           a criterium to select IGES Files to touch up.
    --           Remark : IGES Models noted as version before IGES 5.1 are in
    --           addition changed to 5.1

uses AsciiString from TCollection,
     IGESModel, CopyTool, ContextModif

is

    Create returns UpdateLastChange;
    ---Purpose : Creates an UpdateLastChange, which uses the system Date

    Performing (me; ctx : in out ContextModif;
    	        target  : IGESModel;
                TC      : in out CopyTool);
    ---Purpose : Specific action : only <target> is used : the system Date
    --           is set to Global Section Item n0 25. Also sets IGES Version
    --           (Item n0 23) to IGES5 if it was older.

    Label (me) returns AsciiString from TCollection;
    ---Purpose : Returns a text which is
    --           "Update IGES Header Last Change Date"

end UpdateLastChange;
