-- Created on: 1994-12-12
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Copy from BRepBuilderAPI inherits ModifyShape from BRepBuilderAPI

	---Purpose: Duplication of a shape.
    	-- A Copy object provides a framework for:
    	-- -   defining the construction of a duplicate shape,
    	-- -   implementing the construction algorithm, and
    	-- -   consulting the result.
        
uses
    Shape             from TopoDS,
    Face              from TopoDS,
    ShapeModification from BRepBuilderAPI,
    ListOfShape       from TopTools


is

    Create
	---Purpose: Constructs an empty copy framework. Use the function
    	-- Perform to copy shapes.
       	returns Copy from BRepBuilderAPI;


    Create(S: Shape from TopoDS; copyGeom: Boolean = Standard_True)
	---Purpose: Constructs a copy framework and copies the shape S.
    	-- Use the function Shape to access the result.
    	-- If copyGeom is False, only topological objects will be copied, while 
    	-- geometry will be shared with original shape.
    	-- Note: the constructed framework can be reused to copy
    	-- other shapes: just specify them with the function Perform.
    	returns Copy from BRepBuilderAPI;


    Perform(me: in out; S: Shape from TopoDS; copyGeom: Boolean = Standard_True)
	---Purpose: Copies the shape S.
    	-- Use the function Shape to access the result.
    	-- If copyGeom is False, only topological objects will be copied, while 
    	-- geometry will be shared with original shape.
    	is static;


end Copy;
