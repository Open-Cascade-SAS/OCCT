-- File:	RWStepFEA_RWCurveElementIntervalConstant.cdl
-- Created:	Thu Dec 12 17:51:04 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWCurveElementIntervalConstant from RWStepFEA

    ---Purpose: Read & Write tool for CurveElementIntervalConstant

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    CurveElementIntervalConstant from StepFEA

is
    Create returns RWCurveElementIntervalConstant from RWStepFEA;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : CurveElementIntervalConstant from StepFEA);
	---Purpose: Reads CurveElementIntervalConstant

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: CurveElementIntervalConstant from StepFEA);
	---Purpose: Writes CurveElementIntervalConstant

    Share (me; ent : CurveElementIntervalConstant from StepFEA;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWCurveElementIntervalConstant;
