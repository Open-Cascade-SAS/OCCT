-- Created on: 1997-11-21
-- Created by: Mister rmi
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package UTL
uses Resource, TCollection,Storage, OSD
is

    xgetenv(aCString: CString from Standard)
    returns ExtendedString from TCollection;
    
    OpenFile(aFile: in out BaseDriver from Storage; aName: ExtendedString from TCollection; aMode : OpenMode from Storage)
    returns Error from Storage;
    
    AddToUserInfo(aData: mutable Data from Storage; anInfo: ExtendedString from TCollection);
    
    Path(aFileName: ExtendedString from TCollection) returns Path from OSD;

    Disk(aPath: Path from OSD) returns ExtendedString from TCollection;
    Trek(aPath: Path from OSD) returns ExtendedString from TCollection;
    Name(aPath: Path from OSD) returns ExtendedString from TCollection;
    Extension(aPath: Path from OSD) returns ExtendedString from TCollection;

    FileIterator(aPath: Path from OSD; aMask:ExtendedString from TCollection) returns FileIterator from OSD;
   
    Extension(aFileName: ExtendedString from TCollection) returns ExtendedString from TCollection;
    
    LocalHost returns ExtendedString from TCollection;
    
    ExtendedString(anAsciiString: AsciiString from TCollection) 
    returns ExtendedString from TCollection;


    GUID(anXString: ExtendedString from TCollection)
    returns GUID from Standard;

    Find(aResourceManager: Manager from Resource; aResourceName: ExtendedString from TCollection)
    returns Boolean from Standard;
    
    Value(aResourceManager: Manager from Resource; aResourceName: ExtendedString from TCollection)
    returns ExtendedString from TCollection;
    

    IntegerValue(anExtendedString: ExtendedString from TCollection)
    returns Integer from Standard;
    
    CString(anExtendedString: ExtendedString from TCollection)
    returns CString from Standard;

    IsReadOnly(aFileName: ExtendedString from TCollection)
    returns Boolean from Standard;
    
end UTL;
