-- Created on: 1994-02-07
-- Created by: Modelistation
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Inter from BRepIntCurveSurface 

	---Purpose: Computes the intersection between a face and a
	--          curve. To intersect one curve with shape method
	--          Init(Shape, curve, tTol) should be used.  To
	--          intersect a few curves with specified shape it is
	--          necessary to load shape one time using method
	--          Load(shape, tol) and find intersection points for
	--          each curve using method Init(curve).  For
	--          iteration by intersection points method More() and
	--          Next() should be used.  
	--          
	--- Example:
	---  Inter.Load(shape, tol); 
	---  for( i =1; i <= nbCurves;i++) 
	---   { 
	---    Inter.Init(curve); 
	---    for(  ;Inter.More(); Inter.Next()) 
	---    {
	---     .......
	---    }
	---   }

uses  
--modified by NIZNHY-PKV Sun Dec 15 16:52:33 2002  f 
     TopolTool  from  BRepTopAdaptor, 
     HSurface  from BRepAdaptor, 
--modified by NIZNHY-PKV Sun Dec 15 16:52:34 2002  t
     Shape               from TopoDS,
     FaceClassifier      from BRepClass,
     State               from TopAbs,
     Explorer            from TopExp,
     IntersectionPoint   from IntCurveSurface,
     HInter              from IntCurveSurface,
     Curve               from GeomAdaptor,
     Lin                 from gp,
     Pnt                 from gp,
     TransitionOnCurve   from IntCurveSurface,
     Face                from TopoDS,
     Box                 from Bnd,
     SequenceOfShape     from TopTools,
     HArray1OfBox        from Bnd,
     HCurve               from GeomAdaptor
    
     
raises 
    NotDone from StdFail	  


is

    Create   returns Inter from BRepIntCurveSurface;
    	--- Purpose: Empty constructor;
    	
    Init(me : in out;
    	 theShape : Shape from TopoDS;
	     theCurve : Curve from GeomAdaptor;
	     theTol: Real  from Standard);
	    
	--- Purpose: Load the Shape, the curve  and initialize the
	--           tolerance used for the classification.
    	
    
    Init(me : in out;
    	 theShape : Shape from TopoDS;
	     theLine  : Lin   from gp;
	     theTol: Real  from Standard);
	    
	--- Purpose: Load the Shape, the curve  and initialize the
	--           tolerance used for the classification.
    	

    Load(me : in out; theShape : Shape from TopoDS; theTol: Real  from Standard);
    --- Purpose: Load the Shape,   and initialize the
	  --           tolerance used for the classification.

    Init(me : in out; theCurve : Curve from GeomAdaptor);
    --- Purpose: Method to find intersections of specified curve with loaded shape.
	  
    
    More(me) returns Boolean from Standard;
  	--- Purpose: returns True if there is a current face.
    	    
					     
    Next(me: in out);
    	--- Purpose: Sets the next intersection point to check.
	
	
    Find(me: in out) is protected;
    	---Purpose: Internal function
    	

    Point(me) returns IntersectionPoint from IntCurveSurface
  	  ---Purpose: returns the current Intersection point.
    	raises NotDone from StdFail;
     

    Pnt(me) returns Pnt from gp
    	---Purpose: returns the current geometric Point
    	---C++: return const & 
     	raises NotDone from StdFail;
	
	

    U(me) returns Real from Standard
    	---Purpose: returns the U parameter of the current point 
    	--          on the current face.
   	  raises NotDone from StdFail;


    V(me) returns Real from Standard
    	---Purpose: returns the V parameter of the current point 
    	--          on the current face.
     	raises NotDone from StdFail;
	

    W(me) returns Real from Standard
    	---Purpose: returns the  parameter of the current point 
    	--          on the curve.
   	  raises NotDone from StdFail;


    State(me) returns State from TopAbs
	  ---Purpose: returns the current state  (IN or ON)
    	raises NotDone from StdFail;


    Transition(me) returns TransitionOnCurve   from IntCurveSurface
    	---Purpose: returns the transition of the line on the surface (IN or OUT or UNKNOWN)
    	raises NotDone from StdFail;
	
	
    Face(me) returns Face from TopoDS;
    	---Purpose: returns the current face.
      ---C++: return const &
    	
	 FindPoint(me : in out) returns Boolean from Standard is protected;
    ---Purpose: Method chec found intersection point

    Clear(me : in out) is protected;
    ---Purpose: Method to clear fields of class

fields

    myTolerance      : Real              from Standard;
    myCurve          : HCurve             from GeomAdaptor;
       
    myIntcs          : HInter             from IntCurveSurface;
    
    myCurrentindex   : Integer           from Standard;
    myCurrentnbpoints: Integer           from Standard;  
    myFastClass       :  TopolTool  from  BRepTopAdaptor; 
    
    myCurrentstate    :  State  from  TopAbs; 
    myCurrentU        :  Real  from  Standard;
    myCurrentV        :  Real  from  Standard;
    myCurveBox      : Box from Bnd;
    myIndFace       : Integer from Standard;
    myFaces         : SequenceOfShape from TopTools;
    myFaceBoxes     : HArray1OfBox from Bnd;

end Inter from BRepIntCurveSurface;
