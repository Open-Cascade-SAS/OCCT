-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class CoordinatedUniversalTimeOffset from StepBasic 

inherits TShared from MMgt

uses

	Integer from Standard, 
	AheadOrBehind from StepBasic, 
	Boolean from Standard
is

	Create returns mutable CoordinatedUniversalTimeOffset;
	---Purpose: Returns a CoordinatedUniversalTimeOffset

	Init (me : mutable;
	      aHourOffset : Integer from Standard;
	      hasAminuteOffset : Boolean from Standard;
	      aMinuteOffset : Integer from Standard;
	      aSense : AheadOrBehind from StepBasic) is virtual;

	-- Specific Methods for Field Data Access --

	SetHourOffset(me : mutable; aHourOffset : Integer);
	HourOffset (me) returns Integer;
	SetMinuteOffset(me : mutable; aMinuteOffset : Integer);
	UnSetMinuteOffset (me:mutable);
	MinuteOffset (me) returns Integer;
	HasMinuteOffset (me) returns Boolean;
	SetSense(me : mutable; aSense : AheadOrBehind);
	Sense (me) returns AheadOrBehind;

fields

	hourOffset : Integer from Standard;
	minuteOffset : Integer from Standard;   -- OPTIONAL can be NULL
	sense : AheadOrBehind from StepBasic; -- an Enumeration
	hasMinuteOffset : Boolean from Standard;

end CoordinatedUniversalTimeOffset;
