-- Created on: 1994-06-03
-- Created by: Christian CAILLET
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class WorkLibrary  from IGESSelect  inherits WorkLibrary  from IFSelect

    ---Purpose : Performs Read and Write an IGES File with an IGES Model

uses CString, Transient, 
     InterfaceModel, Protocol from Interface, CheckIterator, ContextWrite,
     Messenger from Message,
     Protocol from IGESData

is

    Create (modefnes : Boolean = Standard_False)
    	returns mutable WorkLibrary from IGESSelect;
    ---Purpose : Creates a IGES WorkLibrary
    --           If <modefnes> is given as True, it will work for FNES

    ReadFile (me; name : CString;
    	      model    : out mutable InterfaceModel;
    	      protocol : Protocol from Interface)
    	  returns Integer;
    ---Purpose : Reads a IGES File and returns a IGES Model (into <mod>),
    --           or lets <mod> "Null" in case of Error
    --           Returns 0 if OK, 1 if Read Error, -1 if File not opened

    WriteFile (me; ctx : in out ContextWrite)  returns Boolean;
    ---Purpose : Writes a File from a IGES Model (brought by <ctx>)
    --           Returns False (and writes no file) if <ctx> is not for IGES

    DefineProtocol (myclass) returns Protocol from IGESData;
    ---Purpose : Defines a protocol to be adequate for IGES
    --           (encompasses ALL the IGES norm including IGESSolid, IGESAppli)

    DumpEntity (me;
    	       model    : InterfaceModel;
    	       protocol : Protocol from Interface;
	       entity   : Transient;
	       S        : Messenger from Message;
	       level    : Integer);
    ---Purpose : Dumps an IGES Entity with an IGES Dumper. <level> is the one
    --           used by IGESDumper.

fields

    themodefnes : Boolean;

end WorkLibrary;
