-- Created on: 2001-01-06
-- Created by: OCC Team
-- Copyright (c) 2001-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PrinterOStream from Message inherits Printer from Message

    ---Purpose: Implementation of a message printer associated with an ostream
    --          The ostream may be either externally defined one (e.g. cout),
    --          or file stream maintained internally (depending on constructor).

uses

    Address        from Standard,
    OStream        from Standard,
    Gravity        from Message,
    AsciiString    from TCollection,
    ExtendedString from TCollection    

is

    Create (theTraceLevel: Gravity from Message = Message_Info)
    returns PrinterOStream from Message;
    	---Purpose: Empty constructor, defaulting to cout
    
    Create (theFileName: CString; theDoAppend: Boolean;
            theTraceLevel: Gravity from Message = Message_Info)
    returns PrinterOStream from Message;
    	---Purpose: Create printer for output to a specified file.
    	--          The option theDoAppend specifies whether file should be
    	--          appended or rewritten.
    	--          For specific file names (cout, cerr) standard streams are used
    
    Close (me: mutable);
        ---C++: alias ~
    	---Purpose: Flushes the output stream and destroys it if it has been
    	--          specified externally with option doFree (or if it is internal
        --          file stream)

    GetUseUtf8 (me) returns Boolean;
    	---Purpose: Returns option to convert non-Ascii symbols to UTF8 encoding
    	---C++: inline

    SetUseUtf8 (me: mutable; useUtf8: Boolean);
    	---Purpose: Sets option to convert non-Ascii symbols to UTF8 encoding
    	---C++: inline

    GetStream (me) returns OStream;
    	---Purpose: Returns reference to the output stream
	---C++: return &
    	---C++: inline
    
    Send (me; theString : CString; theGravity: Gravity from Message;
	      putEndl: Boolean = Standard_True) is redefined;
    	---Purpose: Puts a message to the current stream
	--          if its gravity is equal or greater
	--          to the trace level set by SetTraceLevel()
	      
    Send (me; theString : AsciiString from TCollection;
              theGravity: Gravity from Message;
	      putEndl: Boolean = Standard_True) is redefined;
    	---Purpose: Puts a message to the current stream
	--          if its gravity is equal or greater
	--          to the trace level set by SetTraceLevel()
	      
    Send (me; theString : ExtendedString from TCollection;
              theGravity: Gravity from Message;
	      putEndl: Boolean = Standard_True) is redefined;
    	---Purpose: Puts a message to the current stream
	--          if its gravity is equal or greater
	--          to the trace level set by SetTraceLevel()
	--          Non-Ascii symbols are converted to UTF-8 if UseUtf8
        --          option is set, else replaced by symbols '?'
	      
fields

    myStream:     Address from Standard; -- pointer to OStream 
    myIsFile:     Boolean from Standard;
    myUseUtf8:    Boolean from Standard;

end PrinterOStream;
