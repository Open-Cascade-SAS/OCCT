-- Created on: 1991-01-23
-- Created by: Christophe MARION
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Datum3D from TopLoc inherits TShared from MMgt

	---Purpose: Describes a coordinate transformation, i.e. a change
-- to an elementary 3D coordinate system, or position in 3D space.
-- A Datum3D is always described relative to the default datum.
-- The default datum is described relative to itself: its
-- origin is (0,0,0), and its axes are (1,0,0) (0,1,0) (0,0,1).

uses
    Trsf   from gp

raises
    ConstructionError from Standard
    
is
    Create returns mutable Datum3D;
    	---Purpose: Constructs a default Datum3D.

    Create(T : Trsf from gp) returns mutable Datum3D from TopLoc
	---Purpose: Constructs a Datum3D form a Trsf from gp. An error is
	--          raised if the Trsf is not a rigid transformation.
    raises 
    	ConstructionError from Standard;
    
    Transformation(me) returns Trsf from gp
    	---Purpose: Returns a gp_Trsf which, when applied to this datum,
    	-- produces the default datum.
    	---C++: inline
    	---C++: return const &
    	is static;
    
    ShallowDump(me; S : in out OStream);
	--- Purpose:
    	-- Writes the contents of this Datum3D to the stream S.
	---C++: function call

fields

    myTrsf : Trsf from gp;

end Datum3D;
