-- Created on: 1999-11-26
-- Created by: Andrey BETENEV
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0

class Certification from StepBasic
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity Certification

uses
    HAsciiString from TCollection,
    CertificationType from StepBasic

is
    Create returns Certification from StepBasic;
	---Purpose: Empty constructor

    Init (me: mutable; aName: HAsciiString from TCollection;
                       aPurpose: HAsciiString from TCollection;
                       aKind: CertificationType from StepBasic);
	---Purpose: Initialize all fields (own and inherited)

    Name (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Name
    SetName (me: mutable; Name: HAsciiString from TCollection);
	---Purpose: Set field Name

    Purpose (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Purpose
    SetPurpose (me: mutable; Purpose: HAsciiString from TCollection);
	---Purpose: Set field Purpose

    Kind (me) returns CertificationType from StepBasic;
	---Purpose: Returns field Kind
    SetKind (me: mutable; Kind: CertificationType from StepBasic);
	---Purpose: Set field Kind

fields
    theName: HAsciiString from TCollection;
    thePurpose: HAsciiString from TCollection;
    theKind: CertificationType from StepBasic;

end Certification;
