-- Created on: 1994-09-29
-- Created by: Dieter THIEMANN
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


package UnitsMethods

uses

    Standard, Geom, Geom2d
    
is

    InitializeFactors(LengthFactor :     Real from Standard;
                      PlaneAngleFactor : Real from Standard;
                      SolidAngleFactor : Real from Standard);

       ---Purpose: Initializes the 3 factors for the conversion of
       --          units

    LengthFactor       
    	returns   Real from Standard;

    PlaneAngleFactor   
    	returns   Real from Standard;

    SolidAngleFactor   
    	returns   Real from Standard;

    Set3dConversion(B : Boolean from Standard);
    
    Convert3d          
    	returns   Boolean from Standard;
    
    RadianToDegree(C : Curve from Geom2d; 
    	    	   S : Surface from Geom)
    	returns Curve from Geom2d;
		   
    DegreeToRadian(C : Curve from Geom2d; 
    	    	   S : Surface from Geom)
    	returns Curve from Geom2d;

    MirrorPCurve(C : Curve from Geom2d)
	returns Curve from Geom2d;

    GetLengthFactorValue (param: Integer) returns Real;
    	---Purpose: Returns value of unit encoded by parameter param
        --          (integer value denoting unit, as described in IGES
        --          standard) in millimeters
	
    GetCasCadeLengthUnit returns Real;
    	---Purpose: Returns value of current internal unit for CASCADE
	--          in millemeters
	
    SetCasCadeLengthUnit (param: Integer);
    	---Purpose: Sets value of current internal unit for CASCADE
	--          by parameter param (integer value denoting unit, 
        --          as described in IGES standard) 
	--          GetCasCadeLengthUnit() will then return value 
	--          equal to GetLengthFactorValue(param)
	
end UnitsMethods;
