-- Created on: 1995-12-08
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class CurveExplorer from TopOpeBRepDS

uses

    DataStructure from TopOpeBRepDS,
    Curve from TopOpeBRepDS
    
is

    Create returns CurveExplorer from TopOpeBRepDS;
    Create(DS : DataStructure from TopOpeBRepDS;
           FindOnlyKeep : Boolean from Standard = Standard_True)
     returns CurveExplorer from TopOpeBRepDS;

    Init(me : in out;
    	 DS : DataStructure from TopOpeBRepDS;
         FindOnlyKeep : Boolean from Standard = Standard_True);

    More(me) returns Boolean  is static;
    Next(me : in out) is static;
    Curve(me) returns Curve from TopOpeBRepDS
    ---C++: return const &
    is static;

    IsCurve(me; I : Integer ) returns Boolean  is static;
    IsCurveKeep(me; I : Integer ) returns Boolean  is static;
    Curve(me; I : Integer ) 
    returns Curve from TopOpeBRepDS
    ---C++: return const &
    is static;
    NbCurve(me : in out) returns Integer
    is static;
 
    Index(me) returns Integer 
    is static;

    Find(me : in out) is static private;
        
fields

    myIndex   : Integer ;
    myMax     : Integer ;
    myDS      : Address ; -- (TopOpeBRepDS_DataStructure*)
    myFound   : Boolean ;
    myFindKeep : Boolean;
    
end CurveExplorer from TopOpeBRepDS;
