-- Created on: 1993-04-07
-- Created by: Laurent BUCHARD
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class IntersectionSegment from IntCurveSurface
 

    ---Purpose: A IntersectionSegment describes a segment of curve 
    --          (w1,w2) where distance(C(w),Surface) is less than a  
    --          given tolerances. 
    
    ---Level: Public

uses

    IntersectionPoint    from IntCurveSurface

is

    Create
    	returns IntersectionSegment from IntCurveSurface;
	
    Create(P1: IntersectionPoint from IntCurveSurface;
    	   P2: IntersectionPoint from IntCurveSurface)
	returns IntersectionSegment from IntCurveSurface;
	
    SetValues(me: in out;
    	     P1: IntersectionPoint from IntCurveSurface;
	     P2: IntersectionPoint from IntCurveSurface)
	 is static;
	 
    Values(me;
    	  P1: out IntersectionPoint from IntCurveSurface;
	  P2: out IntersectionPoint from IntCurveSurface)
	 is static;
	 
    FirstPoint(me;
	       P1: out IntersectionPoint from IntCurveSurface)
	 is static;	 

    SecondPoint(me;
	        P2: out IntersectionPoint from IntCurveSurface)
	 is static;

	 
    FirstPoint(me)
	returns IntersectionPoint from IntCurveSurface 
	---C++: return const &
        is static;	 

    SecondPoint(me)
    	 returns IntersectionPoint from IntCurveSurface
	 ---C++: return const &
	 is static;
 
    Dump(me)
          is static;

fields

    myP1 : IntersectionPoint from IntCurveSurface;
    myP2 : IntersectionPoint from IntCurveSurface;
 
end IntersectionSegment;

