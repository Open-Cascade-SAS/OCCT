-- Created on: 1998-06-03
-- Created by: data exchange team
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class WireVertex from ShapeFix 

    ---Purpose: Fixes vertices in the wire on the basis of pre-analysis
    --          made by ShapeAnalysis_WireVertex (given as argument).
    --          The Wire has formerly been loaded in a ShapeExtend_WireData.

uses 
    Wire from TopoDS,
    WireData from ShapeExtend,
    WireVertex from ShapeAnalysis

is

    Create returns WireVertex from ShapeFix;

    Init (me: in out; wire: Wire from TopoDS; preci: Real);
    	---Purpose: Loads the wire, ininializes internal analyzer
	--          (ShapeAnalysis_WireVertex) with the given precision,
	--          and performs analysis

    Init (me: in out; sbwd: WireData from ShapeExtend; preci: Real);
    	---Purpose: Loads the wire, ininializes internal analyzer
	--          (ShapeAnalysis_WireVertex) with the given precision,
	--          and performs analysis

    Init (me: in out; sawv: WireVertex from ShapeAnalysis);
    	---Purpose: Loads all the data on wire, already analysed by 
	--          ShapeAnalysis_WireVertex

    Analyzer (me) returns WireVertex from ShapeAnalysis;
    	---C++: return const &
    	---Purpose: returns internal analyzer

    WireData (me) returns WireData from ShapeExtend;
    	---C++: return const &
    	---Purpose: returns data on wire (fixed)
	---Remark : calls Analyzer().WireData()

    Wire (me) returns Wire from TopoDS;
    	---Purpose: returns resulting wire (fixed)
	---Remark : calls Analyzer().WireData()->Wire()

    FixSame (me: in out) returns Integer;
    	---Purpose: Fixes "Same" or "Close" status (same vertex may be set,
    	--          without changing parameters)
    	--          Returns the count of fixed vertices, 0 if none

    Fix (me: in out) returns Integer;
    	---Purpose: Fixes all statuses except "Disjoined", i.e. the cases in which a
    	--          common value has been set, with or without changing parameters
    	--          Returns the count of fixed vertices, 0 if none

fields

    myAnalyzer: WireVertex from ShapeAnalysis;

end WireVertex;
