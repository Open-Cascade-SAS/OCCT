-- Created on: 1997-02-04
-- Created by: Alexander BRIVIN
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class PointSet from Vrml 

	---Purpose: defines a PointSet node of VRML specifying geometry shapes.

	--  This node represents a set of points located at the current coordinates. PointSet uses the
        --  current coordinates in order, starting at the index specified by the startIndex field. The
       	--  number of points in the set is specified by the numPoints field. A value of -1 for this field
       	--  indicates that all remaining values in the current coordinates are to be used as points. 
       	--  The points are drawn with the current material and texture. 

	--  Treatment of the current material and normal binding is as follows: PER_PART,
       	--  PER_FACE, and PER_VERTEX bindings bind one material or normal to each point. The
       	--  DEFAULT material binding is equal to OVERALL. The DEFAULT normal binding is
       	--  equal to PER_VERTEX. The startIndex is also used for materials or normals when the
       	--  binding indicates that they should be used per vertex. 
is

    Create ( aStartIndex : Integer from Standard = 0;
    	     aNumPoints  : Integer from Standard = -1 )
        returns PointSet from Vrml;

    SetStartIndex ( me : in out; aStartIndex :  Integer from Standard );
    StartIndex ( me ) returns Integer from Standard;
    
    SetNumPoints ( me : in out; aNumPoints :  Integer from Standard );
    NumPoints ( me )  returns Integer from Standard;

    Print  ( me;  anOStream: in out OStream from Standard) returns OStream from Standard;
    ---C++:  return  & 
    
fields

    myStartIndex : Integer from Standard;   -- Index of 1st coordinate of shape
    myNumPoints  : Integer from Standard;   -- Number of points to draw
    
end PointSet;
