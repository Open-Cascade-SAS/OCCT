-- Created on: 1991-07-23
-- Created by: Christophe MARION
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package Primitives 

	---Purpose: This  package   describes   algorithms  to   build
	--          topological primitives.
	--          
	--          The algorithms  in  this package  are  generic. It
	--          contains :
	--          
	--           *   The Builder  signature   class. Describes the
	--           services    required  from    the  Topology  Data
	--           Structure to build the following primitives.
	--          
	--           * The  OneAxis generic class.  Algorithm  used to
	--           build rotational primitives.
	--               
	--           *  The  Wedge  generic  class. Algorithm to build
	--           boxes and wedges.

uses
    gp        -- gp provides all geometrical information

is


    enumeration Direction is 
	---Purpose: 
    	XMin, XMax, YMin, YMax, ZMin, ZMax
    end Direction;
    
    deferred generic class OneAxis;
    	
    generic class Wedge; 
    
end Primitives;
