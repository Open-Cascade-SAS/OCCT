-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class EdgeLoop from StepShape 

inherits Loop from StepShape 
-- WARNING : Multiple EXPRESS inheritance
-- Not yet automaticly managed
-- inherits Path from StepShape 


-- Hand made changes : All the attributes theoricly inherited from the Path
-- entity are explicitly declared in the EdgeLoop entity.
-- The path is not directly referenced by any other entities. As far as
-- Path supertype, topological representation item, is also a 
-- supertype of Edge, this mapping is equivalent.

uses

    	HAsciiString          from TCollection,
	HArray1OfOrientedEdge from StepShape, 
	OrientedEdge          from StepShape

is

	Create returns mutable EdgeLoop;
	---Purpose: Returns a EdgeLoop

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aEdgeList : mutable HArray1OfOrientedEdge from StepShape);

	-- Specific Methods for Field Data Access --

	SetEdgeList(me : mutable; aEdgeList : mutable HArray1OfOrientedEdge);
	EdgeList (me) returns mutable HArray1OfOrientedEdge;
	EdgeListValue (me; num : Integer) returns mutable OrientedEdge;
	NbEdgeList (me) returns Integer;

fields

	edgeList : HArray1OfOrientedEdge from StepShape;

end EdgeLoop;
