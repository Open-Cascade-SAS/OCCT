-- Created on: 1992-02-11
-- Created by: Christian CAILLET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



package StepData

    ---Purpose : Gives basic data definition for Step Interface.
    --           Any class of a data model described in EXPRESS Language
    --           is candidate to be managed by a Step Interface

uses Standard, MMgt, TCollection, TColStd, Dico, LibCtl, Interface, Message

is

    class StepModel;
    class UndefinedEntity;
    deferred class SelectType;

    enumeration Logical  is LFalse, LTrue, LUnknown;
    ---Purpose : A Standard Definition for STEP (which knows Boolean too)

    class Field;
    class SelectMember;
    	class SelectInt;
	class SelectReal;
	class SelectNamed;
	class SelectArrReal;

    class PDescr;
    class FieldList;    -- basic one (no field)
    	class FieldList1;
	class FieldListN;
	class FieldListD;
    deferred class EDescr;
    	class ESDescr;
	class ECDescr;
    deferred class Described;
    	class Simple;
	class Plex;
    class FreeFormEntity;

    class Protocol;                     -- basic protocol for Step
    deferred class GeneralModule;       -- general services

    deferred class FileRecognizer  instantiates
    	Recognizer from Interface (AsciiString from TCollection, Transient);

    class FileProtocol;
    class HeaderTool;
    class EnumTool;

    class DescrProtocol;
    class DescrGeneral;
    class DescrReadWrite;

    class StepReaderData;               -- litteral description of Step File
    class StepReaderTool;
    deferred class ReadWriteModule;
    class StepWriter;                   -- idem but in the other sense
    class StepDumper;

    class WriterLib instantiates  Library from LibCtl
    	(Transient, ReadWriteModule, Protocol from StepData);

    class DefaultGeneral;     -- Default Module which processes UnknownEntity


    	--   General Routines   --
    	--   HeaderProtocol/AddHeaderProtocol are used to handle Header items :
    	--   Reading/Writing but also Copying,Checking,Dumping
    	--   
    	--   
    	-- Init & Protocol encapsulate the general actions required to work with
    	-- this package. While their use is not mandatory, it makes work easier.

    class  Array1OfField  instantiates    Array1 from TCollection
    	(Field from StepData);
    class HArray1OfField  instantiates   HArray1 from TCollection
    	(Field from StepData,Array1OfField from StepData);

    HeaderProtocol  returns Protocol from StepData;
    ---Purpose : Returns the recorded HeaderProtocol, which can be :
    --           - a Null Handle if no Header Protocol was yet defined
    --           - a simple Protocol if only one was defined
    --           - a FileProtocol if more than one Protocol was yet defined

    AddHeaderProtocol (headerproto : Protocol from StepData);
    ---Purpose : Adds a new Header Protocol to the Header Definition

    Init;
    ---Purpose : Prepares General Data required to work with this package,
    --           which are the Protocol and Modules to be loaded into Libraries

    Protocol  returns Protocol from StepData;
    ---Purpose : Returns a Protocol from StepData (avoids to create it)

end StepData;
