-- Created on: 1998-07-29
-- Created by: Christian CAILLET
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



package STEPEdit

    ---Purpose : Provides tools to exploit and edit a set of STEP data :
    --           editors, selections ..

uses Standard, TCollection,
     Interface, IFSelect, StepData

is

    class EditContext;
    -- This class is for global context : ApplicationContext,
    --   ProductRelatedProductCategory

    class EditSDR;
    -- This class allows to edit product data for a SDR


    	--  Some useful operators
    	--  They are not classes, they are just based on general tools

    Protocol returns Protocol from Interface;
    ---Purpose : Returns a Protocol fit for STEP (creates the first time)

    NewModel returns StepModel from StepData;
    ---Purpose : Returns a new empty StepModel fit for STEP
    --           i.e. with its header determined from Protocol

    SignType returns Signature from IFSelect;
    ---Purpose : Returns a SignType fit for STEP (creates the first time)

    NewSelectSDR returns SelectSignature from IFSelect;
    ---Purpose : Creates a Selection for ShapeDefinitionRepresentation
    --           By default searches among root entities

    NewSelectPlacedItem returns SelectSignature from IFSelect;
    ---Purpose : Creates a Selection for Placed Items, i.e. MappedItem or
    --           ContextDependentShapeRepresentation, which itself refers to a
    --           RepresentationRelationship with possible subtypes (Shape...
    --           and/or ...WithTransformation)
    --           By default in the whole StepModel

    NewSelectShapeRepr returns SelectSignature from IFSelect;
    ---Purpose : Creates a Selection for ShapeRepresentation and its sub-types,
    --           plus ContextDependentShapeRepresentation (which is not a
    --           sub-type of ShapeRepresentation)
    --           By default in the whole StepModel

end STEPEdit;
