-- Created on: 1991-09-18
-- Created by: Didier PIFFAULT
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

generic class ToolPolyhedron from Intf (Polyhedron as any)

    ---Purpose: Describes the signature  of  a polyedral surface with  only
    --          triangular facets and the information  necessary to compute
    --          the interferences.


uses    XYZ from gp,
    	Pnt from gp,
    	Box from Bnd,
	HArray1OfBox from Bnd


raises  OutOfRange from Standard


is  Bounding       (myclass; thePolyh : Polyhedron)
    	    	    returns Box from Bnd;
    ---Purpose: Returns the bounding box of the ToolPolyhedron.

    ComponentsBounding
       	    	   (myclass; thePolyh : Polyhedron)
    	    	    returns HArray1OfBox from Bnd;
    ---Purpose: Returns the array of boxes. The box <n> corresponding 
    --          to the triangle <n>.


    DeflectionOverEstimation
		   (myclass; thePolyh : Polyhedron)
    	    	    returns Real from Standard;
    ---Purpose: Returns the tolerance of the polygon.


-- Structure needings :

    NbTriangles	   (myclass; thePolyh : Polyhedron) 
    	    	    returns Integer from Standard;
    ---Purpose: Returns the number of triangles in this polyedron.


    Triangle	   (myclass; thePolyh : Polyhedron;
		    Index     : in Integer from Standard;
		    P1,P2,P3  : out Integer from Standard)
		    raises OutOfRange from Standard;
    ---Purpose: Returns the indices  of  the 3 points of  the triangle of
    --          address Index in the ToolPolyhedron.


    Point	   (myclass; thePolyh : Polyhedron;
		    Index : in Integer)
		    returns Pnt from gp
		    raises OutOfRange from Standard;
    ---Purpose: Returns the point of index i in the polyedron.


    TriConnex	   (myclass; thePolyh : Polyhedron;
		    Triang	 : in Integer;
		    Pivot,Pedge	 : in Integer;
		    TriCon	 : out Integer;
		    OtherPedge	 : out Integer)
		    returns Integer
		    raises OutOfRange from Standard;
    ---Purpose: Returns  the  triangle <Tricon> connected  to  the triangle
    --          <Triang> by  the edge <Pivot><Pedge>.   The  third point of
    --          the connected triangle is returned in <OtherPedge> (Used to
    --          turn  around a vertex).   When the edge  <Pivot><Pedge>  is
    --          free  (no  connected triangle) <Tricon> is  null.   In this
    --          case the function returns the triangle on the free bound of
    --          the polyhedron connected to <Triang> by vertex <Pivot>.



end ToolPolyhedron;
