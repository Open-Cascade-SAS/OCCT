-- Created on: 1999-03-09
-- Created by: data exchange team
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class PersonAndOrganizationItem from StepAP214 inherits ApprovalItem from StepAP214

	-- <PersonAndOrganizationItem> is an EXPRESS Select Type construct translation.
	-- it gathers : ApprovalPersonOrganization, AutoDesignDateAndPersonAssignment

uses

    	AppliedOrganizationAssignment from StepAP214
	
is

	Create returns PersonAndOrganizationItem;
	---Purpose : Returns a PersonAndOrganizationItem SelectType

	CaseNum (me; ent : Transient) returns Integer is redefined;
	---Purpose: Recognizes a APersonAndOrganizationItem Kind Entity that is :
    	--        1 -> AppliedOrganizationAssignment
    	--        2 -> AssemblyComponentUsageSubstitute
	--        3 -> DocumentFile
    	--        4 -> MaterialDesignation
    	--        5 -> MechanicalDesignGeometricPresentationRepresentation
	--        6 -> PresentationArea
    	--        7 -> Product
	--        8 -> ProductDefinition
    	--        9 -> ProductDefinitionFormation
	--    	  10 -> ProductDefinitionRelationship
	--        11 -> PropertyDefinition
    	--        12 -> ShapeRepresentation
    	--        13 -> SecurityClassification
	--        0 else


    	AppliedOrganizationAssignment (me) returns any AppliedOrganizationAssignment;
    	---Purpose : returns Value as a AppliedOrganizationAssignment (Null if another type)

	
end PersonAndOrganizationItem;
