-- Created on: 1993-01-09
-- Created by: CKY / Contract Toubro-Larsen ( SIVA )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class BooleanTree from IGESSolid  inherits IGESEntity

        ---Purpose: defines BooleanTree, Type <180> Form Number <0>
        --          in package IGESSolid
        --          The Boolean tree describes a binary tree structure
        --          composed of regularized Boolean operations and operands,
        --          in post-order notation.

uses

        HArray1OfInteger     from TColStd,
        HArray1OfIGESEntity  from IGESData

raises OutOfRange

is

        Create returns mutable BooleanTree;

        -- Specific Methods pertaining to the class

        Init (me         : mutable;
              operands   : HArray1OfIGESEntity;
              operations : HArray1OfInteger);
        ---Purpose : This method is used to set the fields of the class
        --           BooleanTree
        --       - operands   : Array containing pointer to DE of operands
        --       - operations : Array containing integer type for operations

        Length (me) returns Integer;
        ---Purpose : returns the length of the post-order list

        IsOperand (me; Index: Integer) returns Boolean
        raises OutOfRange;
        ---Purpose : returns True if Index'th value in the post-order list is an Operand;
        -- else returns False if it is an Integer Operations
        -- raises exception if Index < 1 or Index > Length()

        Operand (me; Index : Integer) returns IGESEntity
        raises OutOfRange;
        ---Purpose : returns the Index'th value in the post-order list only if it is 
        -- an operand else returns NULL
        -- raises exception if Index < 1 or Index > Length()

        Operation (me; Index : Integer) returns Integer
        raises OutOfRange;
        ---Purpose : returns the Index'th value in the post-order list only if it is 
        -- an operation else returns 0
        -- raises exception if Index < 1 or Index > Length()

fields

--
-- Class    : IGESSolid_BooleanTree
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class BooleanTree.
--
-- Reminder : A BooleanTree instance is defined by :
--            - a list having operation codes (integers) or pointers to
--            - operands. A positive value in the data entry implies an
--            - operation code; a negative value implies the absolute value
--            - is to be taken as a pointer to an operand.

        theOperands   : HArray1OfIGESEntity;

        theOperations : HArray1OfInteger;

end BooleanTree;
