-- File     : MeshVS_SensitivePolyhedron.cdl
-- Created  : 21 January 2005
-- Author   : Alexander SOLOVYOV
---Copyright: Open CASCADE 2005

class SensitivePolyhedron from MeshVS inherits SensitiveEntity from Select3D

uses
    EntityOwner                from SelectBasics,
    Projector                  from Select3D,
    Location                   from TopLoc,
    Real                       from Standard,
    Boolean                    from Standard,
    Array1OfPnt2d              from TColgp,
    SequenceOfInteger          from TColStd,
    Box2d                      from Bnd,
    Lin                        from gp,
    ListOfBox2d                from SelectBasics,
    Array1OfPnt                from TColgp,
    HArray1OfPnt               from TColgp,
    HArray1OfPnt2d             from TColgp,
    HArray1OfSequenceOfInteger from MeshVS,
    XY                         from gp

is
    Create( Owner : EntityOwner from SelectBasics;
            Nodes : Array1OfPnt from TColgp;
            Topo  : HArray1OfSequenceOfInteger from MeshVS ) returns mutable SensitivePolyhedron from MeshVS;

    Project( me:mutable; aProjector: Projector from Select3D ) is redefined;

    GetConnected( me:mutable; aLocation: Location from TopLoc ) returns SensitiveEntity from Select3D 
       is redefined;
   
    Matches( me   : mutable; 
             X,Y  : Real from Standard;
             aTol : Real from Standard;
             DMin : out Real from Standard ) returns Boolean is redefined;

    Matches( me                  : mutable; 
             XMin,YMin,XMax,YMax : Real from Standard;
             aTol                : Real from Standard ) returns Boolean from Standard is redefined;

    Matches( me       : mutable; 
             Polyline : Array1OfPnt2d from TColgp;
	     aBox     : Box2d from Bnd;
             aTol     : Real from Standard ) returns Boolean from Standard is redefined;

    GetBox2d( me; aBox : out Box2d from Bnd ) is protected;

    FindIntersection( me; NodesIndices : SequenceOfInteger from TColStd;
                          EyeLine      : Lin from gp ) returns Real is protected;

    ComputeDepth( me; EyeLine: Lin from gp ) returns Real from Standard is redefined;

--  ComputeSize( me ) returns Real from Standard is redefined;

    Areas( me: mutable; aResult : in out ListOfBox2d from SelectBasics ) is redefined;

fields
    myNodes   : HArray1OfPnt from TColgp;
    myNodes2d : HArray1OfPnt2d from TColgp;
    myTopo    : HArray1OfSequenceOfInteger from MeshVS;
    myCenter  : XY from gp;

end SensitiveEntity;

