-- Created on: 1993-10-20
-- Created by: Jean-Louis FRENKEL
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PlaneSet from Prs3d inherits TShared from MMgt

uses

    Length from Quantity,
    Pln from gp
is

    Create( Xdir,Ydir,Zdir: Real from Standard;
            Xloc,Yloc,Zloc: Length from Quantity;
    	    anOffset: Length from Quantity)
    returns PlaneSet from Prs3d;

    SetDirection(me: mutable; X,Y,Z: Real from Standard);
    SetLocation(me: mutable; X,Y,Z: Length from Quantity);
    SetOffset(me: mutable; anOffset: Length from Quantity);
    
    Plane(me) returns Pln from gp;
    Offset(me) returns Length from Quantity;
    Location(me; X,Y,Z: out Length from Quantity);
    Direction(me; X,Y,Z: out Length from Quantity);

fields

    myPlane: Pln from gp;
    myOffset: Length from Quantity;
    
end PlaneSet from Prs3d;
