-- File:	BRepBlend_RstRstConstRad.cdl
-- Created:	Thu Feb  6 16:22:22 1997
-- Author:	Jacques GOUSSARD
-- Author:	Laurent BOURESCHE
--		<lbo@pomalox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1997

class RstRstConstRad from BRepBlend
inherits RstRstFunction from Blend

	---Purpose: 

uses Vector          from math,
     Matrix          from math,
     Ax1             from gp,
     Vec             from gp,
     Vec2d           from gp,
     Pnt             from gp,
     Pnt2d           from gp,
     Circ            from gp,
     Array1OfPnt     from TColgp,
     Array1OfVec     from TColgp,
     Array1OfPnt2d   from TColgp,
     Array1OfVec2d   from TColgp,
     Array1OfReal    from TColStd,
     Array1OfInteger from TColStd,
     Shape           from GeomAbs,
     Point           from Blend,
     SectionShape    from BlendFunc,
     HSurface        from Adaptor3d,
     HCurve          from Adaptor3d,
     HCurve2d        from Adaptor2d,
     CurveOnSurface  from Adaptor3d,
     ParameterisationType from Convert,
     DecrochStatus   from Blend

is

    Create(Surf1    : HSurface from Adaptor3d;
           Rst1     : HCurve2d from Adaptor2d;
    	   Surf2    : HSurface from Adaptor3d;
    	   Rst2     : HCurve2d from Adaptor2d; 
    	   CGuide   : HCurve   from Adaptor3d)
    returns RstRstConstRad from BRepBlend;

    NbVariables(me)
    ---Purpose: Returns 2.
    returns Integer from Standard;

    NbEquations(me)
    ---Purpose: Returns 2.
    returns Integer from Standard;

    Value(me: in out; X: Vector; F: out Vector)
    ---Purpose: computes the values <F> of the Functions for the 
    --          variable <X>.
    --          Returns True if the computation was done successfully, 
    --          False otherwise.
    returns Boolean from Standard;
    
    Derivatives(me: in out; X: Vector; D: out Matrix)
    ---Purpose: returns the values <D> of the derivatives for the 
    --          variable <X>.
    --          Returns True if the computation was done successfully, 
    --          False otherwise.
    returns Boolean from Standard;
    
    Values(me: in out; X: Vector; F: out Vector; D: out Matrix)
    ---Purpose: returns the values <F> of the functions and the derivatives
    --          <D> for the variable <X>.
    --          Returns True if the computation was done successfully, 
    --          False otherwise.
    returns Boolean from Standard;

    Set(me      : in out; 
        SurfRef1 : HSurface from Adaptor3d;
    	RstRef1  : HCurve2d from Adaptor2d;
        SurfRef2 : HSurface from Adaptor3d;
    	RstRef2  : HCurve2d from Adaptor2d);
    	   
    Set(me: in out; Param: Real from Standard);

    Set(me: in out; First, Last: Real from Standard);
    ---Purpose: Sets the bounds of the parametric interval on 
    --          the guide line.
    --          This determines the derivatives in these values if the
    --          function is not Cn.

    GetTolerance(me; Tolerance: out Vector from math; Tol: Real from Standard);

    GetBounds(me; InfBound,SupBound: out Vector from math);

    IsSolution(me: in out; Sol: Vector from math; Tol: Real from Standard)
    returns Boolean from Standard;

     GetMinimalDistance(me) 
        ---Purpose: Returns   the    minimal  Distance  beetween   two
        --          extremitys of calculed sections.          
   	returns  Real  from  Standard 
	is redefined;

--- TheFollowing methods are called only when 
--  IsSolution returns Standard_True.

    PointOnRst1(me)
    ---C++: return const&
    returns Pnt from gp;

    PointOnRst2(me)
    ---C++: return const&
    returns Pnt from gp;

    Pnt2dOnRst1(me)
    ---Purpose: Returns U,V coordinates of the point on the surface.
    ---C++: return const&
    returns Pnt2d from gp;

    Pnt2dOnRst2(me)
    ---Purpose: Returns  U,V coordinates of the point  on the curve on
    --          surface.
    ---C++: return const&
    returns Pnt2d from gp;

    ParameterOnRst1(me)
    ---Purpose: Returns parameter of the point on the curve.
    returns Real from Standard;

    ParameterOnRst2(me)
    ---Purpose: Returns parameter of the point on the curve.
    returns Real from Standard;

    IsTangencyPoint(me)
    returns Boolean from Standard;

    TangentOnRst1(me)
    ---C++: return const&
    returns Vec from gp;

    Tangent2dOnRst1(me)
    ---C++: return const&
    returns Vec2d from gp;

    TangentOnRst2(me)
    ---C++: return const&
    returns Vec from gp;

    Tangent2dOnRst2(me)
    ---C++: return const&
    returns Vec2d from gp;

    Decroch(me; 
    	    Sol    : Vector from math;
	    NRst1, TgRst1 : out Vec from gp;
    	    NRst2, TgRst2 : out Vec from gp)
    ---Warning: Peut  etre  appele sans appel prealable   a issolution
    --          mais les valeurs  calculees risquent  de ne pas  avoir
    --          grand  sens.    
    ---Purpose: Permet  d ' implementer   un   critere  de  decrochage
    --          specifique a la fonction.
    returns DecrochStatus from Blend
    is static;

-- methodes hors template (en plus du create)

    Set(me     : in out; 
    	Radius : Real from Standard; 
    	Choix  : Integer from Standard)
    is static;

    Set(me: in out; TypeSection: SectionShape from BlendFunc)
    ---Purpose: Sets  the  type  of   section generation   for the
    --          approximations. 
    is static;

    CenterCircleRst1Rst2(me;
                  	 PtRst1 : Pnt      from gp;
                    	 PtRst2 : Pnt      from gp;
		         np     : Vec      from gp;
		         Center : out Pnt  from gp;
		         VdMed  : out Vec  from gp)		   
    ---Purpose: Give the center of circle define by PtRst1, PtRst2 and
    --          radius ray.
    returns Boolean from Standard         
    is static;		   
		   
    Section(me        : in out; 
            Param     : Real from Standard;
            U,V       : Real from Standard;
            Pdeb,Pfin : out Real from Standard;
            C         : out Circ from gp)
    is static;

-- Methods for the approximation
-- 
    IsRational(me) returns Boolean
    ---Purpose: Returns  if the section is rationnal
    is static;

    GetSectionSize(me) returns Real
    ---Purpose:  Returns the length of the maximum section
    is static;
    
    GetMinimalWeight(me; Weigths  : out Array1OfReal  from TColStd)
    ---Purpose: Compute the minimal value of weight for each poles
    --          of all sections.
    is static;

    NbIntervals(me; S : Shape from GeomAbs) returns Integer
    ---Purpose: Returns  the number  of  intervals for  continuity
    --          <S>. May be one if Continuity(me) >= <S>
    is static;
    
    Intervals(me; T : in out Array1OfReal from TColStd; 
    	          S : Shape from GeomAbs)
    ---Purpose: Stores in <T> the  parameters bounding the intervals
    --          of continuity <S>.        
    --          The array must provide  enough room to  accomodate
    --          for the parameters. i.e. T.Length() > NbIntervals()
    is static;

    GetShape(me        : in out;
             NbPoles   : out Integer from Standard;
    	     NbKnots   : out Integer from Standard;
             Degree    : out Integer from Standard;
             NbPoles2d : out Integer from Standard)
    is static;

    GetTolerance(me; 
    	    	 BoundTol, SurfTol, AngleTol : Real;
		 Tol3d : out Vector;
		 Tol1D : out Vector )
    ---Purpose: Returns the tolerance to reach in approximation
    --          to respecte
    --          BoundTol error at the Boundary
    --          AngleTol tangent error at the Boundary
    --          SurfTol error inside the surface.
    is static;

    Knots(me: in out; TKnots: out Array1OfReal from TColStd)
    is static;

    Mults(me: in out; TMults: out Array1OfInteger from TColStd)
    is static;

    Section(me       : in out ; 
    	    P        : Point from Blend;
            Poles    : out Array1OfPnt   from TColgp;
	    DPoles   : out Array1OfVec   from TColgp;
  	    Poles2d  : out Array1OfPnt2d from TColgp;
	    DPoles2d : out Array1OfVec2d from TColgp;
	    Weigths  : out Array1OfReal  from TColStd;
	    DWeigths : out Array1OfReal  from TColStd)
    ---Purpose: Used for the first and last section 
    returns Boolean from Standard
    is static;

    Section(me       : in out ; 
    	    P        : Point from Blend;
            Poles    : out Array1OfPnt   from TColgp;
    	    Poles2d  : out Array1OfPnt2d from TColgp;
	    Weigths  : out Array1OfReal  from TColStd)
    is static;


    Section(me: in out; P: Point from Blend;
			Poles     : out Array1OfPnt   from TColgp;
			DPoles    : out Array1OfVec   from TColgp;
			D2Poles   : out Array1OfVec   from TColgp;
    	                Poles2d   : out Array1OfPnt2d from TColgp;
			DPoles2d  : out Array1OfVec2d from TColgp;
			D2Poles2d : out Array1OfVec2d from TColgp;
			Weigths   : out Array1OfReal  from TColStd;
			DWeigths  : out Array1OfReal  from TColStd;
                        D2Weigths : out Array1OfReal  from TColStd)
    ---Purpose: Used for the first and last section
    --          The method returns Standard_True if the derivatives
    --          are computed, otherwise it returns Standard_False.
    returns Boolean from Standard
    is static;

    Resolution(me; 
    	       IC2d : Integer from Standard;
	       Tol  : Real from Standard;
	       TolU, TolV : out Real from Standard);

fields

    surf1    : HSurface             from Adaptor3d;
    surf2    : HSurface             from Adaptor3d;
    rst1     : HCurve2d             from Adaptor2d;
    rst2     : HCurve2d             from Adaptor2d;    
    cons1    : CurveOnSurface       from Adaptor3d;
    cons2    : CurveOnSurface       from Adaptor3d;    
    guide    : HCurve               from Adaptor3d; 
    tguide   : HCurve               from Adaptor3d; 
    ptrst1   : Pnt                  from gp;
    ptrst2   : Pnt                  from gp;
    pt2drst1 : Pnt2d                from gp;
    pt2drst2 : Pnt2d                from gp;
    prmrst1  : Real                 from Standard;
    prmrst2  : Real                 from Standard;    
    istangent: Boolean              from Standard;
    tgrst1   : Vec                  from gp;
    tg2drst1 : Vec2d                from gp;
    tgrst2   : Vec                  from gp;
    tg2drst2 : Vec2d                from gp;

    ray      : Real                 from Standard;
    choix    : Integer              from Standard;
    ptgui    : Pnt                  from gp;
    d1gui    : Vec                  from gp;
    d2gui    : Vec                  from gp;
    nplan    : Vec                  from gp;
    normtg   : Real                 from Standard;
    theD     : Real                 from Standard;
       
    surfref1 : HSurface             from Adaptor3d;
    rstref1  : HCurve2d             from Adaptor2d;
    surfref2 : HSurface             from Adaptor3d;
    rstref2  : HCurve2d             from Adaptor2d;
    maxang   : Real                 from Standard;
    minang   : Real                 from Standard;   
    distmin  : Real                 from Standard;   
    mySShape : SectionShape         from BlendFunc;
    myTConv  : ParameterisationType from Convert;

end RstRstConstRad;









