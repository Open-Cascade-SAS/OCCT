-- Created on: 1996-01-25
-- Created by: Frederic MAUPAS
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MakeRectangularTrimmedSurface from GeomToStep  
    inherits Root from GeomToStep
    
    ---Purpose: This class implements the mapping between class
    --          RectangularTrimmedSurface from Geom and the class
    --          RectangularTrimmedSurface from  
    --          StepGeom which describes a 
    --          rectangular_trimmed_surface from ISO-IS 10303-42
  
uses RectangularTrimmedSurface from Geom,
     RectangularTrimmedSurface from StepGeom
     
raises NotDone from StdFail
     
is 

Create ( RTSurf : RectangularTrimmedSurface from Geom ) returns
    MakeRectangularTrimmedSurface;

Value (me) returns
    RectangularTrimmedSurface from StepGeom
    raises NotDone
    is static;
    ---C++: return const&

fields

    theRectangularTrimmedSurface :
    	RectangularTrimmedSurface from StepGeom;
    	-- The solution from StepGeom
    	
end MakeRectangularTrimmedSurface;


