-- Created on: 1995-11-02
-- Created by: Jing Cheng MEI
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class FindPlane from BRepBuilderAPI

	---Purpose: Describes functions to find the plane in which the edges
    	-- of a given shape are located.
    	-- A FindPlane object provides a framework for:
    	-- -   extracting the edges of a given shape,
    	-- -   implementing the construction algorithm, and
    	-- -   consulting the result.
        
uses
    
    Shape    from TopoDS,
    Plane    from Geom

raises

    NoSuchObject from Standard

is

    Create 
    returns FindPlane from BRepBuilderAPI;
    	---Purpose: Initializes an empty algorithm. The function Init is then used to define the shape. 
    
    Create (S         : Shape   from TopoDS; 
    	    Tol       : Real    from Standard = -1)
    returns FindPlane from BRepBuilderAPI;
	---Purpose:  Constructs the plane containing the edges of the shape S.
    	-- A plane is built only if all the edges are within a distance
    	-- of less than or equal to tolerance from a planar surface.
    	-- This tolerance value is equal to the larger of the following two values:
    	-- -   Tol, where the default value is negative, or
    	-- -   the largest of the tolerance values assigned to the individual edges of S.
    	--   Use the function Found to verify that a plane is built.
    	-- The resulting plane is then retrieved using the function Plane.

    Init (me : in out; 
          S         : Shape   from TopoDS; 
    	  Tol       : Real    from Standard = -1);
	---Purpose: Constructs the plane containing the edges of the shape S.
    	-- A plane is built only if all the edges are within a distance
    	-- of less than or equal to tolerance from a planar surface.
    	-- This tolerance value is equal to the larger of the following two values:
    	-- -   Tol, where the default value is negative, or
    	-- -   the largest of the tolerance values assigned to the individual edges of S.
    	--   Use the function Found to verify that a plane is built.
    	-- The resulting plane is then retrieved using the function Plane.
    
    Found(me)
    returns Boolean from Standard;
    	---Purpose: Returns true if a plane containing the edges of the
    	-- shape is found and built. Use the function Plane to consult the result.   
    Plane(me)
    returns mutable Plane from Geom;
    	---Purpose: Returns the plane containing the edges of the shape.
    	-- Warning
    	-- Use the function Found to verify that the plane is built. If
    	-- a plane is not found, Plane returns a null handle.   
        
fields

    myPlane     : Plane from Geom;

end FindPlane;
