-- Created on: 1992-10-19
-- Created by: Laurent BUCHARD
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

generic class IntPolyPolyGen from IntCurve (
    TheCurve       as any;
    TheCurveTool   as any; -- as CurveTool from IntCurve (TheCurve)
    TheProjPCur    as any) -- as ProjPCurGen from IntCurve
    
inherits Intersection from IntRes2d



    ---Level: Internal

uses Domain       from IntRes2d  


    class ThePolygon2d instantiates Polygon2dGen from IntCurve
    	    	    	    	   (TheCurve,
                                    TheCurveTool);
				    
    class TheDistBetweenPCurves instantiates DistBetweenPCurvesGen
    	                           (TheCurve,
                                    TheCurveTool);

    class  ExactIntersectionPoint 

    	uses  Vector        from  math , 
	      ThePolygon2d  from  IntCurve  
    	is  
    	    Create  ( C1  :  TheCurve; 
	    	      C2  :  TheCurve;  
    	    	      Tol :   Real  from  Standard ) 
		returns  ExactIntersectionPoint from  IntCurve    ; 
    	    
    	    Perform ( me: in out ;
    	    	      Poly1       :  ThePolygon2d  from  IntCurve  ; 
	    	      Poly2       :  ThePolygon2d  from  IntCurve  ;  
		      NumSegOn1   :  out  Integer  from  Standard  ; 
		      NumSegOn2   :  out  Integer  from  Standard  ; 
		      ParamOnSeg1 :  out  Real     from  Standard  ; 
		      ParamOnSeg2 :  out  Real     from  Standard );

    	    Perform (  me: in out ;
    	    	       Uo  :  Real  from  Standard  ; 
	    	       Vo  :  Real  from  Standard  ; 
		       UInf  :  Real  from  Standard  ; 
		       VInf  :  Real  from  Standard  ;  
		       USup  :  Real  from  Standard  ;   
		       VSup  :  Real  from  Standard  );
		       
    	    NbRoots  ( me )  
    	    	returns  Integer  from  Standard  ;

    	    Roots  (  me  : in out ; 
    	    	      U   : out  Real from  Standard  ; 
    	    	      V   : out  Real from  Standard  ) ;
    	
	    MathPerform  ( me : in out )  is  private ; 
	    
    	    AnErrorOccurred  (  me  ) 
	     	returns  Boolean                from  Standard  ;
	    	
    	    fields 
	     
	    	done             :  Boolean                from  Standard  ; 
		nbroots          :  Integer                from  Standard  ;  
		myTol            :  Real                   from  Standard  ;  
		FctDist          :  TheDistBetweenPCurves  from  IntCurve  ; 
		ToleranceVector  :  Vector                 from  math  ; 
		BInfVector       :  Vector                 from  math  ;  
		BSupVector       :  Vector                 from  math  ; 
		StartingPoint    :  Vector                 from  math  ;  
		Root             :  Vector                 from  math  ;  
    	        anErrorOccurred  :  Boolean                from  Standard  ;
	     end ExactIntersectionPoint from  IntCurve; 	


is

    Create  
	returns IntPolyPolyGen from IntCurve;
    
    
    Perform(me: in out;
           Curve1 :    TheCurve;
           Domain1:    Domain      from IntRes2d;
	   Curve2 :    TheCurve;
           Domain2:    Domain      from IntRes2d;
	   TolConf:    Real        from Standard;
	   Tol    :    Real        from Standard)
	   
           is static; 

    Perform(me: in out;
           Curve1 :    TheCurve;
           Domain1:    Domain      from IntRes2d;
	   TolConf:    Real        from Standard;
	   Tol    :    Real        from Standard)
	   
           is static; 


    Perform(me: in out;
           Curve1 :    TheCurve;
           Domain1:    Domain      from IntRes2d;
	   Curve2 :    TheCurve;
           Domain2:    Domain      from IntRes2d;
	   TolConf:    Real        from Standard;
	   Tol    :    Real        from Standard;
           NbIter :    Integer     from Standard;
           DeltaU :    Real        from Standard;
           DeltaV :    Real        from Standard)
	   
           is static protected;    


    Perform(me: in out;
           Curve1 :    TheCurve;
           Domain1:    Domain      from IntRes2d;
	   TolConf:    Real        from Standard;
	   Tol    :    Real        from Standard;
           NbIter :    Integer     from Standard;
           DeltaU :    Real        from Standard;
           DeltaV :    Real        from Standard)
	   
           is static protected; 
           
       findIntersect( me: in out ;
           Curve1 :    TheCurve;
           Domain1:    Domain      from IntRes2d;
           Curve2 :    TheCurve;
           Domain2:    Domain      from IntRes2d;
		   TolConf:    Real        from Standard;
	       Tol    :    Real        from Standard;
           NbIter :    Integer     from Standard;
           DeltaU :    Real        from Standard;
           DeltaV :    Real        from Standard;
    	  thePoly1 :  ThePolygon2d  from  IntCurve; 
	      thePoly2 :  ThePolygon2d  from  IntCurve;
	      isFullRepresentation : Boolean from Standard)
	      returns Boolean is private;  
	      ---Purpose : Method to find intersection between two curves
	      --         :  returns false for case when some points of polygon
	      --         : were replaced on line and exact point of intersection was not found
	      --         : for case when point of intersection was found
	      --         : during prelimanary search for line (case of bad paramerization of Bspline for example). 
    
fields    

     DomainOnCurve1 : Domain from IntRes2d;      
     DomainOnCurve2 : Domain from IntRes2d;      
	  
end IntPolyPolyGen;





