-- Created on: 1997-04-17
-- Created by: Christophe MARION
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class FaceIterator from HLRBRep

uses
    Integer     from Standard,
    Boolean     from Standard,
    Orientation from TopAbs,
    WiresBlock  from HLRAlgo,
    EdgesBlock  from HLRAlgo,
    FaceData    from HLRBRep

is
    Create returns FaceIterator from HLRBRep;

    InitEdge(me : in out;
             fd :    out FaceData from HLRBRep)
	---Purpose: Begin an exploration of the edges of the face <fd>
    is static;
    
    MoreEdge(me) returns Boolean from Standard
	---C++: inline
    is static;
    
    NextEdge(me : in out)
    is static;
    
    BeginningOfWire(me) returns Boolean from Standard
	---Purpose: Returns True if the current edge is the first of a
	--          wire.
	--          
	---C++: inline
    is static;
    
    EndOfWire(me) returns Boolean from Standard
	---Purpose: Returns True if the current edge is the  last of a
	--          wire.
	--          
	---C++: inline
    is static;
    
    SkipWire(me : in out)
	---Purpose: Skip the current wire in the exploration.
	--          
	---C++: inline
    is static;
    
    Wire(me) returns any EdgesBlock from HLRAlgo
	---Purpose: Returns the edges of the current wire.
	--          
	---C++: inline
    is static;
    
    Edge(me) returns Integer from Standard
	---C++: inline
    is static;
    
    Orientation(me) returns Orientation from TopAbs
	---C++: inline
    is static;
	
    OutLine(me)
    returns Boolean from Standard
    	---C++: inline
    is static;

    Internal(me)
    returns Boolean from Standard
    	---C++: inline
    is static;

    Double(me)
    returns Boolean from Standard
    	---C++: inline
    is static;

    IsoLine(me)
    returns Boolean from Standard
    	---C++: inline
    is static;

fields
    iWire   : Integer    from Standard;
    nbWires : Integer    from Standard;
    iEdge   : Integer    from Standard;
    nbEdges : Integer    from Standard;
    myWires : WiresBlock from HLRAlgo;
    myEdges : EdgesBlock from HLRAlgo;
    
end FaceIterator;
