-- Created on: 1993-07-28
-- Created by: Martine LANGLOIS
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

private deferred class Root from StepToTopoDS

    ---Purpose : This class implements the common services for
    --           all classes of StepToTopoDS which report error
    --	    	  and sets and returns precision.

is

    Initialize returns Root from StepToTopoDS;

    IsDone(me) returns Boolean is static;
    ---C++: inline
    
    Precision(me) returns Real from Standard is static;
    ---Purpose : Returns the value of "MyPrecision"
    ---C++: inline
        
    SetPrecision(me : in out ; preci : Real from Standard) is static;
    ---Purpose : Sets the value of "MyPrecision"
    ---C++: inline
    
    MaxTol(me) returns Real from Standard is static;
    ---Purpose : Returns the value of "MaxTol"
    ---C++: inline
    
    SetMaxTol(me : in out ; maxpreci : Real from Standard) is static;
    ---Purpose : Sets the value of MaxTol
    ---C++: inline

fields

    done     : Boolean is protected;
    --Equal True if everything is ok, False otherwise.
    myPrecision : Real from Standard;    
    myMaxTol    : Real from Standard;

end Root;



