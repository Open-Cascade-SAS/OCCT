-- Created on: 1999-10-01
-- Created by: Vladislav ROMASHKO
-- Copyright (c) 1999-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ImportShape from QANewBRepNaming inherits TopNaming from QANewBRepNaming

    ---Purpose: This class provides a topological naming 
    --          of a Shape

uses 
 
    Shape     from TopoDS,
    Label     from TDF,
    LabelMap  from TDF,
    TagSource from TDF

is 
 
    Create returns ImportShape from QANewBRepNaming;    

    Create (ResultLabel : Label from TDF) 
    returns ImportShape from QANewBRepNaming;  

    Init (me : in out; ResultLabel : Label from TDF);
    

    Load (me; S : Shape from TopoDS);
    ---Purpose: Use this method for a topological naming of a Shape

    LoadPrime (me; S : Shape from TopoDS);

    LoadFirstLevel (me; S : Shape from TopoDS; Tagger : TagSource from TDF);

    LoadNextLevels (me; S : Shape from TopoDS; Tagger : TagSource from TDF);

    LoadC0Edges(me; S : Shape from TopoDS; 
    	     	       Tagger : TagSource from TDF);
    ---Purpose: Method for internal use. It is used by Load().
    --          It loads the edges which couldn't be uniquely identified as 
    --          an intersection of two faces.


    LoadC0Vertices (me; S : Shape from TopoDS; Tagger : TagSource from TDF);

    NamedFaces (me; theNamedFaces : in out LabelMap from TDF)
    returns Integer from Standard;

    NamedEdges (me; theNamedEdges : in out LabelMap from TDF)
    returns Integer from Standard;

    NamedVertices (me; theNamedVertices : in out LabelMap from TDF)
    returns Integer from Standard;

end ImportShape;	       
