-- File:	RWStepFEA_RWAlignedCurve3dElementCoordinateSystem.cdl
-- Created:	Thu Dec 12 17:51:03 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWAlignedCurve3dElementCoordinateSystem from RWStepFEA

    ---Purpose: Read & Write tool for AlignedCurve3dElementCoordinateSystem

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    AlignedCurve3dElementCoordinateSystem from StepFEA

is
    Create returns RWAlignedCurve3dElementCoordinateSystem from RWStepFEA;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : AlignedCurve3dElementCoordinateSystem from StepFEA);
	---Purpose: Reads AlignedCurve3dElementCoordinateSystem

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: AlignedCurve3dElementCoordinateSystem from StepFEA);
	---Purpose: Writes AlignedCurve3dElementCoordinateSystem

    Share (me; ent : AlignedCurve3dElementCoordinateSystem from StepFEA;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWAlignedCurve3dElementCoordinateSystem;
