-- Created on: 1991-10-04
-- Created by: Remi GILET
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class BParab  from GccInt  

inherits Bisec from GccInt 

     	---Purpose: Describes a parabola as a bisecting curve between two
    	-- 2D geometric objects (such as lines, circles or points).

uses Parab2d from gp,
     IType  from GccInt

is

Create(Parab : Parab2d) returns mutable BParab;
    	---Purpose: Constructs a bisecting curve whose geometry is the 2D parabola Parab.
    
Parabola(me) returns Parab2d from gp
    is redefined;
    	---Purpose: Returns a 2D parabola which is the geometry of this bisecting curve. 
    
ArcType(me) returns IType from GccInt
    is static;
    	---Purpose: Returns GccInt_Par, which is the type of any GccInt_BParab bisecting curve.

fields

    par : Parab2d from gp;
    	---Purpose: The bisecting line.

end BParab;    

