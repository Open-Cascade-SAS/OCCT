-- Created on: 1995-07-18
-- Created by: Modelistation
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

generic class   GenExtCC from Extrema 
(Curve1    as any;
 Tool1     as any;   -- as ToolCurve(Curve1)
 Curve2    as any;
 Tool2     as any;   -- as ToolCurve(Curve2)
 ArrayOfPnt as Transient from Standard; -- as returned by Extrema_CurveCache::Points()
 POnC      as any;
 Pnt       as any;
 Vec       as any)

	---Purpose: It calculates all the distance between two curves.
	--          These distances can be maximum or minimum.
uses SequenceOfReal from TColStd,
	 Vector from math
	
raises  InfiniteSolutions from StdFail,
    	NotDone           from StdFail,
    	OutOfRange        from Standard

is

    Create returns GenExtCC;
    	---Purpose: Calculates all the distances as above
    	--          between Uinf and Usup for C1 and  between Vinf and Vsup 
    	--          for C2.

    Create (C1: Curve1; C2: Curve2) returns GenExtCC;
      	---Purpose: It calculates all the distances.
        --          The function F(u,v)=distance(C1(u),C2(v)) has an 
        --          extremum when gradient(f)=0. The algorithm uses
        --          Evtushenko's global optimization solver.

    Create (C1: Curve1; C2: Curve2; Uinf, Usup, Vinf, Vsup: Real) returns GenExtCC;
    	---Purpose: Calculates all the distances as above
    	--          between Uinf and Usup for C1 and  between Vinf and Vsup 
    	--          for C2.

    SetParams (me: in out; C1: Curve1; C2: Curve2; Uinf, Usup, Vinf, Vsup: Real)
      ---Purpose: Set params in case of empty constructor is usage.
      is static;

    SetTolerance (me: in out; Tol: Real);
      ---Purpose:

    Perform (me: in out) is static;
    	---Purpose: Performs calculations.


    IsDone (me) returns Boolean
    	---Purpose: Returns True if the distances are found.
    	is static;

    NbExt (me) returns Integer
    	---Purpose: Returns the number of extremum distances.
    	raises  NotDone from StdFail,
	    	-- if IsDone(me)=False.
    	    	InfiniteSolutions from StdFail
		-- if IsParallel(me)= True.
    	is static;

    SquareDistance (me; N: Integer =1) returns Real
    	---Purpose: Returns the value of the Nth square extremum distance.
    	raises  NotDone from StdFail,
	    	-- if IsDone(me)=False.
    	    	InfiniteSolutions from StdFail,
		-- if IsParallel(me)= True and N > 1.
    	    	OutOfRange
		-- if N < 1 or N > NbExt(me)
    	is static;

    Points (me; N: Integer; P1,P2: out POnC)
    	---Purpose: Returns the points of the Nth extremum distance.
    	--          P1 is on the first curve, P2 on the second one.
    	raises  NotDone from StdFail,
	    	-- if IsDone(me)=False.
    	    	InfiniteSolutions from StdFail,
		-- if IsParallel(me)= True.
    	    	OutOfRange
		-- if N < 1 or N > NbExt(me)
    	is static;

fields
  myCurveMinTol : Real from Standard;
  myLowBorder : Vector from math;
  myUppBorder : Vector from math;
  myPoints1 : SequenceOfReal from TColStd;
  myPoints2 : SequenceOfReal from TColStd;
  myC : Address from Standard [2];
  myDone : Boolean;

end GenExtCC;
