-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class AutoDesignDateAndPersonItem from StepAP214 inherits SelectType from StepData

	-- <AutoDesignDateAndPersonItem> is an EXPRESS Select Type construct translation.
	-- it gathers : Product, ProductDefinition, ProductDefinitionFormation, Representation
	-- Rev4 adds : AutoDesignOrganizationAssignment


uses
     AutoDesignOrganizationAssignment from StepAP214,
     Product from StepBasic,
     ProductDefinition from StepBasic,
     ProductDefinitionFormation from StepBasic,
     Representation from StepRepr,
     AutoDesignDocumentReference from StepAP214,
     ExternallyDefinedRepresentation from StepRepr,
     ProductDefinitionRelationship from StepBasic,
     ProductDefinitionWithAssociatedDocuments from StepBasic

is

	Create returns AutoDesignDateAndPersonItem;
	---Purpose : Returns a AutoDesignDateAndPersonItem SelectType

	CaseNum (me; ent : Transient) returns Integer;
	---Purpose: Recognizes a AutoDesignDateAndPersonItem Kind Entity that is :
	-- 1     AutoDesignOrganizationAssignment from StepAP214,
	-- 2     Product from StepBasic,
	-- 3     ProductDefinition from StepBasic,
	-- 4     ProductDefinitionFormation from StepBasic,
	-- 5     Representation from StepRepr,
	-- 6     AutoDesignDocumentReference from StepAP214,
	-- 7     ExternallyDefinedRepresentation from StepRepr,
	-- 8     ProductDefinitionRelationship from StepBasic,
	-- 9     ProductDefinitionWithAssociatedDocuments from StepBasic
	--        0 else

     AutoDesignOrganizationAssignment (me) returns AutoDesignOrganizationAssignment from StepAP214;
     Product (me) returns Product from StepBasic;
     ProductDefinition (me) returns ProductDefinition from StepBasic;
     ProductDefinitionFormation (me) returns ProductDefinitionFormation from StepBasic;
     Representation (me) returns Representation from StepRepr;
     AutoDesignDocumentReference (me) returns AutoDesignDocumentReference from StepAP214;
     ExternallyDefinedRepresentation (me) returns ExternallyDefinedRepresentation from StepRepr;
     ProductDefinitionRelationship (me) returns ProductDefinitionRelationship from StepBasic;
     ProductDefinitionWithAssociatedDocuments (me) returns ProductDefinitionWithAssociatedDocuments from StepBasic;

end AutoDesignDateAndPersonItem;

