-- Created on: 2002-11-13
-- Created by: Galina KULIKOVA
-- Copyright (c) 2002-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class RemoveLocations from ShapeUpgrade inherits TShared from MMgt

	---Purpose: Removes all locations sub-shapes of specified shape

uses
    ShapeEnum from TopAbs,
    Shape from TopoDS,
    MapOfShape from TopTools,
    DataMapOfShapeShape from TopTools
is
    Create returns RemoveLocations from ShapeUpgrade;
    	---Purpose:Empy constructor
    
    Remove(me : mutable;theShape : Shape from TopoDS) returns Boolean;
    	---Purpose:Removes all location correspodingly to RemoveLevel.
    
    MakeNewShape(me : mutable;theShape , theAncShape: Shape from TopoDS; 
    	    	 theNewShape:in out Shape from TopoDS;theRemoveLoc : Boolean) 
    	    	     returns Boolean is private;
    
    GetResult(me) returns Shape from TopoDS;
    	---Purpose:Returns shape with removed locatins.
    	---C++: inline
	
    SetRemoveLevel(me: mutable; theLevel : ShapeEnum from TopAbs);
    	---Purpose:sets level starting with that location will be removed, 
    	--         by default TopAbs_SHAPE. In this case locations will be kept for specified shape
    	--         and if specified shape is TopAbs_COMPOUND for sub-shapes of first level.
    	---C++: inline
	
    RemoveLevel(me) returns ShapeEnum from TopAbs;
    	---Purpose:sets level starting with that location will be removed.Value of level can be set to
    	--         TopAbs_SHAPE,TopAbs_COMPOUND,TopAbs_SOLID,TopAbs_SHELL,TopAbs_FACE.By default TopAbs_SHAPE.
	--         In this case location will be removed for all shape types for exception of compound.
    	---C++: inline
    
	
    ModifiedShape (me; theInitShape : Shape from TopoDS) returns Shape from TopoDS;
    	---Purpose: Returns modified shape obtained from initial shape. 
	---C++: inline
    
fields
    myLevelRemoving : ShapeEnum from TopAbs;
    myShape : Shape from TopoDS;
    myMapNewShapes : DataMapOfShapeShape from TopTools;
    
end RemoveLocations;
