-- Created on: 1993-12-23
-- Created by: Gilles DEBARBOUILLE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

generic class MethodInstance from Dynamic (Dictionary as Transient)

inherits

    Method from Dynamic
    
	---Purpose: This  class describes the  facilities available to
	--          manipulate methods  objects. It is a generic class
	--          because the  creation of a MethodInstance requests
	--          a specific dictionary of  definitions. In a method
	--          instance,     it  is  only    possible   to    set
	--          VariableInstance which  are roughtly a copy of the
	--          variable  set in   the  method  definition  and  a
	--          pointer on the  variable, describing the signature
	--          of the complex method  in the process of build  or
	--          addressing the user value.

uses

    CString from Standard,
    OStream from Standard,
    Boolean from Standard,
    ModeEnum     from Dynamic,
    Parameter    from Dynamic,
    Variable     from Dynamic,
    VariableNode from Dynamic,
    AsciiString  from TCollection


is

    Create(atype : CString from Standard) returns mutable MethodInstance from Dynamic;
    
    ---Level: Public 
    
    --- Purpose: Creates a MethodInstance object  of the type <atype>.
    --  If  <atype>  is  not  defined in  the   dictionary, the object
    --  created will have no definition.

    Create(amethodinstance : MethodInstance from Dynamic) returns mutable MethodInstance from Dynamic;
    
    ---Level: Public 
    
    --- Purpose: Creates a MethodInstance with as definition the method 
    --           instance <amethodinstance>.

    Type(me) returns AsciiString from TCollection
    
    ---Level: Public 
    
    ---Purpose: Returns the type of object read in the definition.
    
    is redefined;
    
    Definition(me) returns Method from Dynamic
    
    ---Level: Public 
    
    ---Purpose: Returns   a    reference to  the   definition   of the
    --          MethodInstance.
    
    is static;
    
    Variable(me : mutable ; aparameter : Parameter from Dynamic
                          ; amode      : ModeEnum  from Dynamic
                          ; avariable  : Variable  from Dynamic)
    
    ---Level: Public 
    
    ---Purpose: Creates  and adds to  the  instance <me> the  variable
    --          instance  build  with  <aparameter> and  <amode>   and
    --          adresses the variable .
    
    is static;
    
    Value(me ; aname      : CString from Standard
    	     ; aparameter : out any Parameter from Dynamic 
    	     ; amode      : out ModeEnum      from Dynamic
             ; avariable  : out any Variable  from Dynamic) returns Boolean
    
    ---Level: Public 
    
    ---Purpose: Returns True, if  there is  a variable instance  named
    --          <aname>, False otherwise.   It returns in the argument
    --          <aparameter> the signature of the variable, in <amode>
    --          the variable is  in, out, inout, internal or  constant
    --          and in  <avariable>,  the reference  to the  effective
    --          value   used by the   instance or  a reference  to the
    --          variable defining the  signature of the complex method
    --          using this instance of method.
    
    is static;
    
    Value(me ; aname         : CString from Standard
    	     ; aparameter    : out any Parameter     from Dynamic 
    	     ; amode         : out ModeEnum          from Dynamic
             ; avariablenode : out any VariableNode  from Dynamic) returns Boolean from Standard
    
    ---Level: Public 
    
    ---Purpose: Returns True, if  there is  a variable instance  named
    --          <aname>, False otherwise.   It returns in the argument
    --          <aparameter> the signature of the variable, in <amode>
    --          the  variable is in, out,  inout, internal or constant
    --          and in <avariablenode>,  the  head  of the   effective
    --          referenced value  used by the instance  or the head of
    --          the variables reference  defining the signature of the
    --          complex method using this instance of method.
    
    is static;
    
    Dump(me ; astream : in out OStream from Standard)

    ---Level: Internal 
    
    ---Purpose: Useful for debugging.

    is redefined;
    
fields

    thedefinition : Method from Dynamic;

end MethodInstance;
