-- Created on: 2001-04-24
-- Created by: Christian CAILLET
-- Copyright (c) 2001-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ValueQualifier  from StepShape    inherits SelectType  from StepData

    ---Purpose : Added for Dimensional Tolerances

uses
    PrecisionQualifier from StepShape,
    TypeQualifier from StepShape

is

    Create returns ValueQualifier from StepShape;

    CaseNum (me; ent : Transient) returns Integer;
    ---Purpose : Recognizes a kind of ValueQualifier Select Type :
    --           1 -> PrecisionQualifier from StepShape
    --           2 -> TypeQualifier from StepShape
    --           3 -> UnceraintyQualifier .. not yet implemented

    PrecisionQualifier (me) returns PrecisionQualifier from StepShape;
    ---Purpose : Returns Value as PrecisionQualifier

    TypeQualifier (me) returns TypeQualifier from StepShape;
    ---Purpose : Returns Value as TypeQualifier

end ValueQualifier;
