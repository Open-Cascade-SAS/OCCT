-- Created on: 1993-01-27
-- Created by: Jean-Louis Frenkel
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ShapeTool from Prs3d


uses
    Shape             from TopoDS,
    Face              from TopoDS,
    Edge              from TopoDS,
    Vertex            from TopoDS,
    HSequenceOfShape  from TopTools,
    Box               from Bnd,
    Location          from TopLoc,
    Triangulation     from Poly,
    PolygonOnTriangulation     from Poly,
    Polygon3D         from Poly,
    HArray1OfInteger  from TColStd,
    Explorer          from TopExp,
    IndexedDataMapOfShapeListOfShape from TopTools,
    IndexedMapOfShape                from TopTools

	---Purpose: 
is

    Create ( TheShape: Shape from TopoDS) returns ShapeTool from Prs3d;
    InitFace (me: in out);
    MoreFace (me) returns Boolean from Standard;
    NextFace (me: in out);
    GetFace(me) returns Face from TopoDS;
    	---C++: return const&
    FaceBound(me) returns Box from Bnd;
    IsPlanarFace(me) returns Boolean from Standard;

    InitCurve (me: in out);
    MoreCurve (me) returns Boolean from Standard;
    NextCurve (me: in out);
    GetCurve(me) returns Edge from TopoDS;
    	---C++: return const&
    CurveBound(me) returns Box from Bnd;
    Neighbours(me) returns Integer from Standard;   
    FacesOfEdge(me) returns HSequenceOfShape from TopTools;

    InitVertex(me: in out);
    MoreVertex(me) returns Boolean from Standard;
    NextVertex(me: in out);
    GetVertex(me) returns Vertex from TopoDS;
    	---C++: return const&

    HasSurface(me) returns Boolean;
    
    CurrentTriangulation(me; l: out Location from TopLoc) 
    returns Triangulation from Poly;

    HasCurve(me) returns Boolean;

    PolygonOnTriangulation(me; Indices: out PolygonOnTriangulation from  Poly;
    	    	    	       T:       out Triangulation          from Poly; 
			       l:       out Location               from TopLoc); 
			       
    Polygon3D(me; l: out Location from TopLoc) 
    returns Polygon3D from Poly;

fields
    myShape:        Shape                            from TopoDS;
    myFaceExplorer: Explorer                         from TopExp;
    myEdgeMap:      IndexedDataMapOfShapeListOfShape from TopTools;
    myVertexMap:    IndexedMapOfShape                from TopTools;
    myEdge :        Integer                          from Standard;
    myVertex :      Integer                          from Standard;

end ShapeTool from Prs3d;
