-- Created on: 1994-12-22
-- Created by: Christian CAILLET
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package STEPSelections

    ---Purpose : Step Selections

uses 
    
    MMgt, 
    TCollection, 
    TColStd,
    Interface, 
    IFGraph,
    IFSelect, 
    StepSelect,
    StepBasic,
    StepShape,
    StepGeom,
    StepRepr,
    StepData,
    XSControl

is

    class SelectFaces;
    
    class SelectDerived;
    
    class SelectGSCurves;
    
    class SelectAssembly;
    
    class SelectInstances;
     
    class SelectForTransfer;
    -- Classes that are intended for assembly exploration
    
    class SequenceOfAssemblyLink instantiates
    	Sequence from TCollection (AssemblyLink from STEPSelections);
	
    class HSequenceOfAssemblyLink instantiates
    	HSequence from TCollection (AssemblyLink           from STEPSelections,
	    	    	    	    SequenceOfAssemblyLink from STEPSelections);
				    
    class SequenceOfAssemblyComponent instantiates
    	Sequence from TCollection (AssemblyComponent from STEPSelections);
    
    class AssemblyComponent;
    
    class AssemblyLink;
    
    class AssemblyExplorer;

    class Counter;

end STEPSelections;
