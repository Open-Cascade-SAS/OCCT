-- Created on: 2009-04-06
-- Created by: Sergey ZARITCHNY
-- Copyright (c) 2009-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Point from TDataXtd inherits Attribute from TDF

	---Purpose: 
    	-- The basis to define a point attribute.
    	-- The topological attribute must contain a vertex.
    	-- You use this class to create reference points in a design.
	--          
	--  Warning:  Use TDataXtd_Geometry  attribute  to retrieve the
	--          gp_Pnt of the Point attribute

uses Attribute       from TDF,
     Label           from TDF,
     GUID            from Standard,
     Pnt             from gp,
     DataSet         from TDF,
     RelocationTable from TDF

is    


    ---Purpose: class methods
    --          =============
      
    GetID(myclass)    
    	---C++: return const & 
    returns GUID from Standard;   
    	---Purpose:
    	-- Returns the GUID for point attributes.

    Set (myclass ; label : Label from TDF) 
    	---Purpose: 
    	-- Sets the label Label as a point attribute.
    	-- If no object is found, a point attribute is created.
    returns Point from TDataXtd;      

    Set (myclass ; label : Label from TDF; P : Pnt from gp)
    	---Purpose: 
    	-- Sets the label Label as a point attribute containing the point P.
    	-- If no object is found, a point attribute is created.
    returns Point from TDataXtd;    

    ---Purpose: Point methods
    --          =============    

    Create
    returns Point from TDataXtd;  

    ---Category: TDF_Attribute methods
    --           =====================

    
    ID (me)  
    	---C++: return const & 
    returns GUID from Standard;

    Restore (me: mutable; With : Attribute from TDF);

    NewEmpty (me)
    returns Attribute from TDF;

    Paste (me; Into : Attribute from TDF;
	       RT   : RelocationTable from TDF);  

    Dump (me; anOS : in out OStream from Standard) 
    	returns OStream from Standard
    	is redefined;
	---C++: return &

end Point;

