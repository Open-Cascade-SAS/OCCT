-- Created on: 1995-03-15
-- Created by: Laurent PAINNOT
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PolygonOnClosedTriangulation from BRep 
    
    inherits PolygonOnTriangulation  from  BRep


    	---Purpose: A representation by two arrays of nodes on a 
    	--          triangulation.


uses HArray1OfInteger       from TColStd,
     Array1OfInteger        from TColStd,
     Location               from TopLoc,
     CurveRepresentation    from BRep,
     Triangulation          from Poly,
     PolygonOnTriangulation from Poly


is

    Create(P1, P2 : PolygonOnTriangulation from Poly;
    	   Tr: Triangulation          from Poly;
	   L : Location               from TopLoc)
    returns mutable PolygonOnClosedTriangulation from BRep;


    IsPolygonOnClosedTriangulation(me)    returns Boolean
    	---Purpose: Returns True.
    is redefined;


    PolygonOnTriangulation2(me: mutable; P2: PolygonOnTriangulation from  Poly)
    is redefined;


    PolygonOnTriangulation2(me) returns any PolygonOnTriangulation from  Poly
    	---C++: return const&
    is redefined;


    Copy(me) returns mutable CurveRepresentation from BRep is redefined;
	---Purpose: Return a copy of this representation.


fields

myPolygon2: PolygonOnTriangulation from Poly;

end PolygonOnClosedTriangulation;
