-- File     : Prs2d_Length.cdl
-- Created  : April  2000
-- Author   : Tanya COOL
---Copyright: Matra Datavision 2000

class Length from Prs2d inherits Dimension from Prs2d

 ---Purpose: Constructs the primitive Length

uses

	Drawer	           from Graphic2d,
	GraphicObject      from Graphic2d,
	Pnt2d              from gp,
	Lin2d              from gp,
	ExtendedString     from TCollection,
	ArrowSide          from Prs2d,
	TypeOfDist         from Prs2d,
	TypeOfArrow        from Prs2d,
    	FStream            from Aspect 

is
	Create( aGraphicObject: GraphicObject  from Graphic2d;
	        anAttachPnt1  : Pnt2d          from gp;
            	anAttachPnt2  : Pnt2d          from gp;
          	aText         : ExtendedString from TCollection;
		aTxtScale     : Real           from Standard = 5.0;
		aLength       : Real           from Standard = 0.0;
	        aTypeDist     : TypeOfDist     from Prs2d = Prs2d_TOD_AUTOMATIC;
		anArrAngle    : Real           from Standard = 20.0;
		anArrLength   : Real           from Standard = 25.0;
	    	anArrType     : TypeOfArrow    from Prs2d = Prs2d_TOA_OPENED;
		anArrow       : ArrowSide      from Prs2d = Prs2d_AS_BOTHAR;
		IsReverseArrow: Boolean        from Standard = Standard_False )

	returns mutable Length from Prs2d;

    	---Purpose: Initializes the length dimension between points 
    	--          anAttachPnt1 and anAttachPnt2. 
    	--          aLength is length of the attach lines 
    	--          aTypeDist defines the orientation of the displayed length: 
    	--          AIS2D_TOD_AUTOMATIC
    	--          AIS2D_TOD_OBLIQUE
    	--          AIS2D_TOD_HORIZONTAL
    	--          AIS2D_TOD_VERTICAL
    	--          anArrow defines the number of arrows (one, two or none)

    	Create( aGraphicObject: GraphicObject  from Graphic2d;
	    	anAttachPnt   : Pnt2d          from gp;
            	anAttachLin   : Lin2d          from gp;
            	aText         : ExtendedString from TCollection;
		aTxtScale     : Real           from Standard = 10.0;
	        aLenAttachLin : Real           from Standard = 0.0;
		anArrAngle    : Real           from Standard = 20.0;
		anArrLength   : Real           from Standard = 25.0;
	        anArrType     : TypeOfArrow    from Prs2d = Prs2d_TOA_OPENED;
	        anArrow       : ArrowSide      from Prs2d = Prs2d_AS_BOTHAR;
	        IsReverseArrow: Boolean        from Standard = Standard_False ) 

       returns mutable Length from Prs2d;

    	---Purpose: Initializes the length dimension between point 
    	--          anAttachPnt1 and line defined anAttachLin. 
    	--          aLenAttachLin is length of the attach lines 
    
    	Create( aGraphicObject: GraphicObject  from Graphic2d;
	        anAttachLin1  : Lin2d          from gp;
	        anAttachLin2  : Lin2d          from gp;
            	aText         : ExtendedString from TCollection;
		aTxtScale     : Real           from Standard = 10.0;
	        aLenAttachLin : Real           from Standard = 0.0;
		anArrAngle    : Real           from Standard = 20.0;
		anArrLength   : Real           from Standard = 25.0;
	    	anArrType     : TypeOfArrow    from Prs2d = Prs2d_TOA_OPENED;
	        anArrow       : ArrowSide from Prs2d = Prs2d_AS_BOTHAR;
	        IsReverseArrow: Boolean from Standard = Standard_False ) 

        returns mutable Length from Prs2d;

    	---Purpose: Initializes the length dimension between line 
    	--          anAttachLin1 and line defined anAttachLin2. 
    	--          aLenAttachLin is length of the attach lines 
  
	--------------------------
	-- Category: Draw and Pick
	--------------------------

    Draw( me : mutable; aDrawer: Drawer from Graphic2d ) is static protected;
    	---Level: Internal
    	---Purpose: Draws the length <me>.

    DrawElement( me : mutable; aDrawer: Drawer from Graphic2d;
                 anIndex: Integer from Standard) is redefined protected;
    	---Level: Internal
    	---Purpose: Draws element <anIndex> of the length <me>.

    DrawVertex( me : mutable; aDrawer: Drawer from Graphic2d;
                anIndex: Integer from Standard) is redefined protected;
    	---Level: Internal
    	---Purpose: Draws vertex <anIndex> of the length <me>.

    Pick( me : mutable; X, Y: ShortReal from Standard;
	  aPrecision: ShortReal from Standard;
	  aDrawer: Drawer from Graphic2d) returns Boolean from Standard
	  is static protected;
    	---Level: Internal
    	---Purpose: Returns Standard_True if the length <me> is picked,
    	--	    Standard_False if not.

    GetPntProject( me: mutable; aLength: Real from Standard ) is private;
    ComputeArrows( me: mutable; isnotPoints: Boolean from Standard ) is private;

	--------------------------------------------
	-- Category: Modification of the properties
	--------------------------------------------
	
    SetAttachLinLength( me: mutable; aLength: Real from Standard );
    	    ---Level: Public
	    ---Purpose: Sets the length of attachment lines

    Save( me; aFStream: in out FStream from Aspect ) is virtual;
														
    CalcTxtPos(me:mutable; theFromAbs: 
       	    Boolean from Standard=Standard_False) 
    	---C++: inline
    	is redefined protected;
	
    LineCoord( me ; aFirstPnt, aSecondPnt: in out Pnt2d from gp );
       	---Level: Internal
	---Purpose: returns coordinates of points, which are begining
	--          and end of arrow
	
    CallOutCoord( me ; aFirstPnt, aSecondPnt: in out Pnt2d from gp );
       	---Level: Internal
	---Purpose: returns coordinates of points, which are begining
	--          and end of arrow
    
    TypeOfDist(me) returns TypeOfDist;
      	---Level: Internal
	
	
fields
 
	myX1           : ShortReal         from Standard;
	myY1           : ShortReal         from Standard;
	myX2           : ShortReal         from Standard;
	myY2           : ShortReal         from Standard;
	myAX1          : ShortReal         from Standard;
	myAY1          : ShortReal         from Standard;
	myAX2          : ShortReal         from Standard;
	myAY2          : ShortReal         from Standard;
  	myTypeDist     : TypeOfDist        from Prs2d;
    	myXT1          : ShortReal         from Standard;
    	myYT1          : ShortReal         from Standard;
    	myXT2          : ShortReal         from Standard;
    	myYT2          : ShortReal         from Standard;

end Length from Prs2d;
    
