-- Created on: 1998-05-06
-- Created by: Christian CAILLET
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



package SWDRAW

    ---Purpose: Provides DRAW interface to the functionalities of Shape Healing
    --          toolkit (SHAPEWORKS Delivery Unit).
    --          
    --          Classes prefixed with Shape* corresponds to the packages of
    --          Shape Healing.

uses  TCollection, TColStd, TopoDS, TopTools, Draw, ShapeProcessAPI

is

    class ShapeTool;
    	---Purpose: Contains commands to activate Topology/Geometry not
    	--          Shape Healing

    class ShapeAnalysis;
    	---Purpose: Contains commands to activate package ShapeAnalysis

    class ShapeBuild;
    	---Purpose: Contains commands to activate package ShapeBuild

    class ShapeConstruct;
    	---Purpose: Contains commands to activate package ShapeConstruct

    class ShapeCustom;
    	---Purpose: Contains commands to activate package ShapeCustom

    class ShapeExtend;
    	---Purpose: Contains commands to activate package ShapeExtend

    class ShapeFix;
    	---Purpose: Contains commands to activate package ShapeFix

    class ShapeUpgrade;
    	---Purpose: Contains commands to activate package ShapeUpgrade

    class ShapeProcess;
    	---Purpose: Contains commands to activate package ShapeProcess
    
    class ShapeProcessAPI;
    	---Purpose: Contains commands to activate package ShapeProcessAPI
	
    class ToVRML;
    	---Purpose: A utility which writes a Shape to VRML format
    	---Remark : It can be placed elsewhere, while it depends on
    	--          only BRepMesh i.e. TOPOLOGY

    Init (theCommands: in out Interpretor from Draw);
    	---Purpose: Loads commands defined in SWDRAW

    GroupName returns CString is private;
    	---Purpose: Returns the name of the DRAW group accumulating the
    	--          commands from the classes prefixed with Shape*.
	--          Returns "Shape Healing".
	
end SWDRAW;
