-- Created on: 2001-09-11
-- Created by: Julia DOROVSKIKH
-- Copyright (c) 2001-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class LocationDriver from XmlMXCAFDoc  inherits ADriver from XmlMDF



        ---Purpose: Attribute Driver.

uses    Location         from TopLoc,
        Element          from XmlObjMgt,
        SRelocationTable from XmlObjMgt,
        RRelocationTable from XmlObjMgt,
        Persistent       from XmlObjMgt,
        MessageDriver    from CDM,
        Attribute        from TDF,
        LocationSetPtr   from TopTools

is
    Create (theMessageDriver:MessageDriver from CDM)
        returns mutable LocationDriver from XmlMXCAFDoc;



    NewEmpty (me)  returns mutable Attribute from TDF;




    Paste(me; Source     : Persistent from XmlObjMgt;
              Target     : mutable Attribute from TDF;
              RelocTable : out RRelocationTable from XmlObjMgt)
        returns Boolean from Standard;

    Paste(me; Source     : Attribute from TDF;
              Target     : in out Persistent from XmlObjMgt;
              RelocTable : out SRelocationTable from XmlObjMgt);

    Translate (me; theLoc    : Location from TopLoc;
                        theParent : in out Element from XmlObjMgt;
                        theMap    : in out SRelocationTable from XmlObjMgt);
        ---Purpose: Translate a non storable Location to a storable Location.
        ---Level: Internal

    Translate (me; theParent : Element from XmlObjMgt;
                        theLoc    : in out Location from TopLoc;
                        theMap    : in out RRelocationTable from XmlObjMgt)
    returns Boolean from Standard;
        ---Purpose: Translate a storable Location to a non storable Location.
        ---Level: Internal

    SetSharedLocations(me: mutable;
                       theLocations:  in LocationSetPtr  from TopTools);
    ---C++: inline

fields
    myLocations : LocationSetPtr   from TopTools;
end LocationDriver;
