-- Created on: 1995-01-17
-- Created by: GG
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class MarkMap from Xw inherits Transient

	---Version: 0.0

	---Purpose: This class defines a MarkMap object.

	---Keywords:
	---Warning:
	---References:

uses

	MarkMap		from Aspect,
	MarkMapEntry	from Aspect,
	MarkerStyle 	from Aspect

raises

	MarkMapDefinitionError	from Aspect,
	BadAccess		from Aspect

is

	Create
	returns mutable MarkMap from Xw
	is protected ;
	---Level: Internal

	Create ( Connexion : CString from Standard ) 
	returns mutable MarkMap from Xw 
	---Level: Public
	---Purpose: Creates a MarkMap with unallocated MarkMapEntry.
	--  Warning: Raises if MarkMap creation failed according
	--	    to the supported hardware
	raises MarkMapDefinitionError from Aspect ;

	SetEntry ( me : mutable ; 
		   anEntry : MarkMapEntry from Aspect )
	---Level: Public
	---Purpose: Modifies an entry already defined or Add the Entry
	--	    in the marker map <me> if it don't exist.
	--  Warning: Raises if MarkMap size is exceeded,
	--	    or MarkMap is not defined properly,
	--	    or MarkMapEntry Index is out of range according
	--	    to the supported hardware
	raises BadAccess from Aspect is virtual;

	SetEntries ( me : mutable ; 
		     aMarkmap : MarkMap from Aspect ) 
	---Level: Public
	---Purpose: Modifies all entries from a new Markmap
	--  Warning: Raises if MarkMap size is exceeded,
	--	    or MarkMap is not defined properly,
	--	    or One of new MarkMapEntry Index is out of range according
	--	    to the supported hardware
	raises BadAccess from Aspect is virtual;

	Destroy ( me : mutable ) is virtual;
	---Level: Public
	---Purpose: Destroies the Markmap
	---C++: alias ~

	----------------------------
	-- Category: Inquire methods
	----------------------------

	FreeMarkers ( me )
	returns Integer from Standard 
	---Level: Public
	---Purpose: Returns the Number of Free Marks in the Typemap
	--	    depending of the HardWare
	--  Warning: Raises if MarkMap is not defined properly
	raises BadAccess from Aspect is static;

	ExtendedMarkMap ( me )
	returns Address from Standard
	is static protected ;
	---Level: Internal
	---Purpose: Returns extended data markermap structure pointer.
	---Category: Inquire methods


fields

	MyExtendedDisplay	: Address from Standard ;
	MyExtendedMarkMap 	: Address from Standard ;

friends

	class GraphicDevice from Xw

end MarkMap ;
