-- Created on: 1993-03-10
-- Created by: JCV
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class  SurfaceOfLinearExtrusion from Geom inherits SweptSurface from Geom

        --- Purpose : Describes a surface of linear extrusion ("extruded
        -- surface"), e.g. a generalized cylinder. Such a surface
        -- is obtained by sweeping a curve (called the "extruded
        -- curve" or "basis") in a given direction (referred to as
        -- the "direction of extrusion" and defined by a unit vector).
        -- The u parameter is along the extruded curve. The v
        -- parameter is along the direction of extrusion.
        -- The parameter range for the u parameter is defined
        -- by the reference curve.
        -- The parameter range for the v parameter is ] -
        -- infinity, + infinity [.
        -- The position of the curve gives the origin of the v parameter.
        -- The surface is "CN" in the v parametric direction.
        -- The form of a surface of linear extrusion is generally a
        -- ruled surface (GeomAbs_RuledForm). It can be:
        -- - a cylindrical surface, if the extruded curve is a circle,
        --   or a trimmed circle, with an axis parallel to the
        --   direction of extrusion (GeomAbs_CylindricalForm), or
        -- - a planar surface, if the extruded curve is a line
        --   (GeomAbs_PlanarForm).
        -- Note: The surface of extrusion is built from a copy of
        -- the original basis curve, so the original curve is not
        -- modified when the surface is modified.
        -- Warning
        -- Degenerate surfaces are not detected. A degenerate
        -- surface is obtained, for example, when the extruded
        -- curve is a line and the direction of extrusion is parallel
        -- to that line.

uses Ax1         from gp, 
     Ax2         from gp,
     Dir         from gp,
     Pnt         from gp,
     Trsf        from gp,
     GTrsf2d     from gp,
     Vec         from gp,
     Curve       from Geom,
     Geometry    from Geom,
   BSplineCurve  from  Geom,
     Shape       from GeomAbs,
      CurveType  from  GeomAbs 


raises RangeError          from Standard,
       UndefinedDerivative from Geom

is

  Create (C : Curve; V : Dir)   returns mutable SurfaceOfLinearExtrusion;
        --- Purpose :
        --  V is the direction of extrusion.
        --  C is the extruded curve.
        --  The form of a SurfaceOfLinearExtrusion can be :
        --  . ruled surface (RuledForm),
        --  . a cylindrical surface if the extruded curve is a circle or
        --    a trimmed circle (CylindricalForm),
        --  . a plane surface if the extruded curve is a Line (PlanarForm).
        --  Warnings :
        --  Degenerated surface cases are not detected. For example if the
        --  curve C is a line and V is parallel to the direction of this
        --  line.



  SetDirection (me : mutable; V : Dir);
       --- Purpose : Assigns V as the "direction of extrusion" for this
       -- surface of linear extrusion.

  SetBasisCurve (me : mutable; C : Curve);
        --- Purpose : Modifies this surface of linear extrusion by redefining
        -- its "basis curve" (the "extruded curve").


  UReverse (me : mutable);
        --- Purpose :  Changes the orientation of this surface of linear
        -- extrusion in the u  parametric direction. The
        -- bounds of the surface are not changed, but the given
        -- parametric direction is reversed. Hence the
        -- orientation of the surface is reversed.
        -- In the case of a surface of linear extrusion:
        -- - UReverse reverses the basis curve, and
        -- - VReverse reverses the direction of linear extrusion.


  UReversedParameter (me; U : Real) returns Real;
	---Purpose: Computes the u parameter on the modified
        -- surface, produced by reversing its u  parametric
        -- direction, for any point of u parameter U  on this surface of linear extrusion.
        -- In the case of an extruded surface:
        -- - UReverseParameter returns the reversed
        --   parameter given by the function
        --   ReversedParameter called with U on the basis   curve,
  
  VReverse (me : mutable);
        --- Purpose : Changes the orientation of this surface of linear
        -- extrusion in the v parametric direction. The
        -- bounds of the surface are not changed, but the given
        -- parametric direction is reversed. Hence the
        -- orientation of the surface is reversed.
        -- In the case of a surface of linear extrusion:
        -- - UReverse reverses the basis curve, and
        -- - VReverse reverses the direction of linear extrusion.


  VReversedParameter (me; V : Real) returns Real;
	---Purpose: Computes the v parameter on the modified
        -- surface, produced by reversing its u v parametric
        -- direction, for any point of v parameter V on this surface of linear extrusion.
        -- In the case of an extruded surface VReverse returns -V.
	
  
  Bounds (me; U1, U2, V1, V2 : out Real);
        --- Purpose : Returns the parametric bounds U1, U2, V1 and V2 of
        -- this surface of linear extrusion.
        -- A surface of linear extrusion is infinite in the v
        -- parametric direction, so:
        --     - V1 = Standard_Real::RealFirst()
        -- - V2 = Standard_Real::RealLast().


  IsUClosed (me)   returns Boolean;
        --- Purpose:  IsUClosed returns true if the "basis curve" of this
        -- surface of linear extrusion is closed.


  IsVClosed (me)  returns Boolean;
        --- Purpose : IsVClosed always returns false.


  IsCNu (me; N : Integer)  returns Boolean
        --- Purpose : IsCNu returns true if the degree of continuity for the
        -- "basis curve" of this surface of linear extrusion is at least N.
        --  Raises RangeError if N < 0.
     raises RangeError;


  IsCNv (me; N : Integer)     returns Boolean;
        --- Purpose : IsCNv always returns true.


  IsUPeriodic (me)   returns Boolean;
        --- Purpose : IsUPeriodic returns true if the "basis curve" of this
        -- surface of linear extrusion is periodic.


  IsVPeriodic (me)   returns Boolean;
        --- Purpose : IsVPeriodic always returns false.


  UIso (me; U : Real)  returns mutable Curve;
        --- Purpose : Computes the U isoparametric curve of this surface
        -- of linear extrusion. This is the line parallel to the
        -- direction of extrusion, passing through the point of
        -- parameter U of the basis curve.


  VIso (me; V : Real)   returns mutable Curve;
        --- Purpose : Computes the V isoparametric curve of this surface
        -- of linear extrusion. This curve is obtained by
        -- translating the extruded curve in the direction of
        -- extrusion, with the magnitude V.


  D0 (me; U, V : Real; P : out Pnt);
        --- Purpose :
        --  Computes the  point P (U, V) on the surface.
        --  The parameter U is the parameter on the extruded curve.
        --  The parametrization V is a linear parametrization, and
        --  the direction of parametrization is the direction of
        --  extrusion. If the point is on the extruded curve, V = 0.0


  D1 (me; U, V : Real; P : out Pnt; D1U, D1V : out Vec)
        --- Purpose :
        --  Computes the current point and the first derivatives in the
        --  directions U and V.
        --  Raises UndefinedDerivative if the continuity of the surface is not C1.
     raises UndefinedDerivative;


  D2 (me; U, V : Real; P : out Pnt; D1U, D1V, D2U, D2V, D2UV : out Vec)
        --- Purpose ;
        --  Computes the current point, the first and the second derivatives 
        --  in the directions U and V.
        --  Raises UndefinedDerivative if the continuity of the surface is not C2.
     raises UndefinedDerivative;


  D3 (me; U, V : Real;  P : out Pnt; 
      D1U, D1V, D2U, D2V, D2UV, D3U, D3V, D3UUV, D3UVV : out Vec)
        --- Purpose :
        --  Computes the current point, the first,the second and the third 
        --  derivatives in the directions U and V.
        --  Raises UndefinedDerivative if the continuity of the surface is not C3.
     raises UndefinedDerivative;


  DN (me; U, V : Real; Nu, Nv : Integer)  returns Vec
        --- Purpose :
        --  Computes the derivative of order Nu in the direction u 
        --  and Nv in the direction v.
        --  Raises UndefinedDerivative if the continuity of the surface is not CNu in the u
        --  direction and CNv in the v direction.
        --- Raises RangeError if Nu + Nv < 1 or Nu < 0 or Nv < 0.

     raises UndefinedDerivative,
            RangeError;

 

  LocalD0 (me; U, V : Real; USide : Integer;
    	       P : out Pnt);
   	---Purpose : The following  functions  evaluates the  local
    	-- derivatives on surface. Useful to manage discontinuities
	-- on the surface.
	--           if    Side  =  1  ->  P  =  S( U+,V )
        --           if    Side  = -1  ->  P  =  S( U-,V )
	--           else  P  is betveen discontinuities
	--           can be evaluated using methods  of
    	--           global evaluations    P  =  S( U ,V )
    		
  LocalD1 (me; U, V : Real;  USide : Integer;
          P : out Pnt; D1U, D1V : out Vec);
     	
  LocalD2 (me; U, V : Real; USide : Integer;
           P : out Pnt; D1U, D1V, D2U, D2V, D2UV : out Vec);
     	
  LocalD3 (me; U, V : Real; USide : Integer;
           P : out Pnt; D1U, D1V, D2U, D2V, D2UV, D3U, D3V, D3UUV, D3UVV :
           out Vec);
     	
  LocalDN (me; U, V : Real; USide : Integer; 
           Nu, Nv : Integer)
     returns Vec;
     	 
  Transform(me : mutable; T : Trsf);
        ---Purpose: Applies the transformation T to this surface of linear extrusion.
        
  TransformParameters(me; U,V : in out Real; T : Trsf from gp)
	---Purpose: Computes the  parameters on the  transformed  surface for
	--          the transform of the point of parameters U,V on <me>.
	--          
	--          me->Transformed(T)->Value(U',V')
	--          
	--          is the same point as
	--          
	--          me->Value(U,V).Transformed(T)
	--          
	--          Where U',V' are the new values of U,V after calling
	--          
	--          me->TranformParameters(U,V,T)
	--          
	--          This methods multiplies : 
	--          U by BasisCurve()->ParametricTransformation(T)
	--          V by T.ScaleFactor()
     is redefined;  

  ParametricTransformation(me; T : Trsf from gp) returns GTrsf2d from gp
	---Purpose: Returns a 2d transformation  used to find the  new
	--          parameters of a point on the transformed surface.
	--          
	--          me->Transformed(T)->Value(U',V')
	--          
	--          is the same point as
	--          
	--          me->Value(U,V).Transformed(T)
	--          
	--          Where U',V' are  obtained by transforming U,V with
	--          th 2d transformation returned by
	--          
	--          me->ParametricTransformation(T)
	--          
	--          This  methods  returns  a scale  
	--          U by BasisCurve()->ParametricTransformation(T)
	--          V by T.ScaleFactor()
     is redefined;  
  


  Copy (me)  returns mutable like me;
        ---Purpose: Creates a new object which is a copy of this surface of linear extrusion.
    
end;  
 
