-- Created on: 2000-10-24
-- Created by: Peter KURNEV
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class CompareRange from IntTools 

	---Purpose: Auxiliary class to provide a sorting Ranges, 
        --          taking  into  account a value of Left .   

uses
    Range from IntTools
--raises

is
    Create   
    	returns CompareRange from IntTools; 
	---Purpose:
	--- Empty constructor
	---
	 
    Create  (aTol:Real from Standard) 
    	returns CompareRange from IntTools;
	---Purpose:
	--- Initializes me by tolerance
	---
	 
    IsLower (me; Left, Right: Range from IntTools)
	---Purpose: 
    	--- Returns True if <Left> is lower than <Right>.
	---
    	returns Boolean from Standard;
    
    IsGreater (me; Left, Right: Range from IntTools)
	---Level: Public
	---Purpose: 
    	--- Returns True if <Left> is greater than <Right>.
	---
    	returns Boolean from Standard;

    IsEqual(me; Left, Right: Range from IntTools)
	---Level: Public
	---Purpose: 
    	--- Returns True when <Right> and <Left> are equal.
	---
    	returns Boolean from Standard ;

fields
    myTol: Real from Standard; 

end CompareRange;
