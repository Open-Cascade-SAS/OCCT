-- Created on: 1995-08-25
-- Created by: Remi LEQUETTE
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class HCurve from GeomAdaptor inherits GHCurve from GeomAdaptor

    	---Purpose: An interface between the services provided by any
    	-- curve from the package Geom and those required of
    	-- the curve by algorithms which use it.

uses
    Curve from Geom,
    Curve from GeomAdaptor

raises
    ConstructionError from Standard

is

    Create returns mutable HCurve from GeomAdaptor;
    	---C++: inline
    
    Create( AS : Curve from GeomAdaptor) returns mutable HCurve from GeomAdaptor;
    	---C++: inline

    Create( S : Curve from Geom) returns mutable HCurve from GeomAdaptor;
    	---C++: inline
    
    Create( S : Curve from Geom; UFirst,ULast : Real) 
    returns  mutable HCurve from GeomAdaptor
    	---Purpose: ConstructionError is raised if UFirst>ULast or VFirst>VLast
    	---C++: inline
    raises ConstructionError from Standard;
    
end HCurve;
