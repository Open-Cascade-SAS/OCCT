-- Created on: 2000-09-28
-- Created by: Andrey BETENEV
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ExternFile from STEPCAFControl inherits TShared from MMgt

    ---Purpose: Auxiliary class serving as container for data resulting
    --          from translation of external file

uses
    HAsciiString from TCollection,
    ReturnStatus from IFSelect,
    WorkSession from XSControl,
    Shape from TopoDS,
    Label from TDF

is

    Create returns ExternFile;
    	---Purpose: Creates an empty structure
	
    SetWS (me: mutable; WS: WorkSession from XSControl);
    	---C++: inline
    GetWS (me) returns WorkSession from XSControl;
    	---C++: inline
    
    SetLoadStatus (me: mutable; stat: ReturnStatus from IFSelect);
    	---C++: inline
    GetLoadStatus (me) returns ReturnStatus from IFSelect;
    	---C++: inline
    
    SetTransferStatus (me: mutable; isok: Boolean);
    	---C++: inline
    GetTransferStatus (me) returns Boolean;
    	---C++: inline
    
    SetWriteStatus (me: mutable; stat: ReturnStatus from IFSelect);
    	---C++: inline
    GetWriteStatus (me) returns ReturnStatus from IFSelect;
    	---C++: inline
    
    SetName (me: mutable; name: HAsciiString from TCollection);
    	---C++: inline
    GetName (me) returns HAsciiString from TCollection;
    	---C++: inline
    
--    SetShape (me: mutable; S: Shape from TopoDS);
    	---C++: inline
--    GetShape (me) returns Shape from TopoDS;
    	---C++: inline
    
    SetLabel (me: mutable; L: Label from TDF);
    	---C++: inline
    GetLabel (me) returns Label from TDF;
    	---C++: inline
    
fields

    myWS   : WorkSession from XSControl;
    
    myLoadStatus: ReturnStatus from IFSelect;
    myTransferStatus: Boolean;
    myWriteStatus: ReturnStatus from IFSelect;

    myName: HAsciiString from TCollection;

--    myShape: Shape from TopoDS;
    myLabel: Label from TDF;

end ExternFile;
