-- Created on: 1998-04-09
-- Created by: Andre LIEUTIER
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class NLPlate from NLPlate
---Purpose: 
--
--       

uses 
     XY from gp,
     XYZ from gp, 
     StackOfPlate  from  NLPlate,
     HGPPConstraint  from  NLPlate,
     SequenceOfHGPPConstraint from  NLPlate, 
     Shape   from GeomAbs,
     Surface  from  Geom
is

    Create(InitialSurface  :  Surface  from  Geom) returns NLPlate;
-- 
-- Geometric Constraints
-- 
    Load (me : in out;  GConst : HGPPConstraint);

    Solve(me : in out; ord : Integer = 2;  InitialConsraintOrder  :  Integer=1);

    Solve2(me : in out; ord : Integer = 2;  InitialConsraintOrder  :  Integer=1);

    IncrementalSolve(me : in out; ord : Integer = 2;  InitialConsraintOrder  :  Integer=1; 
    	NbIncrements  :  Integer  =  4;  UVSliding  :  Boolean  =  Standard_False);

    IsDone(me)
        ---Purpose: returns True if all has been correctly done.
    returns Boolean;

    destroy(me : in out);
     ---C++: alias ~
 
    
    Init(me: in out );
    	---Purpose: reset the Plate in the initial state
    	--           ( same as after Create((Surface))
    
    Evaluate(me ; point2d : XY from gp )  
    returns XYZ from gp ; 
    
    EvaluateDerivative(me; point2d: XY  from gp;  
                       iu,iv  : Integer)  
    returns XYZ from gp ; 
         
    Continuity(me)  returns  Integer;

        -- private methods :
    Iterate(me : in out;  
        ConstraintOrder,  ResolutionOrder  :Integer; 
    	IncrementalLoading  : Real  =  1.0) returns Boolean
    is  private;  
     
    ConstraintsSliding(me : in out;  NbIterations  :  Integer  =  3);
    
    MaxActiveConstraintOrder(me) returns Integer;
    
    

fields 
    myInitialSurface  :  Surface  from  Geom;
    myHGPPConstraints : SequenceOfHGPPConstraint; 
    mySOP  :  StackOfPlate;
    OK : Boolean;
end;


