-- Created on: 2001-04-19
-- Created by: Peter KURNEV
-- Copyright (c) 2001-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class PointBetween from BOPTools 

    	---Purpose:  
    	--  class for storing geometry information about  
    	--  a point between neighbouring paves along 
	--  an edge 
      	--- 
uses 
    Pnt from gp
    


is 
    Create  
    	returns PointBetween from BOPTools;  
    	---Purpose:  
    	--- Empty constructor 
    	---
    SetParameter (me:out; 
    	    T:Real  from  Standard); 
    	---Purpose:  
    	--- Modifier 
    	--- sets value of the point's parameter on the edge  
    	---
    SetUV (me:out; 
    	    U:Real  from  Standard;      
    	    V:Real  from  Standard);       
    	---Purpose:  
    	--- Modifier 
    	--- sets values of the point's parameter on the face  
    	---
    SetPnt (me:out; 
    	    aP:Pnt from gp); 
    	---Purpose:  
    	--- Modifier 
    	--- sets the 3D-point   
    	---
    Parameter (me) 
    	returns Real  from  Standard ; 
    	---Purpose:  
    	--- Selector
    	---
    UV  (me; 
    	   U:out Real  from  Standard;      
    	   V:out Real  from  Standard);  
    	---Purpose:  
    	--- Selector
    	---
    Pnt (me) 
    	returns Pnt from gp; 
    	---C++:  return const &    	 
    	---Purpose:  
    	--- Selector
    	---
    
fields 
   
    myT  :  Real  from  Standard;  
    myU  :  Real  from  Standard;  
    myV  :  Real  from  Standard;  
    myPnt:  Pnt   from  gp; 
     
end PointBetween;
