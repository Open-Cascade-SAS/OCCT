-- Created on: 1998-10-15
-- Created by: Denis PASCAL
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Tool from ViewerTest

	---Purpose: to build and initialize ViewerTest static variables.
	--          ====================================================

uses Viewer             from V3d,
     InteractiveContext from AIS


is    

    MakeViewer (myclass; title : CString from Standard) 
    ---Purpose: create a new <context>. ViewerTest variables are not initialized;
    returns Viewer from V3d;

    MakeContext (myclass; title : CString from Standard) 
    ---Purpose: create a new <context>. ViewerTest variables are not initialized;
    returns InteractiveContext from AIS;
    
    InitViewerTest (myclass; current : InteractiveContext from AIS);
    ---Purpose: init variables of ViewerTest with <current>

end Tool;
