-- Created on: 1997-08-22
-- Created by: VAUTHIER Jean-Claude
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Cylinder from QANewBRepNaming inherits TopNaming from QANewBRepNaming

    ---Purpose: To load the Cylinder results

uses 
 
    MakeCylinder from BRepPrimAPI,
    Label        from TDF,
    TypeOfPrimitive3D from QANewBRepNaming

is

    Create returns Cylinder from QANewBRepNaming;

    Create(ResultLabel : Label from TDF) 
    returns Cylinder from QANewBRepNaming; 
     
    Init(me : in out; ResultLabel : Label from TDF);


    Load (me; mkCylinder : in out MakeCylinder from BRepPrimAPI; Type : TypeOfPrimitive3D from QANewBRepNaming);

    Bottom (me)
    ---Purpose: Returns the label of the bottom
    --          face of the cylinder.
    returns Label from TDF;

    Top (me)
    ---Purpose: Returns the label of the top
    --          face of the cylinder.
    returns Label from TDF;

    Lateral (me)
    ---Purpose: Returns the label of the lateral
    --          face of the cylinder.
    returns Label from TDF;

    StartSide (me)
    ---Purpose: Returns the label of the first
    --          side of the cylinder
    returns Label from TDF;
        
    EndSide (me)
    ---Purpose: Returns the label of the second
    --          side of the cylinder.
    returns Label from TDF;


end Cylinder;



