-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class OffsetCurve3d from StepGeom 

inherits Curve from StepGeom 

uses

	Real from Standard, 
	Logical from StepData, 
	Direction from StepGeom, 
	HAsciiString from TCollection
is

	Create returns mutable OffsetCurve3d;
	---Purpose: Returns a OffsetCurve3d


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aBasisCurve : mutable Curve from StepGeom;
	      aDistance : Real from Standard;
	      aSelfIntersect : Logical from StepData;
	      aRefDirection : mutable Direction from StepGeom) is virtual;

	-- Specific Methods for Field Data Access --

	SetBasisCurve(me : mutable; aBasisCurve : mutable Curve);
	BasisCurve (me) returns mutable Curve;
	SetDistance(me : mutable; aDistance : Real);
	Distance (me) returns Real;
	SetSelfIntersect(me : mutable; aSelfIntersect : Logical);
	SelfIntersect (me) returns Logical;
	SetRefDirection(me : mutable; aRefDirection : mutable Direction);
	RefDirection (me) returns mutable Direction;

fields

	basisCurve : Curve from StepGeom;
	distance : Real from Standard;
	selfIntersect : Logical from StepData;
	refDirection : Direction from StepGeom;

end OffsetCurve3d;
