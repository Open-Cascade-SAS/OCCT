-- Created on: 1994-08-25
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Modifier from BRepTools

	---Purpose: 

uses Shape               from TopoDS,
     Modification        from BRepTools,
     DataMapOfShapeShape from TopTools

raises NullObject   from Standard,
       NoSuchObject from Standard

is

    Create returns Modifier from BRepTools;
	---Purpose: Creates an empty Modifier.


    Create(S: Shape from TopoDS)
      	returns Modifier from BRepTools;
	---Purpose: Creates a modifier on the shape <S>.


    Create(S: Shape from TopoDS; M: Modification from BRepTools)
    	returns Modifier from BRepTools;
	---Purpose: Creates a modifier on  the shape <S>, and performs
	--          the modifications described by <M>.


    Init(me: in out; S: Shape from TopoDS)
    	is static;
	---Purpose: Initializes the modifier with the shape <S>.


    Perform(me: in out; M: Modification from BRepTools)
	---Purpose: Performs the modifications described by <M>.
    	raises NullObject from Standard 
        -- if the modifier has not been initialized with a shape.
    	is static;

    IsDone(me)
    
	---Purpose: Returns Standard_True if the modification has
	--          been computed successfully.
	--          
	---C++: inline
    	returns Boolean from Standard
	is static;
    

    ModifiedShape(me; S: Shape from TopoDS)
    	returns Shape from TopoDS
	---Purpose: Returns the modified shape corresponding to <S>.
	---C++: return const&
	---C++: inline
	raises NoSuchObject from Standard
               -- if S is not the initial shape or a sub-shape
               -- of the initial shape.

	is static;

		 
    -- private implementation methods

    Put(me: in out; S: Shape from TopoDS)
    
    	is static private;


    Rebuild(me: in out; S: Shape from TopoDS; M: Modification from BRepTools) 
    	returns Boolean from Standard
    	is static private;


fields

    myMap  : DataMapOfShapeShape from TopTools;
    myShape: Shape               from TopoDS;
    myDone : Boolean             from Standard;

end Modifier;
