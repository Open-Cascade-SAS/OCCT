-- File:        RWStepShape_RWDefinitionalRepresentationAndShapeRepresentation.cdl
-- Created:     Tue Jul 11 19:02:37 2000
-- Author:      Andrey BETENEV
-- Copyright:   Matra-Datavision 2000

class RWDefinitionalRepresentationAndShapeRepresentation from RWStepShape

	---Purpose : Read & Write Module for ConversionBasedUnitAndLengthUnit

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     DefinitionalRepresentationAndShapeRepresentation from StepShape,
     EntityIterator from Interface

is

	Create returns RWDefinitionalRepresentationAndShapeRepresentation;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable DefinitionalRepresentationAndShapeRepresentation from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : DefinitionalRepresentationAndShapeRepresentation from StepShape);

	Share(me; ent : DefinitionalRepresentationAndShapeRepresentation from StepShape; iter : in out EntityIterator);

end RWDefinitionalRepresentationAndShapeRepresentation;
