-- Created on: 1991-06-25
-- Created by: Christophe MARION
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package BRepTest 

	---Purpose: Provides commands to test BRep.
	--          
uses
    Draw,
    TCollection
    
is
   	
    AllCommands(DI : in out Interpretor from Draw);
	---Purpose: Defines all the topology commands.

    BasicCommands(DI : in out Interpretor from Draw);
	---Purpose: Defines the basic commands.

    CurveCommands(DI : in out Interpretor from Draw);
	---Purpose: Defines the commands to build edges and wires.
	
    Fillet2DCommands(DI : in out Interpretor from Draw);
	---Purpose:  Defines the  commands  to perform add  fillets on
	--          wires and  edges.
   
    SurfaceCommands(DI : in out Interpretor from Draw);
	---Purpose: Defines the commands to build faces and shells.

    PrimitiveCommands(DI : in out Interpretor from Draw);
	---Purpose: Defines the commands to build primitives.
	
    FillingCommands(DI : in out Interpretor from Draw);
	---Purpose: Defines the commands to build primitives.
	
    SweepCommands(DI : in out Interpretor from Draw);
	---Purpose: Defines the commands to sweep shapes.
	
    TopologyCommands(DI : in out Interpretor from Draw);
	---Purpose: Defines  the    commands   to perform  topological
	--          operations. 

    FilletCommands(DI : in out Interpretor from Draw);
	---Purpose: Defines  the commands  to perform  add  fillets on
	--          shells.
   
    ChamferCommands(DI : in out Interpretor from Draw);
	---Purpose: Defines  the commands  to perform  add chamfers on
	--          shells.
	
    GPropCommands(DI : in out Interpretor from Draw);
	---Purpose: Defines commands to compute global properties.
	
    MatCommands(DI : in out Interpretor from Draw);
    	---Purpose: Defines commands to compute and to explore the map of the
    	--          Bisecting locus.


    DraftAngleCommands(DI : in out Interpretor from Draw);
	---Purpose: Defines the commands to modify draft angles of the
	--          faces of a shape.


    FeatureCommands(DI : in out Interpretor from Draw);
	---Purpose: Defines the commands to create features on a shape.


    OtherCommands(DI : in out Interpretor from Draw);
	---Purpose: Defines the auxiliary topology commands.
	

    ExtremaCommands(DI : in out Interpretor from Draw);
	---Purpose: Defines the extrema commands.
	

    CheckCommands(DI : in out Interpretor from Draw);
	---Purpose: Defines the checkshape command.

    PlacementCommands(DI : in out Interpretor from Draw);
	---Purpose: Defines the placement  command.
	--          

    ProjectionCommands(DI : in out Interpretor from Draw);
	---Purpose: Defines the commands to project a wire on a shape.
	--          

end BRepTest;

