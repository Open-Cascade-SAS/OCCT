-- Created on: 2003-08-29
-- Created by: data exchange team
-- Copyright (c) 2003-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ShapeMapTool from XCAFDoc inherits Attribute from TDF
    ---Purpose: attribute containing map of sub shapes

uses

    SequenceOfHAsciiString from TColStd,
    Shape from TopoDS,
    IndexedMapOfShape from TopTools,
    Label from TDF,
    RelocationTable from TDF
    
is
    GetID (myclass)   
    ---C++: return const &  
    returns GUID from Standard;    


    Set (myclass; L : Label from TDF) returns ShapeMapTool from XCAFDoc;
    ---Purpose: Create (if not exist) ShapeTool from XCAFDoc on <L>.


    Create returns ShapeMapTool from XCAFDoc;
    	---Purpose: Creates an empty tool
    
    
    ---API: Analysis

    
    IsSubShape (me; sub: Shape from TopoDS) 
    returns Boolean;
    	---Purpose: Checks whether shape <sub> is subshape of shape stored on
        --          label shapeL

    SetShape (me: mutable; S: Shape from TopoDS);
    	---Purpose: Sets representation (TopoDS_Shape) for top-level shape

            ---Category: TDF_Attribute methods
    --           =====================
    
    ID (me)
    	---C++: return const & 
    returns GUID from Standard;

    Restore (me: mutable; with : Attribute from TDF);

    NewEmpty (me)
    returns Attribute from TDF;

    Paste (me; into : Attribute from TDF;
	       RT   : RelocationTable from TDF);    

    GetMap (me) returns IndexedMapOfShape from TopTools;
    ---C++: return const & 

fields

    myMap: IndexedMapOfShape from TopTools;
    
end ShapeTool;
