-- Created on: 1999-04-14
-- Created by: Roman LYGIN
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SplitSurfaceContinuity from ShapeUpgrade inherits SplitSurface from ShapeUpgrade

    ---Purpose: Splits a Surface with a continuity criterion.
    --          At the present moment C1 criterion is used only.
    --          This tool works with tolerance. If C0 surface can be corrected
    --          at a knot with given tolerance then the surface is corrected,
    --          otherwise it is spltted at that knot.

uses

    Shape from GeomAbs

is

    Create returns SplitSurfaceContinuity from ShapeUpgrade; 
        ---Purpose: Empty constructor.
	
    SetCriterion (me: mutable; Criterion: Shape from GeomAbs);
    	---Purpose: Sets criterion for splitting.
	
    SetTolerance (me: mutable; Tol: Real);
    	---Purpose: Sets tolerance.
	
    --Build (me: mutable; Segment: Boolean) is redefined;
    	--Purpose: Performs correction/splitting of the supporting surface(s).
	---         First defines splitting values, then calls inherited method.
    Compute(me: mutable; Segment: Boolean) is redefined;
    --Perform(me: mutable; Segment: Boolean);
fields

    myCriterion: Shape from GeomAbs;
    myTolerance: Real;
    myCont     : Integer;
    
end SplitSurfaceContinuity;
