-- File:	Box2d.cdl
-- Created:	Mon Jan 28 11:51:08 1991
-- Author:	Remi Lequette
--		<rle@topsn3>
---Copyright:	 Matra Datavision 1991, 1992


class Box2d from Bnd 

	---Purpose: Describes a bounding box in 2D space.
    	-- A bounding box is parallel to the axes of the coordinates
    	-- system. If it is finite, it is defined by the two intervals:
    	-- -   [ Xmin,Xmax ], and
    	-- -   [ Ymin,Ymax ].
    	-- A bounding box may be infinite (i.e. open) in one or more
    	-- directions. It is said to be:
    	-- -   OpenXmin if it is infinite on the negative side of the   "X Direction";
    	-- -   OpenXmax if it is infinite on the positive side of the   "X Direction";
    	-- -   OpenYmin if it is infinite on the negative side of the   "Y Direction";
    	-- -   OpenYmax if it is infinite on the positive side of the   "Y Direction";
    	-- -   WholeSpace if it is infinite in all four directions. In
    	--   this case, any point of the space is inside the box;
    	-- -   Void if it is empty. In this case, there is no point included in the box.
    	--  A bounding box is defined by four bounds (Xmin, Xmax, Ymin and Ymax) which
    	--   limit the bounding box if it is finite, six flags (OpenXmin, OpenXmax, OpenYmin,
    	--   OpenYmax, WholeSpace and Void) which describe the bounding box if it is infinite or empty, and
    	-- -   a gap, which is included on both sides in any direction when consulting the finite bounds of the box.


uses    Pnt2d  from gp,
    	Dir2d  from gp,
    	Lin2d  from gp,
    	Trsf2d from gp
    
raises
    ConstructionError from Standard

is

    Create returns Box2d from Bnd;
	---Purpose: Creates an empty 2D bounding box.
    	-- The constructed box is qualified Void. Its gap is null.
	---C++: inline

    SetWhole(me : in out)    is static;
	---Purpose: Sets this bounding box so that it covers the whole 2D
    	-- space, i.e. it is infinite in all directions.
    	---C++: inline

    SetVoid(me : in out)    is static;
	---Purpose: Sets this 2D bounding box so that it is empty. All points are outside a void box.
    	---C++: inline

    Set(me : in out; P : Pnt2d)    is static;
	---Purpose: Sets this 2D bounding box so that it bounds
    	--   the point P. This involves first setting this bounding box
    	--   to be void and then adding the point PThe rectangle bounds   the  point <P>.   
	---C++: inline

    Set(me : in out; P : Pnt2d; D : Dir2d)    is static;
	---Purpose: Sets this 2D bounding box so that it bounds
    	-- the half-line defined by point P and direction D, i.e. all
    	--   points M defined by M=P+u*D, where u is greater than
    	--   or equal to 0, are inside the bounding area. This involves
    	--   first setting this 2D box to be void and then adding the   half-line.
	---C++: inline

    Update(me : in out; aXmin, aYmin, aXmax, aYmax : Real)
	---Purpose: Enlarges this 2D bounding box, if required, so that it
    	--          contains at least:
    	--   -   interval [ aXmin,aXmax ] in the "X Direction",
    	--   -   interval [ aYmin,aYmax ] in the "Y Direction"
    is static;

    Update(me : in out; X,Y : Real)
	---Purpose:    Adds a point of coordinates (X,Y) to this bounding box.
    is static;

    GetGap(me) returns Real
	---Purpose: Returns the gap of this 2D bounding box.
 	---C++: inline
    is static;

    SetGap(me : in out; Tol : Real)
	---Purpose: Set the gap of this 2D bounding box to abs(Tol).
	---C++: inline
    is static;

    Enlarge(me : in out; Tol : Real)
	---Purpose: Enlarges     the  box  with    a  tolerance  value.
	--   This means that the minimum values of its X and Y
    	-- intervals of definition, when they are finite, are reduced by
    	-- the absolute value of Tol, while the maximum values are
    	-- increased by the same amount.
  	---C++: inline
    is static;

    Get(me; aXmin, aYmin, aXmax, aYmax : out Real)
	---Purpose: Returns the bounds of this 2D bounding box. 
    	-- The gap is included. If this bounding box is infinite (i.e. "open"), returned values
    	-- may be equal to +/- Precision::Infinite().
    raises ConstructionError -- if IsVoid()
    is static;
    
    OpenXmin(me : in out)
	---Purpose: The Box will be infinitely long in the Xmin direction.
	---Level: Public 
	---C++: inline
    is static;
    
    OpenXmax(me : in out)
	---Purpose: The Box will be infinitely long in the Xmax direction.
	---Level: Public 
	---C++: inline
    is static;
    
    OpenYmin(me : in out)
	---Purpose: The Box will be infinitely long in the Ymin direction.
	---Level: Public 
	---C++: inline
    is static;
    
    OpenYmax(me : in out)
	---Purpose: The Box will be infinitely long in the Ymax direction.
	---Level: Public 
	---C++: inline
    is static;
    
    IsOpenXmin(me) returns Boolean
	---Purpose: Returns true if this bounding box is open in the Xmin direction.
  	---C++: inline
    is static;
    
    IsOpenXmax(me) returns Boolean
	---Purpose: Returns true if this bounding box is open in the Xmax direction.
  	---C++: inline
    is static;
    
    IsOpenYmin(me) returns Boolean
	---Purpose: Returns true if this bounding box is open in the Ymin direction.
  	---C++: inline
    is static;
    
    IsOpenYmax(me) returns Boolean
	---Purpose: Returns true if this bounding box is open in the Ymax direction.
  	---C++: inline
    is static;
    
    IsWhole(me) returns Boolean    is static;
	---Purpose:
    	-- Returns true if this bounding box is infinite in all 4
    	-- directions (Whole Space flag).
   	---C++: inline
 
    IsVoid(me) returns Boolean    is static;
	---Purpose:
    	-- Returns true if this 2D bounding box is empty (Void flag).
    	---C++: inline

    Transformed(me; T : Trsf2d from gp)
	---Purpose: Returns a bounding box which is the result of applying the
    	-- transformation T to this bounding box.
    	-- Warning
    	-- Applying a geometric transformation (for example, a
    	-- rotation) to a bounding box generally increases its
    	-- dimensions. This is not optimal for algorithms which use it.
    
    returns Box2d from Bnd    is static;

    Add(me : in out; Other : Box2d)    is static;
	---Purpose: Adds the 2d box <Other> to <me>.
	---Level: Public 
    
    Add(me : in out; P : Pnt2d)    is static;
	---Purpose: Adds  the 2d pnt <P> to <me>.
	---Level: Public 
	---C++: inline

    Add(me : in out; P : Pnt2d; D : Dir2d)    is static;
	---Purpose: Extends <me> from the Pnt <P> in the direction <D>.
	---Level: Public 
	---C++: inline
    
    Add(me : in out; D : Dir2d)    is static;
	---Purpose: Extends the Box  in the given Direction, i.e. adds
	--          a half-line. The box may become infinite in 1 or 2
	--          directions. 
	---Level: Public 
    
    IsOut(me; P : Pnt2d) returns Boolean    is static;
	---Purpose: Returns True if the 2d pnt <P> is out <me>.
	---Level: Public 
    
    IsOut(me; Other : Box2d) returns Boolean    is static;
	---Purpose: Returns True if <Box2d> is out <me>.
	---Level: Public 

    IsOut(me; Other : Box2d; T : Trsf2d from gp) returns Boolean    is static;
	---Purpose: Returns True if transformed <Box2d> is out <me>.
	---Level: Public 
	---C++: inline

    IsOut(me; T1 : Trsf2d from gp; Other : Box2d; T2 : Trsf2d from gp)
    returns Boolean    is static;
	---Purpose: Compares  a transformed  bounding with  a    transformed
	--          bounding. The default implementation is  to make a copy
	--          of <me> and <Other>, to transform them and to test.
	---Level: Public 
	---C++: inline

    Dump(me)    is static;


fields  Xmin : Real; 
    	Xmax : Real; 
    	Ymin : Real; 
    	Ymax : Real; 
	Gap  : Real;
    	Flags : Integer;  -- 6 flags

end Box2d;
