-- Created on: 1992-08-26
-- Created by: Jean Louis FRENKEL
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package StdPrs
    	---Purpose: The StdPrs package provides standard display tools
	-- for specific geometries and topologies whereas
	-- Prs3d provides those for generic objects. Among
	-- these classes are definitions of the display of the
	-- specific geometry or topology in various display
	-- modes such as wireframe, shading or hidden line removal mode.
    	       
uses
  Prs3d,
	Geom,
	Geom2d,
	Adaptor3d,
	Adaptor2d,
  GeomAdaptor,
	Geom2dAdaptor,
  BRepAdaptor,
	TopTools,
	TopoDS,
	TopExp,
  TopAbs,
	BRepTools,
	Bnd,
  TColStd,
  HLRAlgo,
  HLRBRep,
  Quantity,
	BRepMesh,
	gp,
	TColgp,
	Poly,
	TopLoc, 
	Graphic3d

is
   class ToolPoint;
   class ToolVertex;
   class ToolRFace;
   class HLRToolShape;
   class ToolShadedShape;
   class ShadedShape;
    
   class PoleCurve;

   class Plane;

   class WFPoleSurface;

   class DeflectionCurve;		      

	---Category: Wireframe algorithms
   
   class WFDeflectionSurface;

   class ShadedSurface;

   -----------------------------------------------
   --- deflection drawing classes :
   -----------------------------------------------

   class WFDeflectionRestrictedFace;

   class Curve;

   class WFSurface;

   ---Category: Hidden lines removal algorithms.
   
   class HLRPolyShape; 

   imported HLRShape;

   imported NListOfSequenceOfPnt from Prs3d; 
   imported NListIteratorOfListOfSequenceOfPnt from Prs3d;
   
   imported WFShape;
   imported WFDeflectionShape;

   imported Vertex;
   imported Point;

   imported WFRestrictedFace;

end StdPrs;



