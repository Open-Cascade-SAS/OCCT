-- Created on: 1994-04-01
-- Created by: Yves FRICAUD
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PolyBis from Bisector 

	---Purpose: Polygon of PointOnBis

uses
    PointOnBis from Bisector,
    Trsf2d     from gp

is
    Create returns PolyBis from Bisector;
    
    Append ( me : in out; Point : PointOnBis from Bisector) 
    is static ;
						    		
    Length (me) returns Integer
    is static ;
    
    IsEmpty (me) returns Boolean
    is static;

    Value (me ; Index : Integer) returns PointOnBis from Bisector
       ---C++: return const&
    is static;
    
    First (me) returns PointOnBis from Bisector
       ---C++: return const&
    is static;
    
    Last (me) returns PointOnBis from Bisector
       ---C++: return const&
    is static;
    
    Interval (me ; U :Real) returns Integer from Standard
    is static;
    
    Transform (me : in out ; T :Trsf2d)
    is static;
    
fields

    thePoints       : PointOnBis from Bisector [30];
    nbPoints        : Integer    from Standard;
    
end PolyBis;

