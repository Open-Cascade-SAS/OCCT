-- Created on: 1991-12-06
-- Created by: Remi LEQUETTE
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package HLRTest 

	---Purpose: This package   is  a test  of  the    Hidden Lines
	--          algorithms instantiated on the BRep Data Structure
	--          and using the Draw package to display the results.

uses
    Standard,
    MMgt,
    TCollection,
    gp,
    TopoDS,
    HLRAlgo,
    HLRBRep,
    HLRTopoBRep,
    Draw

is
    class ShapeData;
    
    class DrawableEdgeTool;
	---Purpose: Used to display the results.

    class DrawablePolyEdgeTool;
	---Purpose: Used to display the results.

    class Projector;
	---Purpose: Draw Variable Projector to test
	
    class OutLiner;
	---Purpose: Draw Variable Outliner to test

    Set(Name : CString;
        P    : Projector from HLRAlgo);
	---Purpose: Set a Projector Variable

    GetProjector(Name : in out CString;
                 P :    in out Projector from HLRAlgo) 
    returns Boolean; 
	---Purpose: Get a projector variable
	--          Returns false if the variable is not a projector

    Set(Name : CString;
        S    : Shape from TopoDS);
	---Purpose: Set a OutLiner Variable

    GetOutLiner(Name : in out CString)  
    	returns OutLiner from HLRTopoBRep;
	---Purpose: Get a outliner variable
	--          Returns a null handle if the variable is not a outliner

    Commands(I : in out Interpretor from Draw);
	---Purpose: Defines commands to test the Hidden Line Removal

end HLRTest;
