-- Created on: 1993-09-28
-- Created by: Bruno DUMORTIER
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Curved from GeomFill inherits Filling from GeomFill

uses
    Array1OfPnt  from TColgp,
    Array1OfReal from TColStd

is
    Create;
    
    Create(P1, P2, P3, P4 : Array1OfPnt from TColgp)
    returns Curved from GeomFill;
    
    Create(P1, P2, P3, P4 : Array1OfPnt  from TColgp;
    	   W1, W2, W3, W4 : Array1OfReal from TColStd)
    returns Curved from GeomFill;
    

    Create(P1, P2, P3 : Array1OfPnt from TColgp)
    returns Curved from GeomFill;
    
    Create(P1, P2, P3 : Array1OfPnt  from TColgp;
    	   W1, W2, W3 : Array1OfReal from TColStd)
    returns Curved from GeomFill;
    

    Create(P1, P2 : Array1OfPnt from TColgp)
    returns Curved from GeomFill;
    
    Create(P1, P2 : Array1OfPnt  from TColgp;
    	   W1, W2 : Array1OfReal from TColStd)
    returns Curved from GeomFill;
    

    Init(me : in out;
    	 P1, P2, P3, P4 : Array1OfPnt from TColgp)
    is static;

    Init(me : in out;
    	 P1, P2, P3, P4 : Array1OfPnt  from TColgp;
    	 W1, W2, W3, W4 : Array1OfReal from TColStd)
    is static;

    Init(me : in out;
    	 P1, P2, P3 : Array1OfPnt from TColgp)
    is static;

    Init(me : in out;
    	 P1, P2, P3 : Array1OfPnt  from TColgp;
    	 W1, W2, W3 : Array1OfReal from TColStd)
    is static;

    Init(me : in out;
    	 P1, P2 : Array1OfPnt from TColgp)
    is static;

    Init(me : in out;
    	 P1, P2 : Array1OfPnt  from TColgp;
    	 W1, W2 : Array1OfReal from TColStd)
    is static;

end Curved;
