-- Created on: 1998-06-03
-- Created by: data exchange team
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Wire from ShapeAnalysis inherits TShared from MMgt

	---Purpose: This class provides analysis of a wire to be compliant to 
    	--          CAS.CADE requirements.
    	--
   	--	    The functionalities provided are the following:
    	--	     1. consistency of 2d and 3d edge curve senses
    	--           2. connection of adjacent edges regarding to: 
    	--	       a. their vertices 
    	--	       b. their pcurves 
    	--	       c. their 3d curves 
    	--           3. adjacency of the edge vertices to its pcurve and 3d curve 
    	--	     4. if a wire is closed or not (considering its 3d and 2d 
    	--              contour) 
    	--	     5. if a wire is outer on its face (considering pcurves)
    	--
    	--
    	-- 	    This class can be used in conjunction with class 
    	--	    ShapeFix_Wire, which will fix the problems detected by this class.
    	--
    	--          The methods of the given class match to ones of the class 
    	--	    ShapeFix_Wire, e.g., CheckSmall and FixSmall. 
    	--          This class also includes some auxilary methods 
    	--          (e.g., CheckOuterBound, etc.),
    	--          which have no pair in ShapeFix_Wire.
    	--
    	--          Like methods of ShapeFix_Wire the ones of this class are 
    	-- 	    grouped into two levels:
    	--          - Public which are recommended for use (the most global 
    	--	      method is Perform),
    	--	    - Advanced, for optional use only
    	--
    	--          For analyzing result of Public API checking methods use
    	--          corresponding Status... method. 
    	--          The 'advanced' functions share the single status field which 
    	--          contains the result of the last performed 'advanced' method. 
    	--          It is quried by the method LastCheckStatus().
	--
	--          In order to prepare an analyzer, it is necessary to load a wire, 
        --          set face and precision.

uses

    Pnt2d     from gp,
    Curve     from Geom2d,
    Surface   from Geom,
    Location  from TopLoc,
    Shape     from TopoDS,
    Wire      from TopoDS,
    Face      from TopoDS,
    SequenceOfIntersectionPoint from IntRes2d,
    SequenceOfPnt               from TColgp,
    SequenceOfReal              from TColStd,
    Status    from ShapeExtend,
    WireData  from ShapeExtend,
    WireOrder from ShapeAnalysis,
    Surface   from ShapeAnalysis,
    IndexedMapOfShape from TopTools,
    DataMapOfShapeListOfShape from TopTools,
    MapOfShape from TopTools
is

    Create returns Wire from ShapeAnalysis;
    	---Purpose: Empty constructor
    
    Create (wire     : Wire from TopoDS;
    	    face     : Face from TopoDS;
    	    precision: Real)
    returns Wire from ShapeAnalysis;
    	---Purpose: Creates object with standard TopoDS_Wire, face
	--          and precision
    
    Create (sbwd     : WireData from ShapeExtend;
    	    face     : Face from TopoDS;
    	    precision: Real)
    returns Wire from ShapeAnalysis;
    	---Purpose: Creates the object with WireData object, face
	--          and precision
	
    Init (me: mutable; wire     : Wire from TopoDS;
    	              face     : Face from TopoDS;
    	              precision: Real);
    	---Purpose: Initializes the object with standard TopoDS_Wire, face
	--          and precision
    
    Init (me: mutable; sbwd     : WireData from ShapeExtend;
    	              face     : Face from TopoDS;
    	              precision: Real);
    	---Purpose: Initializes the object with WireData object, face
	--          and precision
	
    Load (me: mutable; wire: Wire from TopoDS);
    	---Purpose: Loads the object with standard TopoDS_Wire

    Load (me: mutable; sbwd: WireData from ShapeExtend);
    	---Purpose: Loads the object with WireData object
	---Remark : Single WireData object will be shared

    SetFace (me: mutable; face : Face from TopoDS);
    	---Purpose: Loads the face the wire lies on

    SetSurface (me: mutable; surface : Surface from Geom);
    	---Purpose: Loads the surface the wire lies on

    SetSurface (me: mutable; surface : Surface from Geom;
    	    	    	    location: Location from TopLoc);
    	---Purpose: Loads the surface the wire lies on

    SetPrecision (me: mutable; precision: Real);
    	---Precision: Set the precision value

    ClearStatuses (me: mutable);
    	---Purpose: Unsets all the status and distance fields
	--          wire, face and precision are not cleared

    IsLoaded (me) returns Boolean;
        ---C++: inline
    	---Purpose: Returns True if wire is loaded and has number of edges >0
 	
    IsReady (me) returns Boolean;
        ---C++: inline
    	---Purpose: Returns True if IsLoaded and underlying face is not null
	
    Precision (me) returns Real;
        ---C++: inline
    	---Purpose: Returns the value of precision
    
    WireData (me) returns WireData from ShapeExtend;
    	---C++: return const &
        ---C++: inline
    	---Purpose: Returns wire object being analyzed
	
    NbEdges (me) returns Integer;
        ---C++: inline
    	---Purpose: Returns the number of edges in the wire, or 0 if it is not loaded

    Face (me) returns Face from TopoDS;
    	---C++: return const &
        ---C++: inline
    	---Purpose: Returns the working face

    Surface (me) returns Surface from ShapeAnalysis;
    	---C++: return const &
        ---C++: inline
    	---Purpose: Returns the working surface
        
    
    ---Checking methods:
    
    ---Level: Public
    
    ---Return: Check..() methods return True when and only when the situation was
    --         analyzed and the specific case detected. 
    --         This corresponds to the flag DONE (or one of DONE#i) set in Status.

    Perform (me : mutable) returns Boolean; 
    	---Purpose: Performs all the checks in the following order :
    	--	    CheckOrder, CheckSmall, CheckConected, CheckEdgeCurves,
    	--          CheckDegenerated, CheckSelfIntersection, CheckLacking,
    	--          CheckClosed
    	--  Returns: True if at least one method returned True;
    	--          For deeper analysis use Status...(status) methods
    
    CheckOrder (me: mutable; isClosed: Boolean = Standard_True;
    	    	    	     mode3d: Boolean = Standard_True) returns Boolean;
    	---Purpose: Calls CheckOrder and returns False if wire is already
	--          ordered (tail-to-head), True otherwise
	--          Flag <isClosed> defines if the wire is closed or not
	--          Flag <mode3d> defines which mode is used (3d or 2d)
	
    CheckConnected (me : mutable; prec : Real = 0.0) returns Boolean;
    	---Purpose: Calls to CheckConnected for each edge
    	--  Returns: True if at least one pair of disconnected edges (not sharing the 
    	-- 	    same vertex) was detected
    
    CheckSmall (me : mutable; precsmall : Real = 0.0) returns Boolean;
    	---Purpose: Calls to CheckSmall for each edge
    	--  Returns: True if at least one small edge was detected
    
    CheckEdgeCurves (me : mutable) returns Boolean;
    	---Purpose: Checks edges geometry (consitency of 2d and 3d senses, adjasment 
    	--	    of curves to the vertices, etc.).
    	--	    The order of the checks :
	--          Call ShapeAnalysis_Wire to check:
    	--	    ShapeAnalysis_Edge::CheckCurve3dWithPCurve  (1),
        --          ShapeAnalysis_Edge::CheckVertcesWithPCurve  (2), 
    	--	    ShapeAnalysis_Edge::CheckVertcesWithCurve3d (3),
	--          CheckSeam                                   (4)
	--          Additional:
        --          CheckGap3d                                  (5),
	--          CheckGap2d                                  (6),
    	--          ShapeAnalysis_Edge::CheckSameParameter      (7)
    	-- Returns: True if at least one check returned True
	--  Remark:  The numbers in brackets show with what DONEi or FAILi
	--          the status can be queried
    
    CheckDegenerated (me : mutable) returns Boolean;
    	---Purpose: Calls to CheckDegenerated for each edge
    	--  Returns: True if at least one incorrect degenerated edge was detected
    
    CheckClosed (me : mutable; prec : Real = 0.0) returns Boolean;
    	---Purpose: Checks if wire is closed, performs CheckConnected, 
    	--          CheckDegenerated and CheckLacking for the first and the last edges
    	--  Returns: True if at least one check returned True
	--  Status:
    	--          FAIL1 or DONE1: see CheckConnected
	--          FAIL2 or DONE2: see CheckDegenerated

    CheckSelfIntersection (me : mutable) returns Boolean;
    	---Purpose: Checks self-intersection of the wire (considering pcurves)
    	--          Looks for self-intersecting edges and each pair of intersecting 
    	--          edges.
    	--  Warning: It does not check each edge with any other one (only each two 
    	--          adjacent edges)
    	--          The order of the checks :
    	--          CheckSelfIntersectingEdge, CheckIntersectingEdges
    	--  Returns: True if at least one check returned True
	--  Status:  FAIL1 or DONE1 - see CheckSelfIntersectingEdge
	--          FAIL2 or DONE2 - see CheckIntersectingEdges
    
    CheckLacking (me : mutable) returns Boolean;
    	---Purpose: Calls to CheckLacking for each edge
    	--  Returns: True if at least one lacking edge was detected
    
    CheckGaps3d (me : mutable) returns Boolean;
    	---Purpose: 
    	---Returns: 

    CheckGaps2d (me : mutable) returns Boolean;
    	---Purpose: 
    	---Returns: 

    CheckCurveGaps (me : mutable) returns Boolean;
    	---Purpose: 
    	---Returns: 


    ---Level: Advanced

    ---Status: For analyzing the status of the last performed method use method
    --          Status(status)
    --
    --          All the Check...() methods below return False if the problem was 
    --          not detected. If so, Status(ShapeExtend_OK) returns True.
    
    CheckOrder (me: mutable; sawo: out WireOrder from ShapeAnalysis;
    	    	    	     isClosed: Boolean = Standard_True;
    	    	    	     mode3d: Boolean = Standard_True)
    returns Boolean;
    	---Purpose: Analyzes the order of the edges in the wire,
	--          uses class WireOrder for that purpose.
	--          Flag <isClosed> defines if the wire is closed or not
	--          Flag <mode3d> defines which mode is used (3d or 2d)
    	--          Returns False if wire is already ordered (tail-to-head),
    	--          True otherwise.
	--          Use returned WireOrder object for deeper analysis.
	--  Status:
	--          OK   : the same edges orientation, the same edges sequence
        --          DONE1: the same edges orientation, not the same edges sequence
	--          DONE2: as DONE1 and gaps more than myPrecision
	--          DONE3: not the same edges orientation (some need to be reversed)
	--          DONE4: as DONE3 and gaps more than myPrecision
	--          FAIL : algorithm failed (could not detect order)

    CheckConnected (me : mutable; num: Integer; prec: Real = 0.0) returns Boolean;
    	---Purpose: Checks connected edges (num-th and preceeding).
    	--           Tests with starting preci from <SBWD> or  with <prec> if  
    	--	         it is greater.
    	--           Considers Vertices.
    	--  Returns: False if edges are connected by the common vertex, else True
    	--  Status  :
    	-- 	     OK    : Vertices (end of num-1 th edge and start on num-th one) 
    	--                   are already the same
    	--           DONE1 : Absolutely confused (gp::Resolution)
    	--           DONE2 : Confused at starting <preci> from <SBWD>
    	--           DONE3 : Confused at <prec> but not <preci>
    	--           FAIL1 : Not confused
    	--           FAIL2 : Not confused but confused with <preci> if reverse num-th edge
    
    CheckSmall (me : mutable; num      : Integer;
    	    	             precsmall: Real = 0.0)
    returns Boolean;
    	---Purpose: Checks if an edge has a length not greater than myPreci or 
    	--	    precsmall (if it is smaller)
    	--  Returns: False if its length is greater than precision
	--  Status:
	--          OK   : edge is not small or degenerated
	--          DONE1: edge is small, vertices are the same
	--          DONE2: edge is small, vertices are not the same
    	--          FAIL : no 3d curve and pcurve

    CheckSeam (me : mutable; num   : Integer;
    	    	    	    C1, C2: out Curve from Geom2d;
    	    	    	    cf, cl: out Real)
    returns Boolean;
    	---Purpose: Checks if a seam pcurves are correct oriented
    	--  Returns: False (status OK) if given edge is not a seam or if it is OK
	--          C1 - current pcurve for FORWARD edge,
    	--          C2 - current pcurve for REVERSED edge (if returns True they
    	--          should be swapped for the seam),
	--          cf, cl - first and last parameters on curves
    	--  Status: 
    	--          OK   : Pcurves are correct or edge is not seam
    	--          DONE : Seam pcurves should be swapped

    CheckSeam (me : mutable; num: Integer) returns Boolean;
    	---Purpose: Checks if a seam pcurves are correct oriented
	--          See previous functions for details

    CheckDegenerated (me: mutable; num: Integer; dgnr1, dgnr2: out Pnt2d from gp)
    returns Boolean;
    	---Purpose: Checks for degenerated edge between two adjacent ones.
    	--	    Fills parameters dgnr1 and dgnr2 with points in paramterical
    	--          space that correspond to the singularity (either gap that
    	--          needs to be filled by degenerated edge or that already filled)
	--  Returns: False if no singularity or edge is already degenerated,
	--          otherwise True
    	--  Status:
    	--          OK   : No surface singularity, or edge is already degenerated
    	--	    DONE1: Degenerated edge should be inserted (gap in 2D)
    	--          DONE2: Edge <num> should be made degenerated (recompute pcurve 
    	--                 and set the flag)
	--          FAIL1: One of edges neighbouring to degenerated one has 
        --                 no pcurve
	--          FAIL2: Edge marked as degenerated and has no pcurve 
        --                 but singularity is not detected

    CheckDegenerated (me: mutable; num: Integer)
    returns Boolean;
    	---Purpose: Checks for degenerated edge between two adjacent ones.
	--  Remark : Calls previous function
    	--  Status : See the function above for details

    CheckGap3d (me : mutable; num : Integer = 0) returns Boolean;
    	---Purpose: Checks gap between edges in 3D (3d curves).
    	--          Checks the distance between ends of 3d curves of the num-th 
    	--          and preceeding edge. 
    	--	    The distance can be queried by MinDistance3d. 
    	--
    	--  Returns: True if status is DONE
    	--  Status:
    	--	    OK   : Gap is less than myPrecision
    	--          DONE : Gap is greater than myPrecision
    	--          FAIL : No 3d curve(s) on the edge(s)

    CheckGap2d (me : mutable; num : Integer = 0) returns Boolean;
    	---Purpose: Checks gap between edges in 2D (pcurves). 
    	--          Checks the distance between ends of pcurves of the num-th 
    	--          and preceeding edge. 
    	--	    The distance can be queried by MinDistance2d.
    	--         
    	--  Returns: True if status is DONE
    	--  Status:
    	--          OK   : Gap is less than parametric precision out of myPrecision
    	--          DONE : Gap is greater than parametric precision out of myPrecision
    	--          FAIL : No pcurve(s) on the edge(s)

    CheckCurveGap (me : mutable; num : Integer = 0) returns Boolean;
    	---Purpose: Checks gap between points on 3D curve and points on surface
    	--          generated by pcurve of the num-th edge.
    	--	    The distance can be queried by MinDistance3d.
    	--
    	--  Returns: True if status is DONE
    	--  Status:
    	--	    OK   : Gap is less than myPrecision
    	--          DONE : Gap is greater than myPrecision
    	--          FAIL : No 3d curve(s) on the edge(s)
     
    CheckSelfIntersectingEdge (me: mutable; num: Integer;
    	    	    	       points2d: out SequenceOfIntersectionPoint from IntRes2d;
    	    	    	       points3d: out SequenceOfPnt from TColgp)
    returns Boolean;
    	---Purpose: Checks if num-th edge is self-intersecting.
	--          Self-intersection is reported only if intersection point lies outside
	--          of both end vertices of the edge.
    	--  Returns: True if edge is self-intersecting.
    	--	    If returns True it also fills the sequences of intersection points
	--          and corresponding 3d points (only that are not enclosed by a vertices)
    	--  Status:
    	--          FAIL1 : No pcurve
    	--          FAIL2 : No vertices
    	--          DONE1 : Self-intersection found
    
    CheckSelfIntersectingEdge (me: mutable; num: Integer)
    returns Boolean;
    	--  Purpose: Checks num-th edge to be self-intersecting.
	--  Remark : Calls the previous method
    	--  Status : See the function above for details
    
    CheckIntersectingEdges (me : mutable; num: Integer;
    	    	            points2d: out SequenceOfIntersectionPoint from IntRes2d;
    	    	            points3d: out SequenceOfPnt from TColgp;
    	    	            errors: out SequenceOfReal from TColStd)
    returns Boolean;
    	---Purpose: Checks two adjacent edges for intersecting.
	--          Intersection is reported only if intersection point is not enclosed
	--          by the common end vertex of the edges.
    	--  Returns: True if intersection is found.
    	--	    If returns True it also fills the sequences of intersection points,
	--          corresponding 3d points, and errors for them (half-distances between
        --          intersection points in 3d calculated from one and from another edge)
    	--  Status:
    	--          FAIL1 : No pcurve
    	--          FAIL2 : No vertices
    	--          DONE1 : Self-intersection found
     
    CheckIntersectingEdges (me: mutable; num: Integer)
    returns Boolean;
    	---Purpose: Checks two adjacent edges for intersecting.
	--  Remark : Calls the previous method
    	--  Status : See the function above for details
    
    CheckIntersectingEdges(me: mutable; num1: Integer; num2: Integer;
    	    	    	   points2d: out SequenceOfIntersectionPoint from IntRes2d;
    	    	           points3d: out SequenceOfPnt from TColgp;
    	    	           errors: out SequenceOfReal from TColStd)
    returns Boolean;
    	---Purpose: Checks i-th and j-th edges for intersecting. 
	--  Remark : See the previous method for details
	
    CheckIntersectingEdges(me: mutable; num1: Integer; num2: Integer)
    returns Boolean;
    	---Purpose: Checks i-th and j-th edges for intersecting.
	--  Remark : Calls  previous method.
    	--  Status : See the function above for details

    CheckLacking (me: mutable; num: Integer; Tolerance: Real;
                              p2d1, p2d2: out Pnt2d from gp) returns Boolean;
    	---Purpose: Checks if there is a gap in 2d between edges, not comprised by 
        --          the tolerance of their common vertex.
	--          If <Tolerance> is greater than 0. and less than tolerance of
        --          the vertex, then this value is used for check.
    	--  Returns: True if not closed gap was detected
	--          p2d1 and p2d2 are the endpoint of <num-1>th edge and start of
	--          the <num>th edge in 2d.
    	--  Status:
    	--	    OK: No edge is lacking (3d and 2d connection)
	--          FAIL1: edges have no vertices (at least one of them)
	--          FAIL2: edges are neither connected by common vertex, nor have 
        --                 coincided vertices
	--          FAIL1: edges have no pcurves
    	--          DONE1: the gap is detected which cannot be closed by the tolerance
        --                 of the common vertex (or with value of <Tolerance>)
    	--          DONE2: is set (together with DONE1) if gap is detected and the 
        --                 vector (p2d2 - p2d1) goes in direction opposite to the pcurves
        --                 of the edges (if angle is more than 0.9*PI).

    CheckLacking (me : mutable; num: Integer; Tolerance: Real = 0.0) returns Boolean;
    	---Purpose: Checks if there is a gap in 2D between edges and not comprised by vertex tolerance
   	 --         The value of SBWD.thepreci is used.
    	--  Returns: False if no edge should be inserted
    	--  Status:
    	--	     OK    : No edge is lacking (3d and 2d connection)
    	--          DONE1 : The vertex tolerance should be increased only (2d gap is 
    	--                  small)
    	--          DONE2 : Edge can be inserted (3d and 2d gaps are large enough)

    CheckOuterBound (me: mutable; APIMake: Boolean = Standard_True)
    returns Boolean;
    	---Purpose: Checks if wire defines an outer bound on the face
	--          Uses ShapeAnalysis::IsOuterBound for analysis
	--          If <APIMake> is True uses BRepAPI_MakeWire to build the
    	--          wire, if False (to be used only when edges share common
	--          vertices) uses BRep_Builder to build the wire
	--          
    	---Returns: False if wire is an outer bound, else returns True
    	--  Status:
    	--	    OK   : If it is an outer wire
    	--          DONE : If not

    CheckNotchedEdges(me : mutable; num      : Integer; 
    	    	    	    	    shortNum : out Integer;
    	    	    	    	    param    : out Real;
    	    	    	    	    Tolerance: Real = 0.0) returns Boolean;
    	---Purpose: Detects a notch

    CheckSmallArea (me: mutable; theWire : Wire from TopoDS; theIsOuterWire : Boolean)
    returns Boolean;
    	---Purpose: Checks if wire has parametric area less than precision.
		 
    CheckShapeConnect (me : mutable; shape : Shape from TopoDS; prec: Real = 0.0)
    returns Boolean;
    	---Purpose: Checks with what orientation <shape> (wire or edge) can be 
    	--           connected to the wire.
    	--           Tests distances with starting <preci> from <SBWD> (close confusion), 
    	--	     but if given <prec> is greater, tests with <prec> (coarse confusion).
    	--           The smallest found distance can be returned by MinDistance3d
    	--           
    	--  Returns: False if status is FAIL (see below)
    	--  Status:
    	--	     DONE1 : If <shape> follows <SBWD>, direct sense (normal)
    	--           DONE2 : If <shape> follows <SBWD>, but if reversed
    	--           DONE3 : If <shape> preceeds <SBWD>, direct sense
    	--           DONE4 : If <shape> preceeds <SBWD>, but if reversed
    	--           FAIL1 : If <shape> is neither an edge nor a wire 
    	--           FAIL2 : If <shape> cannot be connected to <SBWD>
	--
	--           DONE5 : To the tail of <SBWD> the <shape> is closer with
    	--                   direct sense
	--           DONE6 : To the head of <SBWD> the <shape> is closer with
    	--                   direct sense
	--
	--  Remark:   Statuses DONE1 - DONE4, FAIL1 - FAIL2 are basic and
        --           describe the nearest connection of the <shape> to <SBWD>.
	--           Statuses DONE5 and DONE6 are advanced and are to be used when
	--           analyzing with what sense (direct or reversed) the <shape>
	--           should be connected to <SBWD>:
    	--           For tail of <SBWD> if DONE4 is True <shape> should be direct,
        --           otherwise reversed.
    	--           For head of <SBWD> if DONE5 is True <shape> should be direct,
        --           otherwise reversed.
	
    CheckShapeConnect (me : mutable; tailhead: out Real;
    	    	                    tailtail: out Real;
    	    	                    headtail: out Real;
    	    	                    headhead: out Real;
    	    	                    shape   : Shape from TopoDS;
                                    prec    : Real = 0.0)
    returns Boolean;
    	---Purpose: The same as previous CheckShapeConnect but is more advanced.
	--          It returns the distances between each end of <sbwd> and each
	--          end of <shape>. For example, <tailhead> stores distance
    	--          between tail of <sbwd> and head of <shape>
	--  Remark:  First method CheckShapeConnect calls this one

    CheckLoop (me : mutable; aMapLoopVertices : out IndexedMapOfShape from TopTools;
    	    	    	     aMapVertexEdges :out DataMapOfShapeListOfShape from TopTools;
    	    	    	     aMapSmallEdges : out MapOfShape from TopTools;
    	    	    	     aMapSeemEdges : out MapOfShape from TopTools) returns Boolean;
    	---Purpose: Checks existance of loop on wire and return vertices wich are loop vertices 
-- (vertices belonging to a few pairs of edges)
	
    	
    	---Status after checking :
    
    	---Level  : Public

    	-- Querying the status of perfomed API checking procedures
    StatusOrder            (me; Status: Status from ShapeExtend) returns Boolean;
    	---C++: inline
    StatusConnected        (me; Status: Status from ShapeExtend) returns Boolean;
    	---C++: inline
    StatusEdgeCurves       (me; Status: Status from ShapeExtend) returns Boolean;
    	---C++: inline
    StatusDegenerated      (me; Status: Status from ShapeExtend) returns Boolean;
    	---C++: inline
    StatusClosed           (me; Status: Status from ShapeExtend) returns Boolean;
    	---C++: inline
    StatusSmall            (me; Status: Status from ShapeExtend) returns Boolean;
    	---C++: inline
    StatusSelfIntersection (me; Status: Status from ShapeExtend) returns Boolean;
    	---C++: inline
    StatusLacking          (me; Status: Status from ShapeExtend) returns Boolean;
    	---C++: inline
    StatusGaps3d           (me; Status: Status from ShapeExtend) returns Boolean;
    	---C++: inline
    StatusGaps2d           (me; Status: Status from ShapeExtend) returns Boolean;
    	---C++: inline
    StatusCurveGaps        (me; Status: Status from ShapeExtend) returns Boolean;
    	---C++: inline

    StatusLoop             (me; Status: Status from ShapeExtend) returns Boolean;
    	---C++: inline
    	---Level  : Advanced

    LastCheckStatus        (me; Status: Status from ShapeExtend) returns Boolean;
    	---C++: inline
    	---Purpose:  Querying the status of the LAST perfomed 'Advanced' checking procedure

    	---Querying fields
    
    MinDistance3d (me) returns Real;
    	---C++: inline
    	---Purpose: Returns the last lowest distance in 3D computed by
    	--           CheckOrientation, CheckConnected, CheckContinuity3d, 
    	--	         CheckVertex, CheckNewVertex

    MinDistance2d (me) returns Real;
    	---C++: inline
    	---Purpose: Returns the last lowest distance in 2D-UV computed by
    	--           CheckContinuity2d

    MaxDistance3d (me) returns Real;
    	---C++: inline
    	---Purpose: Returns the last maximal distance in 3D computed by
    	--           CheckOrientation, CheckConnected, CheckContinuity3d, 
    	--	         CheckVertex, CheckNewVertex, CheckSameParameter

    MaxDistance2d (me) returns Real;
    	---C++: inline
    	---Purpose: Returns the last maximal distance in 2D-UV computed by
    	--           CheckContinuity2d
    
fields

    myWire: WireData from ShapeExtend is protected;
    myFace: Face from TopoDS is protected;
    mySurf: Surface from ShapeAnalysis is protected;
    myPrecision : Real is protected;

    myMin3d: Real is protected; -- lower computed distance 3d
    myMin2d: Real is protected; -- lower computed distance 2d
    myMax3d: Real is protected; -- upper computed distance 3d
    myMax2d: Real is protected; -- upper computed distance 2d
    
    	-- statuses corresponding to API methods, queried by Status..(status) methods
    myStatusOrder:            Integer is protected;
    myStatusConnected:        Integer is protected;
    myStatusEdgeCurves:       Integer is protected;
    myStatusDegenerated:      Integer is protected;
    myStatusClosed:           Integer is protected;
    myStatusSmall:            Integer is protected;
    myStatusSelfIntersection: Integer is protected;
    myStatusLacking:          Integer is protected;
    myStatusGaps3d:           Integer is protected; -- szvsh
    myStatusGaps2d:           Integer is protected; -- szvsh
    myStatusCurveGaps:        Integer is protected; -- szvsh
    myStatusLoop  :           Integer is protected;
    
    myStatus: Integer is protected; -- for internal use, queried by LastCheckStatus(status) method

end Wire;
