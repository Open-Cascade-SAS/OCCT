-- Created on: 1991-05-13
-- Created by: Laurent PAINNOT
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.





deferred class MultipleVarFunctionWithGradient from math

inherits MultipleVarFunction
---Purpose:
-- The abstract class MultipleVarFunctionWithGradient
-- describes the virtual functions associated with a multiple variable function.
uses Vector from math

is

    Delete(me:out) is virtual;
    ---C++: alias "Standard_EXPORT virtual ~math_MultipleVarFunctionWithGradient(){Delete();}"
    
    NbVariables(me)
    	---Purpose: Returns the number of variables of the function.

    returns Integer
    is deferred;


    Value(me: in out; X: Vector; F: out Real)
    	---Purpose: Computes the values of the Functions <F> for the   variable <X>.
    	--          Returns True if the computation was done successfully, 
    	--          False otherwise.

    returns Boolean
    is deferred;
    
    
    Gradient(me: in out; X: Vector; G: out Vector)
    	---Purpose: Computes the gradient <G> of the functions for the   variable <X>.
    	--         Returns True if the computation was done successfully, 
    	--         False otherwise.

    returns Boolean
    is deferred;
    
    
    Values(me: in out; X: Vector; F: out Real; G: out Vector)
    	---Purpose: computes the value <F> and the gradient <G> of the 
    	--          functions for the variable <X>.
    	--          Returns True if the computation was done successfully, 
    	--          False otherwise.

    returns Boolean
    is deferred;
    
end MultipleVarFunctionWithGradient;
