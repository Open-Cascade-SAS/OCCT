-- File:        SurfaceStyleFillArea.cdl
-- Created:     Mon Dec  4 12:02:31 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWSurfaceStyleFillArea from RWStepVisual

	---Purpose : Read & Write Module for SurfaceStyleFillArea

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     SurfaceStyleFillArea from StepVisual,
     EntityIterator from Interface

is

	Create returns RWSurfaceStyleFillArea;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable SurfaceStyleFillArea from StepVisual);

	WriteStep (me; SW : in out StepWriter; ent : SurfaceStyleFillArea from StepVisual);

	Share(me; ent : SurfaceStyleFillArea from StepVisual; iter : in out EntityIterator);

end RWSurfaceStyleFillArea;
