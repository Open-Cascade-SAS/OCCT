-- Created on: 1993-07-08
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class HBoxTool from TopOpeBRepTool inherits TShared from MMgt

uses

    Box from Bnd,
    Shape from TopoDS,
    ShapeEnum from TopAbs,
    IndexedDataMapOfShapeBox from TopOpeBRepTool
    
is
    
    Create returns mutable HBoxTool from TopOpeBRepTool;
    Clear(me:mutable);
    AddBoxes(me:mutable;S:Shape;TS:ShapeEnum;TA:ShapeEnum=TopAbs_SHAPE);
    AddBox(me:mutable;S:Shape);

    ComputeBox(myclass;S:Shape;B:out Box from Bnd);
    ComputeBoxOnVertices(myclass;S:Shape;B:out Box from Bnd);
    DumpB(myclass;B:Box from Bnd);

    Box(me:mutable;S:Shape) returns Box from Bnd;---C++: return const &
    Box(me; I:Integer) returns Box from Bnd;---C++: return const &
    HasBox(me; S:Shape) returns Boolean;
    Shape(me; I:Integer) returns Shape;---C++: return const &
    Index(me; S:Shape) returns Integer;
    Extent(me) returns Integer;
    ChangeIMS(me:mutable) returns IndexedDataMapOfShapeBox;---C++:return &
    IMS(me) returns IndexedDataMapOfShapeBox;---C++:return const &
    
fields

    myIMS:IndexedDataMapOfShapeBox from TopOpeBRepTool;

end HBoxTool;
