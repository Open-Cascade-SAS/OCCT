-- Created on: 1994-05-31
-- Created by: Christian CAILLET
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SelectName  from IGESSelect  inherits  SelectExtract

    ---Purpose : Selects Entities which have a given name.
    --           Consider Property Name if present, else Short Label, but
    --           not the Subscript Number
    --           First version : keeps exact name
    --           Later : regular expression

uses AsciiString from TCollection, HAsciiString from TCollection,
     Transient, InterfaceModel

is

    Create returns mutable SelectName;
    ---Purpose : Creates an empty SelectName : every entity is considered
    --           good (no filter active)

    Sort (me; rank : Integer; ent : Transient; model : InterfaceModel)
    	returns Boolean;
    ---Purpose : Returns True if Name of Entity complies with Name Filter

    SetName (me : mutable; name : HAsciiString from TCollection);
    ---Purpose : Sets a Name as a criterium : IGES Entities which have this name
    --           are kept (without regular expression, there should be at most
    --           one). <name> can be regarded as a Text Parameter

    Name (me) returns HAsciiString from TCollection;
    ---Purpose : Returns the Name used as Filter

    ExtractLabel (me) returns AsciiString from TCollection;
    ---Purpose : Returns the Selection criterium : "IGES Entity, Name : <name>"

fields

    thename : HAsciiString from TCollection;

end SelectName;
