-- Created on: 1997-08-13
-- Created by: Jean-Louis Frenkel
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class DirectoryIterator from CDF

uses
    Directory from CDF,
    Document from CDM,
    ListIteratorOfListOfDocument from CDM
raises
    NoSuchObject from Standard

is

    Create
    returns DirectoryIterator from CDF;
    ---Purpose: creates an Iterator with the directory 
    --          of the current CDF.

    Create(aDirectory: Directory from CDF) 
    returns  DirectoryIterator from CDF;

    MoreDocument (me: in out) returns Boolean from Standard;
    ---Purpose : Returns True if there are more entries to return
    
    NextDocument (me: in out);
    ---Purpose : Go to the next entry
    --           (if there is not, Value will raise an exception)
    
    Document (me: in out) returns Document from CDM
    ---Purpose : Returns item value of current entry
    raises NoSuchObject  from Standard;

fields

    myIterator: ListIteratorOfListOfDocument from CDM;
end DirectoryIterator from CDF;
