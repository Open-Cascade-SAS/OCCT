-- Created on: 1995-12-04
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package RWStepRepr 

uses

	StepData, Interface, TCollection, TColStd, StepRepr

is


--class ReadWriteModule;

--class GeneralModule;

class RWDefinitionalRepresentation;
class RWDescriptiveRepresentationItem;
class RWFunctionallyDefinedTransformation;
class RWGlobalUncertaintyAssignedContext;
class RWGlobalUnitAssignedContext;
class RWItemDefinedTransformation;
--moved to StepBasic: class RWGroup;
--moved to StepBasic: class RWGroupRelationship;
class RWMappedItem;
class RWParametricRepresentationContext;
class RWProductDefinitionShape;
class RWPropertyDefinition;
class RWPropertyDefinitionRepresentation;
--moved to StepAP214: class RWRepItemGroup;
class RWRepresentation;
class RWRepresentationContext;
class RWRepresentationItem;
class RWRepresentationMap;
class RWRepresentationRelationship;

class RWShapeAspect;
class RWShapeAspectRelationship;
class RWShapeAspectTransition;
-- class RWShapeDefinitionRepresentation;  moved to StepShape

    	-- Added from AP214 CC1 to CC2

class RWMakeFromUsageOption;
class RWAssemblyComponentUsage;
class RWQuantifiedAssemblyComponentUsage;
class RWSpecifiedHigherUsageOccurrence;

class RWAssemblyComponentUsageSubstitute;

class RWRepresentationRelationshipWithTransformation;
class RWShapeRepresentationRelationshipWithTransformation;

class RWMaterialDesignation;

-- ABV added for CAX TRJ 2 validation properties
class RWMeasureRepresentationItem;

    -- Added for AP203
    class RWConfigurationDesign;
    class RWConfigurationEffectivity;
    class RWConfigurationItem;
    class RWProductConcept;

    -- Added for Dimensional Tolerancing (CKY 25 APR 2001 for TR7J)
    class RWCompoundRepresentationItem;

	---Package Method ---

--- added for AP209
    class RWDataEnvironment;
    class RWMaterialPropertyRepresentation;
    class RWPropertyDefinitionRelationship;
    class RWMaterialProperty;
    class RWStructuralResponseProperty;
    class RWStructuralResponsePropertyDefinitionRepresentation;

--- added for TR12J (GD&T) 
    class RWCompositeShapeAspect;
    class RWDerivedShapeAspect;
    class RWExtension;
    class RWShapeAspectDerivingRelationship;
    class RWReprItemAndLengthMeasureWithUnit;
    
--	Init;
	---Purpose: enforced the initialisation of the  libraries

end RWStepRepr;
