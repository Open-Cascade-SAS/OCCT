-- Created on: 1997-06-25
-- Created by: Philippe MANGIN
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred  class SweepFunction from Approx inherits TShared from MMgt  

	---Purpose: defined the function used by SweepApproximation to
	--          perform sweeping application.
          

uses 
 Shape            from GeomAbs,
 Pnt              from gp, 
 Array1OfPnt      from TColgp,
 Array1OfPnt2d    from TColgp,
 Array1OfVec      from TColgp,
 Array1OfVec2d    from TColgp, 
 Array1OfInteger  from TColStd,
 Array1OfReal     from TColStd

raises NotImplemented , 
       OutOfRange from  Standard

is   

-- 
--========== To compute Sections and derivatives Sections
--   
   D0(me : mutable; 
      Param: Real;
      First, Last : Real; 
      Poles    : out Array1OfPnt   from TColgp;
      Poles2d  : out Array1OfPnt2d from TColgp;
      Weigths  : out Array1OfReal  from TColStd)
      ---Purpose: compute the section for v = param           
   returns Boolean  is  deferred;
	
   D1(me : mutable;
      Param: Real;
      First, Last : Real; 
      Poles    : out Array1OfPnt   from TColgp;
      DPoles   : out Array1OfVec   from TColgp;
      Poles2d  : out Array1OfPnt2d from TColgp;
      DPoles2d : out Array1OfVec2d from TColgp;
      Weigths  : out Array1OfReal  from TColStd;
      DWeigths : out Array1OfReal  from TColStd)
      ---Purpose: compute the first  derivative in v direction  of the
      --           section for v =  param 
      --  Warning : It used only for C1 or C2 aproximation
   returns Boolean  
   raises  NotImplemented 
   is  virtual; 
   
    D2(me : mutable;
      Param: Real;
      First, Last : Real; 
      Poles     : out Array1OfPnt   from TColgp;
      DPoles    : out Array1OfVec   from TColgp;
      D2Poles   : out Array1OfVec   from TColgp;
      Poles2d   : out Array1OfPnt2d from TColgp;
      DPoles2d  : out Array1OfVec2d from TColgp;
      D2Poles2d : out Array1OfVec2d from TColgp;
      Weigths   : out Array1OfReal  from TColStd;
      DWeigths  : out Array1OfReal  from TColStd;
      D2Weigths : out Array1OfReal  from TColStd)      
      ---Purpose: compute the second derivative  in v direction of the
      --          section  for v = param  
      --  Warning : It used only for C2 aproximation
   returns Boolean 
   raises  NotImplemented  
   is  virtual; 
    
-- 
--   =================== General Information On The Function  ===================
--                                         
   Nb2dCurves(me)     
     ---Purpose: get the number of 2d curves to  approximate.
   returns Integer  is  deferred;  

   SectionShape(me; NbPoles   : out Integer from Standard;
                    NbKnots   : out Integer from Standard;
                    Degree    : out Integer from Standard) 
	---Purpose: get the format of an  section
    is  deferred;  
    
    Knots(me; TKnots: out Array1OfReal from TColStd)
	---Purpose: get the Knots of the section 
	is deferred;

    Mults(me; TMults: out Array1OfInteger from TColStd)
	---Purpose: get the Multplicities of the section          
	is deferred;   

    IsRational(me)
	---Purpose: Returns if the sections are rationnal or not         
    returns Boolean  is deferred; 

          
--
--  =================== Management  of  continuity  ===================
--                 
    NbIntervals(me; S : Shape from GeomAbs) 
	---Purpose: Returns  the number  of  intervals for  continuity
	--          <S>. 
        --          May be one if Continuity(me) >= <S>
   returns Integer  is  deferred;

   Intervals(me; T : in out Array1OfReal from TColStd; 
    	         S : Shape from GeomAbs)
	---Purpose: Stores in <T> the  parameters bounding the intervals
	--          of continuity <S>.
	--          
	--          The array must provide  enough room to  accomodate
	--          for the parameters. i.e. T.Length() > NbIntervals()
    raises
    	OutOfRange from Standard 
    is deferred;  
     
    	
   SetInterval(me: mutable; First, Last: Real from Standard)    
	---Purpose: Sets the bounds of the parametric interval on 
	--          the fonction
	--          This determines the derivatives in these values if the
	--          function is not Cn.
    	is deferred; 
   

--  ===================== To  help  computation  of  Tolerance ======
--      Evaluation of error, in 2d space, or on rational function, is
--      difficult.  The following methods can help the approximation to
--      make good evaluation and use good tolerances.
--      
--       It is not necessary for the following informations to be very
--       precise. A fast evaluation is sufficient.
     
   Resolution(me;   
              Index       :  Integer  from  Standard;
   	      Tol         : Real from Standard;   
              TolU,  TolV :  out Real  from Standard)  
   ---Purpose: Returns the resolutions in the  sub-space 2d <Index>
   --          This information is usfull to find an good tolerance in
   --          2d approximation.              
  ---Warning: Used only if Nb2dCurve > 0          
  raises  NotImplemented   
  is virtual;
    
 
   GetTolerance(me;  
    	    	BoundTol, SurfTol, AngleTol : Real;
		Tol3d : out Array1OfReal)
	---Purpose: Returns the tolerance to reach in approximation
	--          to satisfy.
	--          BoundTol error at the Boundary
	--          AngleTol tangent error at the Boundary (in radian)
	--          SurfTol error inside the surface.         
  is  deferred; 
   
  
  SetTolerance(me :  mutable; Tol3d,  Tol2d  :  Real) 
        ---Purpose: Is usefull, if (me) have to run numerical
        --           algorithm to perform D0, D1 or D2        
  is  deferred; 
   
  BarycentreOfSurf(me) 
   ---Purpose:  Get the barycentre of Surface.   
   --          An   very  poor estimation is sufficent. 
   --          This information is usefull to perform well 
   --          conditioned rational approximation. 
   --  Warning: Used only if <me> IsRational         
   returns Pnt from gp    
   raises  NotImplemented   
   is  virtual; 
      
	
   MaximalSection(me) returns Real
    	---Purpose: Returns the   length of the greater section. This
    	--          information is usefull to G1's control.
        --  Warning: With an little value, approximation can be slower.          
   raises  NotImplemented   
   is virtual;
    
   GetMinimalWeight(me; Weigths  : out Array1OfReal  from TColStd)
    	---Purpose: Compute the minimal value of weight for each poles
    	--          in all  sections.  
        --          This information is  usefull to control error
    	--          in rational approximation.
        --  Warning: Used only if <me> IsRational        
   raises  NotImplemented   
   is virtual;
   
end SweepFunction;
