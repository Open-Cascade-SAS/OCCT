-- Created on: 1998-06-30
-- Created by: Christian CAILLET
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class RepresentationRelationshipWithTransformation  from StepRepr
    inherits ShapeRepresentationRelationship

    -- in principle, inherits RepresentationRelationship
    -- But <Shape>... only adds a constraint on a field, this allows to
    -- simplify the multiple inheritance between ShapeRR and RRWithTransf...

uses
     HAsciiString from TCollection,
     Representation from StepRepr,
     Transformation from StepRepr

is

    Create returns mutable RepresentationRelationshipWithTransformation;

    Init (me : mutable;
              aName : mutable HAsciiString from TCollection;
              aDescription : mutable HAsciiString from TCollection;
              aRep1 : mutable Representation from StepRepr;
              aRep2 : mutable Representation from StepRepr;
	      aTransf : Transformation);

    TransformationOperator (me) returns Transformation;
    SetTransformationOperator (me : mutable; aTrans : Transformation);

fields

    theTrans : Transformation;

end RepresentationRelationshipWithTransformation;
