-- Created on: 1993-12-02
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

generic class PointOnRst from Blend
    (TheArc    as any)


	---Purpose: Definition of an intersection point between a line
	--          and a restriction on a surface.
	--          Such a point is contains geometrical informations (see
	--          the Value method) and logical informations.


uses Transition from IntSurf
     
raises DomainError from Standard

is


    Create
    
	---Purpose: Empty constructor.

    	returns PointOnRst from Blend;


    Create( A: TheArc; Param: Real from Standard;
            TLine, TArc: Transition from IntSurf)

	---Purpose: Creates the PointOnRst on the arc A, at parameter Param,
	--          with the transition TLine on the walking line, and
	--          TArc on the arc A.

    	returns PointOnRst from Blend;



    SetArc(me: in out; A: TheArc; Param: Real from Standard;
                       TLine, TArc: Transition from IntSurf)

	---Purpose: Sets the values of a point which is on the arc
	--          A, at parameter Param.


    	is static;



    Arc(me)
    
	---Purpose: Returns the arc of restriction containing the
	--          vertex.

    	returns any TheArc
	---C++: return const&
	---C++: inline
	
	is static;


    TransitionOnLine(me)
    
	---Purpose: Returns the transition of the point on the
	--          line on surface.

    	returns Transition from IntSurf
	---C++: return const&
	---C++: inline
	
	is static;


    TransitionOnArc(me)
    
	---Purpose: Returns the transition of the point on the arc
	--          returned by Arc().

    	returns Transition from IntSurf
	---C++: return const&
	---C++: inline
	
	is static;


    ParameterOnArc(me)
    
	---Purpose: Returns the parameter of the point on the
	--          arc returned by the method Arc().

    	returns Real from Standard
	---C++: inline
	
	is static;


fields

    arc       : TheArc;
    traline   : Transition from IntSurf;
    traarc    : Transition from IntSurf;
    prm       : Real       from Standard;

end PointOnRst;
