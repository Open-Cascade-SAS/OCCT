-- Created on: 1999-09-17
-- Created by: Denis PASCAL
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PathParser from TDocStd 

	---Purpose: parse an OS path

uses ExtendedString from TCollection

is 
    Create (path : ExtendedString from TCollection) returns PathParser from TDocStd;
    Parse (me : in out);
    Trek(me) returns ExtendedString from TCollection;
    Name(me) returns ExtendedString from TCollection;
    Extension(me) returns ExtendedString from TCollection;
    Path(me) returns ExtendedString from TCollection;  
    Length (me) returns Integer from Standard;
    
fields 
    myPath      : ExtendedString from TCollection;
    myExtension : ExtendedString from TCollection;
    myTrek      : ExtendedString from TCollection;
    myName      : ExtendedString from TCollection;
end;
