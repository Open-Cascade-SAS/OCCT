-- Created on: 1994-10-03
-- Created by: Yves FRICAUD
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package BRepMAT2d 

	---Purpose: 

uses
    MAT2d,
    MAT,
    TCollection,
    TColStd,
    TColGeom2d,
    Geom2d,
    gp,	
    TopoDS,
    TopTools
    
is
    class Explorer;
    	---Purpose: Construct an  explorer for  the computation of the 
    	--          bisecting locus  from a Wire, a  Face, or a set of 
    	--          curves from Geom2d.

    class BisectingLocus instantiates BisectingLocus from MAT2d 
    	    	    	    	    	  (Explorer  from BRepMAT2d);
	---Purpose: the map of bisecting locus.
					  
    class LinkTopoBilo;
    	---Purpose: Constucts links between the Wire or the Face and
    	--          the BasicElts contained in the bisecting locus.


    class SequenceOfBasicElt instantiates Sequence from TCollection
                                                         (BasicElt from MAT); 
							 
    class DataMapOfShapeSequenceOfBasicElt instantiates DataMap from TCollection 
    		    		    	      (Shape               from TopoDS, 
					       SequenceOfBasicElt  from  BRepMAT2d, 
					       ShapeMapHasher      from TopTools); 
    
    class DataMapOfBasicEltShape  instantiates
    	DataMap from TCollection (BasicElt            from MAT,
    	    	    	    	  Shape               from TopoDS,
    	    	    	    	  MapTransientHasher  from TColStd);				       

end BRepMAT2d;




