-- Created on: 1993-01-27
-- Created by: Jean-Louis Frenkel
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.





class ShapeTool from Prs3d


uses
    Shape             from TopoDS,
    Face              from TopoDS,
    Edge              from TopoDS,
    Vertex            from TopoDS,
    HSequenceOfShape  from TopTools,
    Box               from Bnd,
    Location          from TopLoc,
    Triangulation     from Poly,
    PolygonOnTriangulation     from Poly,
    Polygon3D         from Poly,
    HArray1OfInteger  from TColStd,
    Explorer          from TopExp,
    IndexedDataMapOfShapeListOfShape from TopTools,
    IndexedMapOfShape                from TopTools

	---Purpose: 
is

    Create ( TheShape: Shape from TopoDS) returns ShapeTool from Prs3d;
    InitFace (me: in out);
    MoreFace (me) returns Boolean from Standard;
    NextFace (me: in out);
    GetFace(me) returns Face from TopoDS;
    	---C++: return const&
    FaceBound(me) returns Box from Bnd;
    IsPlanarFace(me) returns Boolean from Standard;

    InitCurve (me: in out);
    MoreCurve (me) returns Boolean from Standard;
    NextCurve (me: in out);
    GetCurve(me) returns Edge from TopoDS;
    	---C++: return const&
    CurveBound(me) returns Box from Bnd;
    Neighbours(me) returns Integer from Standard;   
    FacesOfEdge(me) returns HSequenceOfShape from TopTools;

    InitVertex(me: in out);
    MoreVertex(me) returns Boolean from Standard;
    NextVertex(me: in out);
    GetVertex(me) returns Vertex from TopoDS;
    	---C++: return const&

    HasSurface(me) returns Boolean;
    
    CurrentTriangulation(me; l: out Location from TopLoc) 
    returns Triangulation from Poly;

    HasCurve(me) returns Boolean;

    PolygonOnTriangulation(me; Indices: out PolygonOnTriangulation from  Poly;
    	    	    	       T:       out Triangulation          from Poly; 
			       l:       out Location               from TopLoc); 
			       
    Polygon3D(me; l: out Location from TopLoc) 
    returns Polygon3D from Poly;

fields
    myShape:        Shape                            from TopoDS;
    myFaceExplorer: Explorer                         from TopExp;
    myEdgeMap:      IndexedDataMapOfShapeListOfShape from TopTools;
    myVertexMap:    IndexedMapOfShape                from TopTools;
    myEdge :        Integer                          from Standard;
    myVertex :      Integer                          from Standard;

end ShapeTool from Prs3d;
