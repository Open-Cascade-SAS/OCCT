-- Created on: 1999-11-26
-- Created by: Andrey BETENEV
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0

class CcDesignDateAndTimeAssignment from StepAP203
inherits DateAndTimeAssignment from StepBasic

    ---Purpose: Representation of STEP entity CcDesignDateAndTimeAssignment

uses
    DateAndTime from StepBasic,
    DateTimeRole from StepBasic,
    HArray1OfDateTimeItem from StepAP203

is
    Create returns CcDesignDateAndTimeAssignment from StepAP203;
	---Purpose: Empty constructor

    Init (me: mutable; aDateAndTimeAssignment_AssignedDateAndTime: DateAndTime from StepBasic;
                       aDateAndTimeAssignment_Role: DateTimeRole from StepBasic;
                       aItems: HArray1OfDateTimeItem from StepAP203);
	---Purpose: Initialize all fields (own and inherited)

    Items (me) returns HArray1OfDateTimeItem from StepAP203;
	---Purpose: Returns field Items
    SetItems (me: mutable; Items: HArray1OfDateTimeItem from StepAP203);
	---Purpose: Set field Items

fields
    theItems: HArray1OfDateTimeItem from StepAP203;

end CcDesignDateAndTimeAssignment;
