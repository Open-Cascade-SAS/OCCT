-- Created on: 2003-06-04
-- Created by: Galina KULIKOVA
-- Copyright (c) 2003-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class DatumReference from StepDimTol
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity DatumReference

uses
    Datum from StepDimTol

is
    Create returns DatumReference from StepDimTol;
	---Purpose: Empty constructor

    Init (me: mutable; aPrecedence: Integer;
                       aReferencedDatum: Datum from StepDimTol);
	---Purpose: Initialize all fields (own and inherited)

    Precedence (me) returns Integer;
	---Purpose: Returns field Precedence
    SetPrecedence (me: mutable; Precedence: Integer);
	---Purpose: Set field Precedence

    ReferencedDatum (me) returns Datum from StepDimTol;
	---Purpose: Returns field ReferencedDatum
    SetReferencedDatum (me: mutable; ReferencedDatum: Datum from StepDimTol);
	---Purpose: Set field ReferencedDatum

fields
    thePrecedence: Integer;
    theReferencedDatum: Datum from StepDimTol;

end DatumReference;
