-- File:	RWStepElement_RWSurface3dElementDescriptor.cdl
-- Created:	Thu Dec 12 17:29:04 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWSurface3dElementDescriptor from RWStepElement

    ---Purpose: Read & Write tool for Surface3dElementDescriptor

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    Surface3dElementDescriptor from StepElement

is
    Create returns RWSurface3dElementDescriptor from RWStepElement;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : Surface3dElementDescriptor from StepElement);
	---Purpose: Reads Surface3dElementDescriptor

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: Surface3dElementDescriptor from StepElement);
	---Purpose: Writes Surface3dElementDescriptor

    Share (me; ent : Surface3dElementDescriptor from StepElement;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWSurface3dElementDescriptor;
