-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


---Version:	 1.2 

--  Version	Date		Purpose
--         	Feb  3 1995	Creation
--         	Dec  15 1996    Version CSFDB

package ObjMgt 

---Purpose: This package defines services to manage the storage grain of data 
--          produced by applications and those classes to manage persistent 
--          extern reference.

uses

    PCollection,
    Storage,
    CDM,PCDM, TCollection

is

    --deferred class RetrievalDriver;
    ---Purpose: to retrieve ExternShareable objects in the framework.
 

    deferred class ExternShareable;
    ---Purpose: Defines the root persistent object which can be persistent 
    --          extern reference.

    private class ExternRef;
    ---Purpose: Defines (objet-relais) to implement extern reference.

    private class PSeqOfExtRef instantiates HSequence from 
    	    PCollection (ExternRef from ObjMgt);

end ObjMgt;
