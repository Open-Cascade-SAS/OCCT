-- Created on: 1999-06-17
-- Created by: data exchange team
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package ShapeProcessAPI

    ---Purpose: Provides tools for converting shapes for data exchange
    --          between various systems (CATIA, EUCLID3 etc.)

uses

    TopAbs,
    TopoDS,
    TopTools,
    Message,
    ShapeProcess,
    TCollection
    
is

    class ApplySequence;
    	---Purpose: Applies one of the sequence of calls from resource file.
    
end ShapeProcessAPI;
