-- Created on: 1995-03-09
-- Created by: Laurent PAINNOT
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Polygon3D from BRep inherits CurveRepresentation from BRep

	---Purpose: 

uses
    Polygon3D           from Poly,
    CurveRepresentation from BRep,
    Location            from TopLoc

raises DomainError from Standard

is

    Create(P: Polygon3D from Poly;
    	   L: Location  from TopLoc) 
    	---Purpose:

    returns mutable Polygon3D from BRep;
    
    
    IsPolygon3D(me) returns Boolean
    	---Purpose: Returns True.
    is redefined;
    
    Polygon3D(me) returns any Polygon3D from Poly
    	---C++: return const&
    is redefined;
    
    Polygon3D(me: mutable; P: Polygon3D from Poly)
    raises
    	DomainError from Standard
    is redefined;

    Copy(me) returns mutable CurveRepresentation from BRep;
	---Purpose: Return a copy of this representation.


fields

myPolygon3D: Polygon3D from Poly;


end Polygon3D;
