-- Created on: 1997-02-21
-- Created by: Laurent BOURESCHE
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


deferred class SurfCurvFuncInv from Blend

inherits FunctionSetWithDerivatives from math


    ---Purpose: Deferred   class  for a  function  used  to compute  a
    --          blending surface between a  surface and a curve, using
    --          a  guide  line.   This   function is  used  to find  a
    --          solution on a done restriction of the surface.
    --          
    --          The vector  <X> used in  Value, Values and Derivatives
    --          methods  has   to  be the   vector  of  the parametric
    --          coordinates  wguide, wcurv, wrst  where  wguide is the
    --          parameter on the guide line, wcurv is the parameter on
    --          the curve, wrst is the parameter on the restriction on
    --          the surface.

uses
    HCurve2d from Adaptor2d,
    Vector   from math,
    Matrix   from math


is

    NbVariables(me)
    ---Purpose: Returns 3.
    returns Integer from Standard
    is static;

    NbEquations(me)
    ---Purpose: returns the number of equations of the function.
    returns Integer from Standard
    is deferred;

    Value(me: in out; X: Vector; F: out Vector)
    ---Purpose: computes the values <F> of the Functions for the 
    --          variable <X>.
    --          Returns True if the computation was done successfully, 
    --          False otherwise.
    returns Boolean from Standard
    is deferred;
    
    Derivatives(me: in out; X: Vector; D: out Matrix)
    ---Purpose: returns the values <D> of the derivatives for the 
    --          variable <X>.
    --          Returns True if the computation was done successfully, 
    --          False otherwise.
    returns Boolean from Standard
    is deferred;
    
    Values(me: in out; X: Vector; F: out Vector; D: out Matrix)
    ---Purpose: returns the values <F> of the functions and the derivatives
    --          <D> for the variable <X>.
    --          Returns True if the computation was done successfully, 
    --          False otherwise.
    returns Boolean from Standard
    is deferred;

    Set(me: in out; Rst : HCurve2d from Adaptor2d)
    ---Purpose: Set the Point on which a solution has to be found. 
    is deferred;

    GetTolerance(me; Tolerance: out Vector from math; Tol: Real from Standard)
    ---Purpose: Returns in the vector Tolerance the parametric tolerance
    --          for each of the 3 variables;
    --          Tol is the tolerance used in 3d space.
    is deferred;

    GetBounds(me; InfBound,SupBound: out Vector from math)
    ---Purpose: Returns in the vector InfBound the lowest values allowed
    --          for each of the 3 variables.
    --          Returns in the vector SupBound the greatest values allowed
    --          for each of the 3 variables.
    is deferred;


    IsSolution(me: in out; Sol: Vector from math; Tol: Real from Standard)
    ---Purpose: Returns Standard_True if Sol is a zero of the function.
    --          Tol is the tolerance used in 3d space.
    returns Boolean from Standard
    is deferred;


end SurfCurvFuncInv;
