-- Created by: DAUTRY Philippe
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

--      	------------

---Version:	0.0
--Version	Date		Purpose
--		0.0	Feb 10 1997	Creation


class Data from DDF inherits Drawable3D from Draw

	---Purpose : Encapsulates a data framework in a drawable object

uses

    Data        from TDF,
    Interpretor from Draw,
    Display     from Draw

is


    Create  (aDF : Data from TDF)
    returns mutable Data from DDF;
    
    
    DrawOn (me; dis : in out Display);
    
    
    Copy (me) 
    returns mutable Drawable3D from Draw
    is redefined;

	
    Dump (me; S : in out OStream) 
    is redefined;


    DataFramework (me : mutable; aDF : Data from TDF);


    DataFramework (me)
    returns Data from TDF;
    

    Whatis (me; I : in out Interpretor from Draw)
    is redefined;

	
fields

    myDF : Data from TDF;

end Data;


