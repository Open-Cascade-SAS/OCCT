-- Created on: 2007-07-31
-- Created by: Sergey ZARITCHNY
-- Copyright (c) 2007-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class AsciiString from TDataStd inherits Attribute from TDF

        ---Purpose: Used to define an AsciiString attribute containing a TCollection_AsciiString

uses 
    Attribute         from TDF,
    Label             from TDF,
    GUID              from Standard,
    AsciiString       from TCollection,
    RelocationTable   from TDF

is
    ---Purpose: class methods
    --          =============

    GetID (myclass)   
        ---C++: return const & 
        ---Purpose: Returns the GUID of the attribute.  
    returns GUID from Standard;    

    Set (myclass; label : Label from TDF; string  : AsciiString from TCollection)
    ---Purpose: Finds, or creates an AsciiString attribute and sets the string.
    --          the AsciiString attribute is returned.
    returns AsciiString from TDataStd;
    
    ---Purpose: AsciiString methods
    --          ===================
    
    Create 
    returns mutable AsciiString from TDataStd;
    -- Constructor    
    
    Set (me : mutable; S : AsciiString from TCollection);
    -- Sets the ascii string <S>
    
    Get (me)
    returns AsciiString from TCollection;         
    -- Returns the AsciiString  <myString>
    ---C++: return const &
     
    IsEmpty(me) 
    returns Boolean from Standard;
    -- Returns True if the string of <me> contains zero characters. 
    
    ---Category: TDF_Attribute methods
    --           =====================
    
    ID (me)
        ---C++: return const & 
    returns GUID from Standard;

    Restore (me: mutable; with : Attribute from TDF);
    --  Restores the backuped content from <with> into this one. 
    
    NewEmpty (me)
    returns mutable Attribute from TDF;
    -- Returns an new empty AsciiString attribute. 
    
    Paste (me; into : mutable Attribute from TDF;
               RT   : mutable RelocationTable from TDF);    
    -- This method is used when copying an attribute from a source structure 
    -- into a target structure. 
    
    Dump(me; anOS : in out OStream from Standard)
        returns OStream from Standard
        is redefined;
        ---C++: return &
    -- This method dumps the attribute value into the stream
fields
    myString : AsciiString from TCollection; 
    
end AsciiString;
