-- Created on: 1991-10-03
-- Created by: Jean Claude VAUTHIER
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


package Geom2dConvert

        --- Purpose : 
        --  This package provides an implementation of algorithmes to do
        --  the conversion between equivalent geometric entities from 
        --  package Geom2d.
        --  It gives the possibility : 
        --   . to obtain the B-spline representation of bounded curves.
        --   . to split a B-spline curve into several B-spline curves 
        --     with some constraints of continuity,
        --   . to convert a B-spline curve into several Bezier curves
        --     or surfaces.
        --  All the geometric entities used in this package are bounded.
    	--   References :
        --  . Generating the Bezier Points of B-spline curves and surfaces
        --    (Wolfgang Bohm) CAGD volume 13 number 6 november 1981
        --  . On NURBS: A Survey  (Leslie Piegl) IEEE Computer Graphics and
        --    Application January 1991
        --  . Curve and surface construction using rational B-splines 
        --    (Leslie Piegl and Wayne Tiller) CAD Volume 19 number 9 november
        --    1987
        --  . A survey of curve and surface methods in CAGD (Wolfgang BOHM)
        --    CAGD 1 1984

uses Standard, TColStd, TColGeom2d,gp, Geom2d, Convert,GeomAbs

is


  class BSplineCurveKnotSplitting;
        --- Purpose :
        --  This algorithm searches the knot values corresponding to the 
        --  splitting of a given B-spline curve into  several arcs with
        --  the same continuity. The continuity order is given at the
        --  construction time. It is possible to compute the curve arcs
        --  corresponding to this splitting with the method of package 
        --  SplitBSplineCurve.



  class BSplineCurveToBezierCurve;
        --- Purpose : 
        --  This algorithm converts a B-spline curve from the package Geom
        --  into several Bezier curves.

  class CompCurveToBSplineCurve;
        --- Purpose : 
        --  This algorithm converts and concat sevral curve in a 
        --  B-spline curve.
  class  ApproxCurve;   
        ---Purpose : -- Convert a curve to BSpline  by Approximation
        --         
    
  SplitBSplineCurve (C               : BSplineCurve from Geom2d; 
                     FromK1, ToK2    : Integer;
                     SameOrientation : Boolean = Standard_True)
     returns mutable BSplineCurve from Geom2d
        --- Purpose : 
        --  This method computes the arc of B-spline curve between the two 
        --  knots FromK1 and ToK2.  If C is periodic the arc has the same
        --  orientation as C if SameOrientation = Standard_True.  
        --  If C is not periodic  SameOrientation is not used for the
        --  computation and C is oriented from the knot fromK1 to the
        --  knot toK2.  
        --  We just keep the local definition of C between the knots
        --  FromK1 and ToK2.  The returned B-spline curve has its first
        --  and last knots with a multiplicity equal to degree + 1, where
        --  degree is the polynomial degree of C.
        --  The indexes of the knots FromK1 and ToK2 doesn't include the
        --  repetition of multiple knots in their definition.
     raises OutOfRange from Standard,
        --- Purpose :  
        --  Raised if FromK1 or ToK2 are out of the bounds 
        --  [FirstUKnotIndex, LastUKnotIndex]
            DomainError from Standard;
      --- Purpose :  Raised if FromK1 = ToK2



  SplitBSplineCurve (C                   : BSplineCurve from Geom2d; 
                     FromU1, ToU2        : Real;
                     ParametricTolerance : Real;
                     SameOrientation     : Boolean = Standard_True)
     returns mutable BSplineCurve from Geom2d
        --- Purpose :
        --  This function computes the segment of B-spline curve between the 
        --  parametric values FromU1, ToU2.
        --  If C is periodic the arc has the same orientation as C if
        --  SameOrientation = True.  
        --  If C is not periodic SameOrientation is not used for the 
        --  computation and C is oriented fromU1 toU2. 
        --  If U1 and U2 and two parametric values we consider that 
        --  U1 = U2 if Abs (U1 - U2) <= ParametricTolerance and 
        --  ParametricTolerance must  be greater or equal to Resolution
        --  from package gp.
     raises DomainError from Standard;
        --- Purpose :
        --  Raised if FromU1 or ToU2 are out of the parametric bounds of the
        --  curve (The tolerance criterion is ParametricTolerance).
        --  Raised if Abs (FromU1 - ToU2) <= ParametricTolerance
        --  Raised if ParametricTolerance < Resolution from gp.



  CurveToBSplineCurve (C : Curve from Geom2d ;
    	    	       Parameterisation : ParameterisationType from Convert 
    	    	    	= Convert_TgtThetaOver2)
     returns mutable BSplineCurve from Geom2d
        --- Purpose : This function converts a non infinite curve from
        --   Geom into a  B-spline curve.  C must  be  an ellipse or a
        --   circle or a trimmed conic  or a trimmed  line or a Bezier
        --  curve or a trimmed  Bezier curve or a  BSpline curve or  a
        --  trimmed BSpline   curve  or an  Offset  curve or a  trimmed
        --  Offset curve.
         --  The returned B-spline is not periodic except if C is a 
        --  Circle or an Ellipse.
        --  ParameterisationType applies only if the curve is a Circle
        --  or an ellipse : 
        --      TgtThetaOver2,
    	--    TgtThetaOver2_1,
    	--    TgtThetaOver2_2,
    	--    TgtThetaOver2_3,
    	--    TgtThetaOver2_4,
	-- Purpose: this is the classical rational parameterisation
	--                    2
	--               1 - t
	--  cos(theta) = ------
	--                    2
	--               1 + t
	--                   
	--                 2t
	--  sin(theta) = ------
	--                     2
	--                1 + t
	--                   
	--  t = tan (theta/2)        
	-- 
	--  with TgtThetaOver2  the routine will compute the number of spans
	--  using the rule num_spans = [ (ULast - UFirst) / 1.2 ] + 1 
	--  with TgtThetaOver2_N, N  spans will be forced: an error will 
	--  be raized if (ULast - UFirst) >= PI and N = 1,
	--  ULast - UFirst >= 2 PI and N = 2
	--   
	-- QuasiAngular,
	--  here t is a rational function that approximates  
	--  theta ----> tan(theta/2).
	--  Neverthless the composing with above function yields exact
	--  functions whose square sum up to 1
	-- RationalC1 ;
	--  t is replaced by a polynomial function of u so as to grant
	--  C1 contiuity across knots.
	--  Exceptions
    	-- Standard_DomainError if the curve C is infinite.
    	-- Standard_ConstructionError:
    	-- -   if C is a complete circle or ellipse, and if
    	--   Parameterisation is not equal to
    	--   Convert_TgtThetaOver2 or to Convert_RationalC1, or
    	-- -   if C is a trimmed circle or ellipse and if
    	--   Parameterisation is equal to
    	--   Convert_TgtThetaOver2_1 and if U2 - U1 >
    	--   0.9999 * Pi where U1 and U2 are
    	--   respectively the first and the last parameters of the
    	--   trimmed curve (this method of parameterization
    	--   cannot be used to convert a half-circle or a
    	--   half-ellipse, for example), or
    	-- -   if C is a trimmed circle or ellipse and
    	--   Parameterisation is equal to
    	--   Convert_TgtThetaOver2_2 and U2 - U1 >
    	--   1.9999 * Pi where U1 and U2 are
    	--   respectively the first and the last parameters of the
    	--   trimmed curve (this method of parameterization
    	--   cannot be used to convert a quasi-complete circle or ellipse).
     raises DomainError;
    
       
       
    ConcatG1(ArrayOfCurves          : in out Array1OfBSplineCurve from TColGeom2d;
    	     ArrayOfToler           : in           Array1OfReal   from TColStd;
    	     ArrayOfConcatenated    : out  HArray1OfBSplineCurve from TColGeom2d;
	     ClosedFlag             : in   Boolean   from Standard ;
    	     ClosedTolerance        : in   Real                  from Standard);
    	--- Purpose : This Method concatenates G1 the ArrayOfCurves as far
    	--  as it is possible.
    	--  ArrayOfCurves[0..N-1]
    	--  ArrayOfToler contains the  biggest tolerance of the two
    	--               points shared by two consecutives curves.
    	--               Its dimension: [0..N-2]
    	--  ClosedTolerance     indicates if the ArrayOfCurves is closed.
    	--               In this case ClosedTolerance contains the biggest tolerance
    	--               of the two points which are at the closure.
    	--               Otherwise its value is 0.0
    
    
    ConcatC1(ArrayOfCurves          : in out Array1OfBSplineCurve from TColGeom2d;
    	     ArrayOfToler           : in           Array1OfReal   from TColStd;
	     ArrayOfIndices         : out        HArray1OfInteger from TColStd;
    	     ArrayOfConcatenated    : out  HArray1OfBSplineCurve from TColGeom2d;
	     ClosedFlag             : in   Boolean   from Standard ;
    	     ClosedTolerance        : in   Real                  from Standard);
    	--- Purpose : This Method concatenates C1 the ArrayOfCurves as far
    	--  as it is possible.
    	--  ArrayOfCurves[0..N-1]
    	--  ArrayOfToler contains the  biggest tolerance of the two
    	--               points shared by two consecutives curves.
    	--               Its dimension: [0..N-2]
    	--  ClosedTolerance     indicates if the ArrayOfCurves is closed.
    	--               In this case ClosedTolerance contains the biggest tolerance
    	--               of the two points which are at the closure.
    	--               Otherwise its value is 0.0
    	--               
        ConcatC1(ArrayOfCurves      : in out Array1OfBSplineCurve from TColGeom2d;
    	     ArrayOfToler           : in           Array1OfReal   from TColStd;
	     ArrayOfIndices         : out        HArray1OfInteger from TColStd;
    	     ArrayOfConcatenated    : out  HArray1OfBSplineCurve from TColGeom2d;
	     ClosedFlag             : in   Boolean   from Standard ;
    	     ClosedTolerance        : in   Real                  from Standard;
	     AngularTolerance       : in Real                  from Standard) ;
    	--- Purpose : This Method concatenates C1 the ArrayOfCurves as far
    	--  as it is possible.
    	--  ArrayOfCurves[0..N-1]
    	--  ArrayOfToler contains the  biggest tolerance of the two
    	--               points shared by two consecutives curves.
    	--               Its dimension: [0..N-2]
    	--  ClosedTolerance     indicates if the ArrayOfCurves is closed.
    	--               In this case ClosedTolerance contains the biggest tolerance
    	--               of the two points which are at the closure.
    	--               Otherwise its value is 0.0

    C0BSplineToC1BSplineCurve(BS              : in out BSplineCurve from Geom2d;
    	    	    	      Tolerance       : in Real from Standard);
    	--- Purpose :  This Method reduces as   far as it  is possible the
    	--  multiplicities of  the  knots of  the BSpline BS.(keeping  the geometry).
    	--  It returns a new BSpline which could still be C0.
    	--  tolerance is a geometrical tolerance


    C0BSplineToArrayOfC1BSplineCurve(BS        : in  BSplineCurve from Geom2d;
    	    	    	    	     tabBS     : out HArray1OfBSplineCurve from TColGeom2d;
				     Tolerance :in Real from Standard);
    	--- Purpose :This Method   reduces as far  as  it is possible  the
    	--  multiplicities  of  the knots  of the BSpline  BS.(keeping the geometry).
    	--  It returns an array of BSpline C1.
    	--  Tolerance is a geometrical tolerance
    
    C0BSplineToArrayOfC1BSplineCurve( BS               : in  BSplineCurve from Geom2d;
    	    	    	    	     tabBS             : out HArray1OfBSplineCurve from TColGeom2d;
				     AngularTolerance  : in Real from Standard;
				     Tolerance         : in Real from Standard) ;
    	--- Purpose :This Method   reduces as far  as  it is possible  the
    	--  multiplicities  of  the knots  of the BSpline  BS.(keeping the geometry).
    	--  It returns an array of BSpline C1.
    	--  tolerance is a geometrical tolerance
     

    
end Geom2dConvert;









