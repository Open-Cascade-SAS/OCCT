-- Created on: 1993-03-03
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Update:      fma


class Datum3D from PTopLoc inherits Persistent from Standard

	---Purpose: An  elementary local coordinate system. It  may be
	--          shared in the Database.

uses
    Trsf from gp

raises
    ConstructionError from Standard

is
    Create(T : Trsf from gp) returns Datum3D from PTopLoc
	---Purpose: Creates a   local coordinate  system    with   the
	--          transformation.  An   error   is raised  if    the
	--          transformation is not rigid.
	---Level: Internal 
    raises
    	ConstructionError from Standard;
	
    Transformation(me) returns Trsf from gp
    	---Purpose: Returns the transformation defining the coordinate
    	--          system.
	---Level: Internal 
    is static;
    
fields

    myTrsf : Trsf from gp;

end Datum3D;
