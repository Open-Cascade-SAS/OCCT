-- Created on: 1992-09-11
-- Created by: Stephan GARNAUD
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.





class EnvironmentIterator from OSD   

 ---Purpose: This allows consultation of every environment variable.
 --          There is no specific order of results.

uses Environment, Error, AsciiString from TCollection
raises OSDError

is
 Create returns EnvironmentIterator;
    ---Purpose: Instantiates Object as Iterator;
    ---Level: Public

 Destroy ( me : out );
	---C++: alias ~
	-- Only implemented on Windows NT system

 More (me : in out) returns Boolean  is static;
    ---Purpose: Returns TRUE if there are other environment variables.
    ---Level: Public

 Next (me : in out)  is static;
    ---Purpose: Sets the iterator to the next item.
    --          Returns the item value corresponding to the current
    --          position of the iterator.
    ---Level: Public

 Values (me : in out) returns Environment is static;
    ---Purpose: Returns the next environment variable found.
    ---Level: Public

 Failed (me) returns Boolean is static;
   ---Purpose: Returns TRUE if an error occurs
    ---Level: Public

 Reset (me : in out) is static;
   ---Purpose: Resets error counter to zero
    ---Level: Public
      
 Perror (me : in out)
   ---Purpose: Raises OSD_Error
    ---Level: Public
   raises OSDError is static ;

 Error (me) returns Integer is static ;
   ---Purpose: Returns error number if 'Failed' is TRUE.
    ---Level: Public

 fields
      myEnv        : Address;         -- Windows NT specific
      myCount      : Integer;         -- Count in list of variables
      myError      : Error;
end EnvironmentIterator from OSD;

