-- Created on: 1997-03-19
-- Created by: Yves FRICAUD
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Modified     by  SZY  Wed  Aug  18  1999


class Name from TNaming 
    
uses

    NameType         from TNaming,
    NamedShape       from TNaming,
    ListOfNamedShape from TNaming,
    ShapeEnum        from TopAbs,
    Orientation      from TopAbs,     
    Shape            from TopoDS,
    Label            from TDF, 
    LabelMap         from TDF,
    RelocationTable  from TDF 

is

    ---Category: Construction
    --           ============
    
    Create returns Name from TNaming;
    
    Type           (me : in out; aType : NameType  from TNaming);
    
    ShapeType      (me : in out; aType : ShapeEnum from TopAbs);
     
    Shape          (me : in out; theShape : Shape from TopoDS);
    
    Append         (me : in out; arg : NamedShape  from TNaming);
    
    StopNamedShape (me : in out; arg : NamedShape  from TNaming);
    
    Index          (me : in out; I : Integer   from Standard);  
     
    ContextLabel   (me : in out; theLab : Label from TDF);  
   
    Orientation    (me : in out; theOrientation : Orientation from TopAbs);
  

   ---Category: Queriyng
   --           ========

    Type (me) returns NameType from TNaming;
    
    ShapeType (me)  returns ShapeEnum from TopAbs;  
    
    Shape     (me)   returns Shape from TopoDS; 
    
    Arguments (me) returns ListOfNamedShape from TNaming;
    ---Purpose: 
    ---C++: return const&

    StopNamedShape (me) returns NamedShape from TNaming ;
    
    Index          (me) returns Integer    from Standard; 
         
    ContextLabel   (me) returns Label from TDF;  
    ---C++: return const&  

    Orientation    (me) returns Orientation from TopAbs;
    ---C++: inline
    ---C++: return const
    

    ---Category: Resolution
    --           ==========
    
    Solve(me; 
    	  aLab   : Label        from TDF;
    	  Valid  : LabelMap     from TDF)
    returns Boolean from Standard;		    	    	  
	    	
    Paste (me; 
    	   into : in out  Name from TNaming; 
    	   RT   : mutable RelocationTable from TDF);
    	    	
fields

    myType      : NameType         from TNaming;
    myShapeType : ShapeEnum        from TopAbs; 
    myArgs      : ListOfNamedShape from TNaming;
    myStop      : NamedShape       from TNaming;    
    myIndex     : Integer          from Standard; 
    myShape     : Shape            from TopoDS;
    myContextLabel : Label         from TDF;
    myOrientation  : Orientation   from TopAbs;
    
end Name;
