-- File:	Extrema_FuncExtCS.cdl
-- Created:	Mon Jan 22 17:06:01 1996
-- Author:	Laurent PAINNOT
--		<lpa@nonox>
---Copyright:	 Matra Datavision 1996


private class FuncExtCS from Extrema

 inherits FunctionSetWithDerivatives from math
    ---Purpose: Function to find extrema of the 
    --          distance between a curve and a surface.

uses    POnSurf           from Extrema,
    	POnCurv           from Extrema,
	SequenceOfPOnSurf from Extrema,
	SequenceOfPOnCurv from Extrema,
	SequenceOfReal    from TColStd,
	Pnt               from gp,
	Vector            from math,
	Matrix            from math,
	Curve             from Adaptor3d,
    	CurvePtr          from Adaptor3d,
	Surface           from Adaptor3d,
    	SurfacePtr        from Adaptor3d

raises  OutOfRange from Standard

is
    Create returns FuncExtCS;

    Create (C: Curve from Adaptor3d; S: Surface from Adaptor3d) returns FuncExtCS;
    	---Purpose:

    Initialize(me: in out; C: Curve from Adaptor3d; S: Surface from Adaptor3d)
    	---Purpose: sets the field mysurf of the function.
    is static;
    
    ------------------------------------------------------------
    -- In all next methods, an exception is raised if the fields 
    -- were not initialized.

    NbVariables (me) returns Integer;

    NbEquations (me) returns Integer;

    Value (me: in out; UV: Vector; F: out Vector) returns Boolean;
    	---Purpose: Calculation of Fi(U,V).

    Derivatives (me: in out; UV: Vector; DF: out Matrix)
    	returns Boolean;
    	---Purpose: Calculation of Fi'(U,V).

    Values (me: in out; UV: Vector; F: out Vector; DF: out Matrix)
    	returns Boolean;
    	---Purpose: Calculation of Fi(U,V) and Fi'(U,V).

    GetStateNumber (me: in out) returns Integer
    	---Purpose: Save the found extremum.
    	is redefined;

    NbExt (me) returns Integer;
    	---Purpose: Return the number of found extrema.

    SquareDistance (me; N: Integer) returns Real
    	---Purpose: Return the value of the Nth distance.
    	raises  OutOfRange;
	    	-- if N < 1 or N > NbExt(me).

    PointOnCurve (me; N: Integer) returns POnCurv
    	---Purpose: Returns the Nth extremum on C.
    	---C++: return const&
    	raises  OutOfRange;
	    	-- if N < 1 or N > NbExt(me).

    PointOnSurface (me; N: Integer) returns POnSurf
    	---Purpose: Return the Nth extremum on S.
    	---C++: return const&
    	raises  OutOfRange;
	    	-- if N < 1 or N > NbExt(me).

    Bidon1(me) returns SurfacePtr from Adaptor3d
    is static private;

    Bidon2(me) returns CurvePtr from Adaptor3d
    is static private;


fields
    myC    : CurvePtr from Adaptor3d;
    myS    : SurfacePtr from Adaptor3d;
    
    myP1   : Pnt from gp;
    myP2   : Pnt from gp;

    myt    : Real;          -- current value of U on C
    myU    : Real;          -- current value of U on S
    myV    : Real;          -- current value of V on S

    mySqDist:  SequenceOfReal    from TColStd;
    myPoint1: SequenceOfPOnCurv from Extrema;
    myPoint2: SequenceOfPOnSurf from Extrema;
    
    myCinit: Boolean;
    mySinit: Boolean;

end FuncExtCS;
