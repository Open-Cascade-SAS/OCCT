-- Created on: 1997-05-21
-- Created by: Christian CAILLET
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DescrReadWrite  from StepData    inherits ReadWriteModule  from StepData

uses Transient,
     SequenceOfAsciiString    from TColStd,
     AsciiString              from TCollection,
     Check                    from Interface,
     StepReaderData           from StepData,
     StepWriter               from StepData,
     Protocol                 from StepData

is

    Create (proto : Protocol from StepData) returns DescrReadWrite from StepData;

    CaseStep (me; atype : AsciiString from TCollection) returns Integer;

    CaseStep(me; types : SequenceOfAsciiString from TColStd) returns Integer
    	is redefined;

    IsComplex (me; CN : Integer) returns Boolean is redefined;

    StepType (me; CN : Integer) returns AsciiString from TCollection;
    ---C++ : return const &

    ComplexType (me; CN : Integer;
            	 types : in out SequenceOfAsciiString from TColStd)
        returns Boolean  is redefined;

    ReadStep (me; CN : Integer; data : StepReaderData; num : Integer;
               ach : in out Check; ent : mutable Transient);

    WriteStep (me; CN : Integer; SW : in out StepWriter; ent : Transient);

fields

    theproto : Protocol from StepData;

end DescrReadWrite;
