-- File:	BooleanOperations.cdl
-- Created:	Mon Jul 10 10:19:21 2000
-- Author:	Vincent DELOS
--		<vds@bulox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 2000


package BooleanOperations 

	---Purpose: package to perform  Boolean Operations between two
	--          solids called Object and Tool.

uses
    gp,
    Bnd,
    math,
    BRep,
    Geom,
    TopAbs,
    TopExp,
    TopoDS,
    TColStd,
    TopTools,
    Standard,
    TCollection,
    BRepAdaptor,
    GeomAdaptor, 
    IntTools, 
    BOPTColStd	     
is

    class AncestorsAndSuccessors;
    ---Purpose: to have a fast access in the class ShapesDataStructure
    --          to  the   upper and  lower  shapes of  a  given shape.
    --          e.g. : ancestors of an edge are the wires that contain
    --          it and its successors are the vertices that it holds.

 
--modified by NIZNHY-PKV Wed Feb  2 14:47:51 2005f     
--    class InterferenceResult;
    --Purpose: to describe a single interference between two shapes
    --          in the class ShapesDataStructure.
    
--    pointer PInterferenceResult to InterferenceResult from BooleanOperations;
    
--    class InterferencesList;
    --Purpose:  if the considered shape  S belongs to the Object this
    --          class  will  list all  the shapes   of the Tool  whose
    --          bounding boxes intersects with the  bounding box of S;
    --          if S belongs  to the Tool we  store all the shapes  of
    --          the Object whose intersection with S is not empty.
--modified by NIZNHY-PKV Wed Feb  2 14:48:00 2005t 

   class ShapeAndInterferences;
    ---Purpose: contains   a  shape S,  its  bounding  box,  its state
    --           according  to   the other  solid,   its ancestors and
    --          successors, all of   its interferences with the  other
    --          solid.
    
    pointer PShapeAndInterferences to ShapeAndInterferences from BooleanOperations;
    
    class ShapesDataStructure;
    ---Purpose:  contains all the  shapes of the  Object and Tool, all
    --          the  shapes created  by  intersection,  their bounding
    --          boxes,  their states, their ancestors  and successors,
    --          and all of their interferences.

    pointer PShapesDataStructure to ShapesDataStructure from BooleanOperations;
    
    class Explorer;
    ---Purpose: to find subshapes of a given shape of the Data Structure.

    class OnceExplorer;
    ---Purpose: the derived class of Explorer to find subshapes only once.

    --class BooleanOperations;
    ---Purpose: is to be  deferred with inherited classes Cut, Common,
    --          Fuse to perform boolean operations .


    enumeration StateOfShape is 
	---Purpose: State of a Shape of the 1st solid according to the
	--          2nd one.  State INOROUT is  used when we know that
	--           a shape  is  totally IN or   totally  OUT.  State
	--          INTERSECTED refers to a shape of the 1st solid cut
	--          by   the  2nd solid.   When a  shape has  a  state
	--          different  of  INTERSECTED or UNKNOWN   all of its
	--          subshapes have the same state.
	IN,
	OUT,
	ON,
	UNKNOWN,
	INOROUT,
	INTERSECTED
    end StateOfShape;
    
    enumeration KindOfInterference is 
	---Purpose: Interferences describe an intersection between two
	--          shapes. They  are classified following a hierarchy
	--          from the lower until the  upper.
    	SurfaceSurface,
	EdgeSurface,
	VertexSurface,
	EdgeEdge,
	VertexEdge,
	VertexVertex, 
	UnknownInterference  
    end StateOfShape;

    enumeration KindOfIntersection is
	---Purpose:  Describes the    fact   that  we    can  have  no
	--           intersection between two shapes, or   a true or a
	--          tangent one.
    	NoIntersection,
	TrueIntersection,
	SameDomain
    end KindOfIntersection;
    
    
    ------------------------
    -- For internal needs --
    ------------------------

    class AncestorsSeqAndSuccessorsSeq;

    class IndexedDataMapOfShapeAncestorsSuccessors instantiates IndexedDataMap from TCollection
    (Shape from TopoDS,AncestorsSeqAndSuccessorsSeq from BooleanOperations,ShapeMapHasher from TopTools);


     
    class IndexedDataMapOfShapeInteger instantiates 
    	    IndexedDataMap from TCollection(Shape          from TopoDS,
	    	    	    	    	    Integer        from Standard,
                                            ShapeMapHasher from TopTools);  

end BooleanOperations;



