-- File:        ManifoldSurfaceShapeRepresentation.cdl
-- Created:     Mon Dec  4 12:02:27 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWManifoldSurfaceShapeRepresentation from RWStepShape

	---Purpose : Read & Write Module for ManifoldSurfaceShapeRepresentation

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     ManifoldSurfaceShapeRepresentation from StepShape,
     EntityIterator from Interface

is

	Create returns RWManifoldSurfaceShapeRepresentation;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable ManifoldSurfaceShapeRepresentation from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : ManifoldSurfaceShapeRepresentation from StepShape);

	Share(me; ent : ManifoldSurfaceShapeRepresentation from StepShape; iter : in out EntityIterator);

end RWManifoldSurfaceShapeRepresentation;
