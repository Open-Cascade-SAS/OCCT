-- File:        LocalTime.cdl
-- Created:     Mon Dec  4 12:02:27 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWLocalTime from RWStepBasic

	---Purpose : Read & Write Module for LocalTime

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     LocalTime from StepBasic,
     EntityIterator from Interface

is

	Create returns RWLocalTime;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable LocalTime from StepBasic);

	WriteStep (me; SW : in out StepWriter; ent : LocalTime from StepBasic);

	Share(me; ent : LocalTime from StepBasic; iter : in out EntityIterator);

end RWLocalTime;
