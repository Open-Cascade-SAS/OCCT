-- File:	StepBasic_SourceItem.cdl
-- Created:	Wed May 10 15:09:05 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class SourceItem from StepBasic
inherits SelectType from StepData

    ---Purpose: Representation of STEP SELECT type SourceItem

uses
    HAsciiString from TCollection,
    SelectMember from StepData

is
    Create returns SourceItem from StepBasic;
	---Purpose: Empty constructor

    CaseNum (me; ent: Transient) returns Integer;
	---Purpose: Recognizes a kind of SourceItem select type
	--          1 -> HAsciiString from TCollection
	--          0 else
	
    NewMember (me) returns SelectMember is redefined;

    Identifier (me) returns HAsciiString from TCollection;
	---Purpose: Returns Value as Identifier (or Null if another type)

end SourceItem;
