-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ConversionBasedUnitAndLengthUnit from StepBasic inherits ConversionBasedUnit from StepBasic 

	--- This classe is an implementation of EXPRESS
	--  ANDOR Subtype Declaration.
uses

    LengthUnit from StepBasic, 
    DimensionalExponents from StepBasic, 
    HAsciiString from TCollection, 
    MeasureWithUnit from StepBasic
    
is

    Create returns ConversionBasedUnitAndLengthUnit;
	---Purpose: Returns a ConversionBasedUnitAndLengthUnit

    Init (me: mutable; aDimensions: DimensionalExponents from StepBasic)
    is redefined;

    Init (me: mutable; aDimensions: DimensionalExponents from StepBasic;
	               aName      : HAsciiString from TCollection;
	               aConversionFactor: MeasureWithUnit from StepBasic) is redefined;

    -- Specific Methods for Field Data Access --

    SetLengthUnit(me: mutable; aLengthUnit: LengthUnit);
    
    LengthUnit (me) returns LengthUnit;

    -- Specific Methods for ANDOR Field Data Access --

fields

    lengthUnit: LengthUnit from StepBasic;

end ConversionBasedUnitAndLengthUnit;
