-- Created on: 1995-06-06
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


package BRepApprox 

	---Purpose: This package provides services on intersection curves
	--          dealt by topological operations on BRep objects.
	--          Services are approximation services.


uses

    MMgt,
    TColStd,
    gp,
    GeomAbs,
    Adaptor3d,
    Geom,
    Geom2d,
    BRepAdaptor,
    IntSurf,
    ApproxInt
    
is

    generic class ApproxLineGen;
    
    class ApproxLine instantiates ApproxLineGen from BRepApprox
    	(BSplineCurve from Geom,
     	 BSplineCurve from Geom2d);

    generic class SurfaceToolGen;

    class SurfaceTool instantiates SurfaceToolGen from BRepApprox 
    	(Surface from BRepAdaptor);
    
    class Approx instantiates Approx from ApproxInt
    	(Surface                 from BRepAdaptor,
	 SurfaceTool             from BRepApprox,
	 Quadric                 from IntSurf,
	 QuadricTool             from IntSurf,
	 ApproxLine              from BRepApprox);

end BRepApprox;
