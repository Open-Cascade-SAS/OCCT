-- Created on: 1994-11-08
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class EdgeInterferenceTool from TopOpeBRepDS 

	---Purpose: a tool computing complex transition on Edge.

uses

    Orientation from TopAbs,
    CurveTransition from TopTrans,
    Interference from TopOpeBRepDS,
    Point from TopOpeBRepDS,
    Shape from TopoDS

is

    Create returns EdgeInterferenceTool from TopOpeBRepDS;
    
    Init(me : in out; 
         E : Shape from TopoDS; 
         I : Interference from TopOpeBRepDS)
    is static;
    
    Add(me : in out; 
        E : Shape from TopoDS;
        V : Shape from TopoDS;
        I : Interference from TopOpeBRepDS)
    is static;
    
    Add(me : in out; 
        E : Shape from TopoDS;
	P : Point from TopOpeBRepDS;
        I : Interference from TopOpeBRepDS)
    is static;
    
    Transition(me; I : mutable Interference from TopOpeBRepDS)
    is static;
    
fields
    
    myEdgeOrientation : Orientation from TopAbs;
    myEdgeOriented    : Integer from Standard;
    myTool            : CurveTransition from TopTrans;

end EdgeInterferenceTool from TopOpeBRepDS;
