-- Created on: 1996-11-21
-- Created by: Joelle CHAUVET
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Modified:	Wed Mar  5 09:45:42 1997
--    by:	Joelle CHAUVET
--              G1134 : new methods RealBounds and Constraints

class Surface from GeomPlate inherits Surface from Geom

    	---Purpose:
    	-- Describes the characteristics of plate surface objects
    	-- returned by BuildPlateSurface::Surface. These can be
    	-- used to verify the quality of the resulting surface before
    	-- approximating it to a Geom_BSpline surface generated
    	-- by MakeApprox. This proves necessary in cases where
    	-- you want to use the resulting surface as the support for
    	-- a shape. The algorithmically generated surface cannot
    	-- fill this function as is, and as a result must be converted first.
        
uses  Pnt     from gp,
      Vec     from gp,
      Trsf    from gp,
      GTrsf2d from gp,
      Shape   from GeomAbs,
      Curve   from Geom,
      Surface from Geom,
      Plate from Plate,
      Array2OfPnt2d from TColgp, 
      Array2OfPnt from TColgp,
      SequenceOfXY from TColgp 
      
raises RangeError          from Standard,
       NoSuchObject        from Standard,
       UndefinedDerivative from Geom,
       UndefinedValue      from Geom

is
      
       
    
  Create ( Surfinit : Surface from  Geom; Surfinter :  Plate  from  Plate)   
  returns  Surface  from  GeomPlate ;
  
  UReverse (me : mutable)
        ---Purpose :
        --  Reverses the U direction of parametrization of <me>. 
        --  The bounds of the surface are not modified.
    ;




  UReversedParameter (me; U : Real) returns Real
	---Purpose: Return the  parameter on the  Ureversed surface for
	--          the point of parameter U on <me>.
	--          
	--          me->UReversed()->Value(me->UReversedParameter(U),V)
	--          
	--          is the same point as
	--          
	--          me->Value(U,V)
    ;

  VReverse (me : mutable)
        ---Purpose :
        --  Reverses the V direction of parametrization of <me>. 
        --  The bounds of the surface are not modified.
    ;


  VReversedParameter (me; V : Real) returns Real
	---Purpose: Return the  parameter on the  Vreversed surface for
	--          the point of parameter V on <me>.
	--          
	--          me->VReversed()->Value(U,me->VReversedParameter(V))
	--          
	--          is the same point as
	--          
	--          me->Value(U,V)
    ;
    
  TransformParameters(me; U,V : in out Real; T : Trsf from gp)
	---Purpose: Computes the  parameters on the  transformed  surface for
	--          the transform of the point of parameters U,V on <me>.
	--          
	--          me->Transformed(T)->Value(U',V')
	--          
	--          is the same point as
	--          
	--          me->Value(U,V).Transformed(T)
	--          
	--          Where U',V' are the new values of U,V after calling
	--          
	--          me->TranformParameters(U,V,T)
	--          
	--          This methods does not change <U> and <V>
	--          
	--          It  can be redefined.  For  example on  the Plane,
	--          Cylinder, Cone, Revolved and Extruded surfaces.
    is redefined;
    
  ParametricTransformation(me; T : Trsf from gp) returns GTrsf2d from gp
	---Purpose: Returns a 2d transformation  used to find the  new
	--          parameters of a point on the transformed surface.
	--          
	--          me->Transformed(T)->Value(U',V')
	--          
	--          is the same point as
	--          
	--          me->Value(U,V).Transformed(T)
	--          
	--          Where U',V' are  obtained by transforming U,V with
	--          th 2d transformation returned by
	--          
	--          me->ParametricTransformation(T)
	--          
	--          This methods returns an identity transformation
	--          
	--          It  can be redefined.  For  example on  the Plane,
	--          Cylinder, Cone, Revolved and Extruded surfaces.
	--          
    is redefined;
    
  Bounds(me; U1, U2, V1, V2 : out Real)
        -- To get the parametric bounds of the surface.
        -- Returned values can be RealFirst or RealLast if the surface is
        -- infinite.
    ;

  IsUClosed (me)   returns Boolean
        ---Purpose : 
        --  Is the surface closed in the parametric direction U ?
        --  Returns True if for each parameter V  the distance
        --  between the point P (UFirst, V) and P (ULast, V) is
        --  lower or equal to Resolution from gp.  UFirst and ULast
        --  are the parametric bounds in the U direction.
    ;

  IsVClosed (me)   returns Boolean
        ---Purpose : 
        --  Is the surface closed in the parametric direction V ?
        --  Returns True if for each parameter U  the distance
        --  between the point P (U, VFirst) and  P (U, VLast) is
        --  lower or equal to Resolution from gp.  VFirst and VLast
        --  are the parametric bounds in the V direction.
    ;

  IsUPeriodic (me)   returns Boolean
        ---Purpose :
        --  Is the parametrization of a surface periodic in the 
        --  direction U ?
        --  It is possible only if the surface is closed in this
        --  parametric direction and if the following relation is
        --  satisfied : 
        --  for each parameter V the distance between the point 
        --  P (U, V)  and the point  P (U + T, V) is lower or equal
        --  to Resolution from package gp. T is the parametric period
        --  and must be a constant.
    ;
    
  UPeriod (me)  returns Real from Standard
	---Purpose: returns the Uperiod.
  raises
    	NoSuchObject from Standard
	---Purpose: raises if the surface is not uperiodic.
    is redefined;

  IsVPeriodic (me)   returns Boolean
        ---Purpose :
        --  Is the parametrization of a surface periodic in the 
        --  direction U ?
        --  It is possible only if the surface is closed in this
        --  parametric direction and if the following relation is
        --  satisfied : 
        --  for each parameter V the distance between the point 
        --  P (U, V)  and the point  P (U + T, V) is lower or equal
        --  to Resolution from package gp. T is the parametric period
        --  and must be a constant.
    ;

  VPeriod (me)    returns Real from Standard
	---Purpose: returns the Vperiod.
  raises
    	NoSuchObject from Standard
	---Purpose: raises if the surface is not vperiodic.
    is redefined;

  UIso (me; U : Real)  returns Curve
        ---Purpose : Computes the U isoparametric curve.
     	;

  VIso (me; V : Real)  returns Curve
        ---Purpose : Computes the V isoparametric curve.
    ;

  Continuity (me)   returns Shape from GeomAbs
        ---Purpose :
        --  Global Continuity of the surface in direction U and V : 
        --  C0 : only geometric continuity,
        --  C1 : continuity of the first derivative all along the surface,
        --  C2 : continuity of the second derivative all along the surface,
        --  C3 : continuity of the third derivative all along the surface,
        --  G1 : tangency continuity all along the surface,
        --  G2 : curvature continuity all along the surface,
        --  CN : the order of continuity is infinite.
        --- Example :
        --  If the surface is C1 in the V parametric direction and C2
        --  in the U parametric direction Shape = C1.
    ;

  IsCNu (me; N : Integer)   returns Boolean
        ---Purpose :
        --- Returns the order of continuity of the surface in the 
        --  U parametric direction. 
     raises RangeError
        ---Purpose : Raised if N < 0.
    ;

  IsCNv (me; N : Integer)   returns Boolean
        ---Purpose :
        --- Returns the order of continuity of the surface in the 
        --  V parametric direction. 
     raises RangeError
        ---Purpose : Raised if N < 0.
    ;

  D0 (me; U, V : Real; P : out Pnt)
        ---Purpose :
        --  Computes the point of parameter U,V on the surface.
     raises UndefinedValue
        ---Purpose : 
        --  Raised only for an "OffsetSurface" if it is not possible to
        --  compute the current point. 
    ;

  D1 (me; U, V : Real; P : out Pnt; D1U, D1V : out Vec)
        ---Purpose :
        --  Computes the point P and the first derivatives in the
        --  directions U and V at this point.
     raises UndefinedDerivative
        ---Purpose : Raised if the continuity of the surface is not C1.
    ;

  D2 (me; U, V : Real; P : out Pnt; D1U, D1V, D2U, D2V, D2UV : out Vec)
        ---Purpose :
        --  Computes the point P, the first and the second derivatives in
        --  the directions U and V at this point.
     raises UndefinedDerivative
        ---Purpose : Raised if the continuity of the surface is not C2.
    ;

  D3 (me; U, V : Real; P : out Pnt; 
      D1U, D1V, D2U, D2V, D2UV, D3U, D3V, D3UUV, D3UVV :out Vec)
        ---Purpose :
        --  Computes the point P, the first,the second and the third 
        --  derivatives in the directions U and V at this point.
     raises UndefinedDerivative
        ---Purpose : Raised if the continuity of the surface is not C2.
    ;

  DN (me; U, V : Real; Nu, Nv : Integer)   returns Vec
        ---Purpose ;
        --  Computes the derivative of order Nu in the direction U and Nv
        --  in the direction V at the point P(U, V).
     raises UndefinedDerivative,
        ---Purpose : 
        --  Raised if the continuity of the surface is not CNu in the U
        --  direction or not CNv in the V direction.
            RangeError
        ---Purpose : Raised if Nu + Nv < 1 or Nu < 0 or Nv < 0.
    ;  

  Copy (me)  returns like me; 

  Transform (me : mutable; T : Trsf) ;
        ---Purpose :
        --  Transformation of a geometric object. This tansformation 
        --  can be a translation, a rotation, a symmetry, a scaling
        --  or a complex transformation obtained by combination of
        --  the previous elementaries transformations.
        --  (see class Transformation of the package Geom).
  
   CallSurfinit (me) returns Surface from Geom;
   
   SetBounds (me : mutable ; Umin,Umax,Vmin,Vmax : in Real from Standard );         
   
   RealBounds(me; U1, U2, V1, V2 : out Real);
        -- To get the real parametric bounds of the surface.

   Constraints(me; Seq : out SequenceOfXY);
        -- To get the 2d constraints used by Plate


fields
    	mySurfinter : Plate from Plate; 
    	mySurfinit : Surface from  Geom;
    	myUmin,myUmax,myVmin,myVmax : Real from Standard;   

end;
