-- Created on: 1995-01-24
-- Created by: Mister rmi
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SensitiveSegment   from Select3D 
inherits SensitiveEntity from Select3D

	---Purpose: A framework to define sensitive zones along a segment
	--          One gives the 3D start and end point;
	--          the maximum number of 2D boxes given
	--          by this entity may be set by the user
	--          if the projected segment is 
	--          vertical or horizontal, one needs only 1 box. 
	--          for a pi/4 angle -> MaxNumber 2D boxes

uses
    Pnt              from gp,
    Pnt2d            from gp,
    Projector        from Select3D,
    Lin              from gp,
    EntityOwner      from SelectBasics,
    ListOfBox2d      from SelectBasics,
    PickArgs         from SelectBasics,
    Array1OfPnt2d    from TColgp,
    Box2d            from Bnd,
    Location         from TopLoc,
    Pnt              from Select3D,
    Pnt2d            from Select3D


is


    Create (OwnerId      : EntityOwner from SelectBasics;
    	    FirstP,LastP : Pnt from gp;
    	    MaxRect      : Integer = 1)
     returns mutable SensitiveSegment;
	---Purpose: Constructs the sensitive segment object defined by
    	-- the owner OwnerId, the points FirstP, LastP and the
    	-- maximum number of sensitive bounding boxes MaxRect.     
	    
    Set (me:mutable; MaxRect : Integer) is static;
    	---Purpose:  Sets the maximum number of sensitive rectangles MaxRect.
    	---C++: inline
    
    
    
    StartPoint (me : mutable ; aPt : Pnt from gp) is static;
    	---Level: Public 
    	---Purpose: changes the start Point of the Segment;
    	---C++: inline
    


    EndPoint (me : mutable ; aPt : Pnt from gp) is static;
    	---Level: Public 
    	---Purpose: changes the end point of the segment
    	---C++: inline
    
    
    StartPoint (me) returns Pnt from gp is static;
    	---Level: Public 
    	---Purpose: gives the 3D start Point of the Segment
    	---C++: inline
    
    
    EndPoint(me) returns Pnt from gp is static;
    	---Level: Public 
    	---Purpose: gives the 3D End Point of the Segment
    	---C++: inline 
	 
    StartPoint2d (me) returns Pnt2d from gp is static;
    	---Level: Public 
    	---Purpose: gives the 3D start Point of the Segment
    	---C++: inline
    
    
    EndPoint2d(me) returns Pnt2d from gp is static;
    	---Level: Public 
    	---Purpose: gives the 3D End Point of the Segment
    	---C++: inline
    
    Project (me:mutable;aProjector : Projector from Select3D) 
    is redefined virtual;
    	---Level: Public 
    	---Purpose: projection of the sensitive primitive in order to
    	--          get 2D boxes for the Sort Algorithm

    
    Areas   (me:mutable ; boxes : in out ListOfBox2d from SelectBasics) 
    is redefined static;
    	---Level: Public 
    	---Purpose: gives the 2D boxes which represent the segment in the 
    	--          selection process...

    GetConnected(me:mutable;aLocation: Location from TopLoc)
    returns SensitiveEntity from Select3D is redefined static;

    Matches (me : mutable;
             thePickArgs : PickArgs from SelectBasics;
             theMatchDMin, theMatchDepth : out Real from Standard)
    returns Boolean is redefined static;
    ---Level: Public
    ---Purpose: Checks whether the sensitive entity matches the picking
    -- detection area (close to the picking line).
    -- For details please refer to base class declaration.

    Matches (me  :mutable; 
             XMin,YMin,XMax,YMax : Real from Standard;
             aTol: Real from Standard) 
    returns Boolean
    is static;
     
    Matches (me  :mutable; 
             Polyline:Array1OfPnt2d from TColgp;
	     aBox:Box2d from Bnd;
             aTol: Real from Standard) 
    returns Boolean
    is redefined virtual;
    	---Level: Public 
    
        
    ComputeDepth(me;EyeLine: Lin from gp) 
    returns Real from Standard;

    MaxBoxes(me) returns Integer is redefined static;    
    	---Level: Public 
    	---Purpose:returns <mymaxrect>
    	---C++: inline

    Dump(me; S: in out OStream;FullDump : Boolean from Standard = Standard_True) is redefined virtual;

fields

    mymaxrect : Integer;
    mystart   : Pnt from Select3D;
    myend     : Pnt from Select3D;

    myprojstart : Pnt2d from Select3D; -- computed at convert time
    myprojend   : Pnt2d from Select3D; -- computed at convert time

end SensitiveSegment;








