-- Created on: 1991-01-10
-- Created by: Arnaud BOUZY
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


deferred class UnaryExpression from Expr

inherits GeneralExpression from Expr

uses NamedUnknown from Expr

raises OutOfRange from Standard, 
    NumericError from Standard,
    InvalidOperand from Expr

is

    Operand(me)
    ---Purpose: Returns the operand used
    ---C++: inline
    ---C++: return const &
    ---Level : Internal
    returns any GeneralExpression
    is static;

    SetOperand(me : mutable; exp : GeneralExpression)
    ---Purpose: Sets the operand used
    --          Raises InvalidOperand if <exp> contains <me>.
    ---Level : Internal
    raises InvalidOperand
    is static;
    
    CreateOperand(me : mutable; exp : GeneralExpression)
    ---Purpose: Sets the operand used during creation
    ---Level : Internal
    is static protected;
    
    NbSubExpressions(me)
    ---Purpose: Returns the number of sub-expressions contained
    --          in <me> ( >= 0)
    returns Integer
    is static;

    SubExpression(me; I : Integer)
    ---Purpose: Returns the <I>-th sub-expression of <me>.
    --          Raises OutOfRange if <I> > NbSubExpressions(me)
    ---C++: return const &
    returns any GeneralExpression
    raises OutOfRange
    is static;

    ContainsUnknowns(me) 
    ---Purpose: Does <me> contains NamedUnknown ?
    returns Boolean
    is static;

    Contains(me; exp : GeneralExpression)
    ---Purpose: Tests if <exp> is contained in <me>.
    returns Boolean
    is static;

    Replace(me : mutable ; var : NamedUnknown ; with : GeneralExpression)
    ---Purpose: Replaces all occurences of <var> with <with> in <me>
    --          Raises InvalidOperand if <with> contains <me>.
    raises InvalidOperand
    is static;
    
    Simplified(me) 
    ---Purpose: Returns a GeneralExpression after replacement of
    --          NamedUnknowns by an associated expression, and after
    --          values computation.
    returns any GeneralExpression
    raises NumericError;
    
fields

    myOperand : GeneralExpression;

end UnaryExpression;

