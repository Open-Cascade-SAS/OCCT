-- File:	RWStepBasic_RWProductDefinitionFormationRelationship.cdl
-- Created:	Sun Dec 15 10:59:25 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWProductDefinitionFormationRelationship from RWStepBasic

    ---Purpose: Read & Write tool for ProductDefinitionFormationRelationship

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    ProductDefinitionFormationRelationship from StepBasic

is
    Create returns RWProductDefinitionFormationRelationship from RWStepBasic;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : ProductDefinitionFormationRelationship from StepBasic);
	---Purpose: Reads ProductDefinitionFormationRelationship

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: ProductDefinitionFormationRelationship from StepBasic);
	---Purpose: Writes ProductDefinitionFormationRelationship

    Share (me; ent : ProductDefinitionFormationRelationship from StepBasic;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWProductDefinitionFormationRelationship;
