-- Created on: 1994-07-12
-- Created by: Bruno DUMORTIER
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class MakePipe from BRepOffsetAPI inherits MakeSweep from BRepPrimAPI

    	---Purpose: Describes functions to build pipes.
    	-- A pipe is built a basis shape (called the profile) along
    	-- a wire (called the spine) by sweeping.
    	-- The profile must not contain solids.
    	-- A MakePipe object provides a framework for:
    	-- - defining the construction of a pipe,
    	-- - implementing the construction algorithm, and
    	-- - consulting the result.
    	-- Warning
    	-- The MakePipe class implements pipe constructions
    	-- with G1 continuous spines only.
uses
    Pipe        from BRepFill,
    Wire        from TopoDS,
    Shape       from TopoDS,
    Edge        from TopoDS,
    ListOfShape from TopTools

is
 
    
    Create( Spine   : Wire  from TopoDS;
    	    Profile : Shape from TopoDS )
	---Purpose: Constructs a pipe by sweeping the shape Profile along
    	-- the wire Spine.The angle made by the spine with the profile is
    	-- maintained along the length of the pipe.
    	-- Warning
    	-- Spine must be G1 continuous; that is, on the connection
    	-- vertex of two edges of the wire, the tangent vectors on
    	-- the left and on the right must have the same direction,
    	-- though not necessarily the same magnitude.
        -- Exceptions
    	-- Standard_DomainError if the profile is a solid or a
    	-- composite solid.
    returns MakePipe from BRepOffsetAPI;
    

    Pipe(me) returns Pipe from BRepFill
	---C++: return const &
	---Level: Advanced
    is static;


    Build(me : in out)
    is redefined;
	---Purpose: Builds the resulting shape (redefined from MakeShape).
	---Level: Public    


    FirstShape (me : in out)
    ---Purpose: Returns the  TopoDS  Shape of the bottom of the prism.
    returns Shape from TopoDS;


    LastShape (me : in out)
    ---Purpose: Returns the TopoDS Shape of the top of the prism.
    returns Shape from TopoDS;


    Generated (me: in out; SSpine, SProfile : Shape from TopoDS)
        ---Level: Public
    returns Shape from TopoDS;


fields

    myPipe : Pipe from BRepFill;

end MakePipe; 
