-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SurfaceModel from StepShape inherits SelectType from StepData

	-- <SurfaceModel> is an EXPRESS Select Type construct translation.
	-- it gathers : ShellBasedSurfaceModel, FaceBasedSurfaceModel
	-- Rev4 : only remains ShellBasedSurfaceModel

uses

	ShellBasedSurfaceModel
--	FaceBasedSurfaceModel
is

	Create returns SurfaceModel;
	---Purpose : Returns a SurfaceModel SelectType

	CaseNum (me; ent : Transient) returns Integer;
	---Purpose: Recognizes a SurfaceModel Kind Entity that is :
	--        1 -> ShellBasedSurfaceModel
	--        2 -> FaceBasedSurfaceModel
	--        0 else

	ShellBasedSurfaceModel (me) returns any ShellBasedSurfaceModel;
	---Purpose : returns Value as a ShellBasedSurfaceModel (Null if another type)

end SurfaceModel;

