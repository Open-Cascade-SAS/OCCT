-- Created by: DAUTRY Philippe
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

--      	------------------

---Version:	0.0
--Version	Date		Purpose
--		0.0	Feb  4 1998	Creation


class Shape1 from PTopoDS inherits Storable from Standard

    ---Purpose: The PTopoDS_Shape1 is the Persistent view of a TopoDS_Shape.
    --          
    --  a  Shape1 contains :
    --          
    --          - a reference to a TShape1.
    --          
    --          - a Location  to put the TShape1 in  a local coordinate
    --          system.
    --          
    --          - an Orientation.
    --          
    --          It inherits from ExternShareable, so that it can be shared
    --          by other objects located outside the container.
    
uses

    Orientation   from TopAbs,
    TShape1       from PTopoDS,
    Location      from PTopLoc
    
is
    Create returns Shape1 from PTopoDS;
    ---Level: Internal 

    Nullify(me : in out)
    is static;

    TShape(me) returns any TShape1 from PTopoDS
    ---Level: Internal 
    ---C++: return const &
    is static;

    TShape(me : in out; T : TShape1 from PTopoDS)
    ---Level: Internal 
    is static;

    Location(me) returns Location from PTopLoc
    ---Level: Internal 
    is static;
	
    Location(me : in out; L : Location from PTopLoc)
    ---Level: Internal 
    is static;
	
    Orientation(me) returns Orientation from TopAbs
    ---Level: Internal 
    is static;

    Orientation(me: in out; O : Orientation from TopAbs)
    ---Level: Internal 
    is static;
    
fields

    myTShape   : TShape1     from PTopoDS;
    myLocation : Location    from PTopLoc;
    myOrient   : Orientation from TopAbs;

end Shape1;
