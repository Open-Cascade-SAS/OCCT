-- Created on: 2001-12-28
-- Created by: Andrey BETENEV
-- Copyright (c) 2001-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1

class ConnectedEdgeSet from StepShape
inherits TopologicalRepresentationItem from StepShape

    ---Purpose: Representation of STEP entity ConnectedEdgeSet

uses
    HAsciiString from TCollection,
    HArray1OfEdge from StepShape

is
    Create returns ConnectedEdgeSet from StepShape;
	---Purpose: Empty constructor

    Init (me: mutable; aRepresentationItem_Name: HAsciiString from TCollection;
                       aCesEdges: HArray1OfEdge from StepShape);
	---Purpose: Initialize all fields (own and inherited)

    CesEdges (me) returns HArray1OfEdge from StepShape;
	---Purpose: Returns field CesEdges
    SetCesEdges (me: mutable; CesEdges: HArray1OfEdge from StepShape);
	---Purpose: Set field CesEdges

fields
    theCesEdges: HArray1OfEdge from StepShape;

end ConnectedEdgeSet;
