-- Created on: 2008-05-21
-- Created by: Vladislav ROMASHKO
-- Copyright (c) 2008-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class BooleanOperation from Voxel

    ---Purpose: Boolean operations (fuse, cut)
    --          for voxels of the same dimension.

uses

    DS from Voxel,
    BoolDS from Voxel,
    ColorDS from Voxel,
    FloatDS from Voxel

is

    Create
    ---Purpose: An empty constructor.
    returns BooleanOperation from Voxel;

    
    ---Category: Fusion
    --           ======

    Fuse(me;
    	 theVoxels1 : in out BoolDS from Voxel;
    	 theVoxels2 : in     BoolDS from Voxel)
    ---Purpose: Fuses two cubes of voxels.
    --          It modifies the first cube of voxels.
    --          It returns false in case of different dimension of the cube,
    --          different number of voxels.
    returns Boolean from Standard;

    Fuse(me;
    	 theVoxels1 : in out ColorDS from Voxel;
    	 theVoxels2 : in     ColorDS from Voxel)
    ---Purpose: Fuses two cubes of voxels.
    --          It modifies the first cube of voxels.
    --          It returns false in case of different dimension of the cube,
    --          different number of voxels.
    --          It summerizes the value of corresponding voxels and puts the result to theVoxels1.
    --          If the result exceeds 15 or becomes greater, it keeps 15.
    returns Boolean from Standard;

    Fuse(me;
    	 theVoxels1 : in out FloatDS from Voxel;
    	 theVoxels2 : in     FloatDS from Voxel)
    ---Purpose: Fuses two cubes of voxels.
    --          It modifies the first cube of voxels.
    --          It returns false in case of different dimension of the cube,
    --          different number of voxels.
    --          It summerizes the value of corresponding voxels and puts the result to theVoxels1.
    returns Boolean from Standard;

    
    ---Category: Cut
    --           ===

    Cut(me;
    	theVoxels1 : in out BoolDS from Voxel;
    	theVoxels2 : in     BoolDS from Voxel)
    ---Purpose: Cuts two cubes of voxels.
    --          It modifies the first cube of voxels.
    --          It returns false in case of different dimension of the cube,
    --          different number of voxels.
    returns Boolean from Standard;
    
    Cut(me;
    	theVoxels1 : in out ColorDS from Voxel;
    	theVoxels2 : in     ColorDS from Voxel)
    ---Purpose: Cuts two cubes of voxels.
    --          It modifies the first cube of voxels.
    --          It returns false in case of different dimension of the cube,
    --          different number of voxels.
    --          It subtracts the value of corresponding voxels and puts the result to theVoxels1.
    returns Boolean from Standard;

    Cut(me;
    	theVoxels1 : in out FloatDS from Voxel;
    	theVoxels2 : in     FloatDS from Voxel)
    ---Purpose: Cuts two cubes of voxels.
    --          It modifies the first cube of voxels.
    --          It returns false in case of different dimension of the cube,
    --          different number of voxels.
    --          It subtracts the value of corresponding voxels and puts the result to theVoxels1.
    returns Boolean from Standard;

    
    ---Category: Private area
    --           ============
    
    Check(me;
    	  theVoxels1 : DS from Voxel;
    	  theVoxels2 : DS from Voxel)
    returns Boolean from Standard
    is private;
    
end BooleanOperation;
