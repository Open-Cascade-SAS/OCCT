-- Created on: 1992-03-26
-- Created by: Laurent BUCHARD
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




private class PConicTool from IntCurve

	---Purpose: Implementation of the ParTool from IntImpParGen
	--          for conics of gp, using the class PConic from IntCurve.

        ---Level: Internal

uses Pnt2d    from gp,
     Vec2d    from gp,
     Lin2d    from gp,
     XY       from gp,
     PConic from IntCurve

is


    EpsX (myclass; C: PConic)
    	--Purpose: Tolerance used by mathematical algorithms 
    	--         usually about 1e-10
    	returns Real from Standard;


    NbSamples(myclass; C: PConic)
    	--Purpose: returns the number of samples on the parametric curve
    	returns Integer from Standard;

    NbSamples(myclass; C: PConic; U0,U1: Real from Standard)
    	--Purpose: returns the number of samples on the parametric curve
    	returns Integer from Standard;
 

    Value (myclass; C: PConic from IntCurve; X: Real from Standard)
    	--Purpose: Returns the   geometric  point which  lies   at the
    	--         parameter x on the parametric curve.
    	returns Pnt2d from gp;


    D1 (myclass; C: PConic from IntCurve; U: Real from Standard ; 
                 P: out Pnt2d; T: out Vec2d);
    	--Purpose: Computes the Value, First and  Second Derivative at
    	--         the parameter U on the curve.


    D2 (myclass; C: PConic from IntCurve; U: Real from Standard ; 
                 P: out Pnt2d; T,N: out Vec2d);
		 
    	--Purpose: Computes the Value, First and  Second Derivative at
    	--         the parameter U on the curve.
	 		 
end PConicTool;









