-- File:	StepAP203_StartWork.cdl
-- Created:	Fri Nov 26 16:26:40 1999 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0
-- Copyright:	Matra Datavision 1999

class StartWork from StepAP203
inherits ActionAssignment from StepBasic

    ---Purpose: Representation of STEP entity StartWork

uses
    Action from StepBasic,
    HArray1OfWorkItem from StepAP203

is
    Create returns StartWork from StepAP203;
	---Purpose: Empty constructor

    Init (me: mutable; aActionAssignment_AssignedAction: Action from StepBasic;
                       aItems: HArray1OfWorkItem from StepAP203);
	---Purpose: Initialize all fields (own and inherited)

    Items (me) returns HArray1OfWorkItem from StepAP203;
	---Purpose: Returns field Items
    SetItems (me: mutable; Items: HArray1OfWorkItem from StepAP203);
	---Purpose: Set field Items

fields
    theItems: HArray1OfWorkItem from StepAP203;

end StartWork;
