-- Created on: 1993-07-21
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class Command from BRepBuilderAPI 

	---Purpose: Root class for all commands in BRepBuilderAPI.  
	--          
	--          Provides :
	--          
	--          * Managements of the notDone flag.
	--          
	--          * Catching of exceptions (not implemented).
	--          
	--          * Logging (not implemented).

raises
    NotDone from StdFail
    
is
    Delete(me:out) is virtual;
    ---C++: alias "Standard_EXPORT virtual ~BRepBuilderAPI_Command(){Delete() ; }"
    
    Initialize;
	---Purpose: Set done to False.
    
    IsDone(me) returns Boolean is virtual;
	---Level: Public
    
    Done(me : in out)
	---Purpose: Set done to true.
	---Level: Public
    is static protected;
    
    NotDone(me : in out)
	---Purpose: Set done to false.
	---Level: Public
    is static protected;
    
    
    
    Check(me)
	---Purpose: Raises NotDone if done is false.
	---Level: Public
    raises NotDone from StdFail
    is static;

fields 
    myDone : Boolean;

end Command;
