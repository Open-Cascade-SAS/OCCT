-- Created on: 1991-10-09
-- Created by: Michel CHAUVAT
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

generic class   ExtPSOfRev from Extrema (SurfaceOfRevolution as any;
    	    	    	    	    	 Tool                as any ; -- as ToolSurfaceOfRevolution(SurfaceOfRevolution)
					 Curve               as any;
					 ToolCurve           as any; -- as ToolCurve(Curve)
					 TheExtPC            as any
					)
    	---Purpose: It calculates all the extremum distances
    	--          between a point and a surface.
    	--          These distances can be minimum or maximum.

uses   	POnSurf           from Extrema,
    	SequenceOfPOnSurf from Extrema,
    	Pnt               from gp,
    	SequenceOfReal    from TColStd
	
raises  NotDone    from StdFail,
    	OutOfRange from Standard

is
    Create (P: Pnt; S: SurfaceOfRevolution; Tol: Real; NbV: Integer;
    	    TolV: Real) returns ExtPSOfRev;
      	---Purpose: It calculates all the distances between a point 
      	--          and a surface of revolution.
      	--          Tol is used to test if the point is on the axis.
      	--          NbV and TolV are used to compute the extrema on a 
      	--          meridian (see ExtPC.cdl).

    IsDone (me) returns Boolean
    	---Purpose: Returns True if the distances are found.
    	is static;
    
    NbExt (me) returns Integer
    	---Purpose: Returns the number of extremum distances.
    	raises  NotDone from StdFail
	    	-- if IsDone(me)=False.
    	is static;

    SquareDistance (me; N: Integer) returns Real
    	---Purpose: Returns the value of the Nth resulting square distance.
    	raises  NotDone from StdFail,
    	    	-- if IsDone(me)=False.
    	        OutOfRange
		-- if N < 1 or N > NbPoints(me).
    	is static;

    Point (me; N: Integer) returns POnSurf
        ---C++: return const &
    	---Purpose: Returns the point of the Nth resulting distance.
    	raises  NotDone from StdFail,
    	    	-- if IsDone(me)=False.
    	        OutOfRange
		-- if N < 1 or N > NbPoints(me).
    	is static;

fields
    myDone : Boolean;
    mySqDist: SequenceOfReal from TColStd;
    myPoint: SequenceOfPOnSurf from Extrema;

end ExtPSOfRev;
