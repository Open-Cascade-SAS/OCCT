-- Created on: 1994-07-06
-- Created by: Laurent PAINNOT
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

generic class GLocateExtCC2d from Extrema (Curve1    as any;
    	    	    	    	    	   Tool1     as any;
					   Curve2    as any;
					   Tool2     as any)
					
    	---Purpose: It calculates the distance between two curves with
    	--          a close point; these distances can be maximum or 
    	--          minimum.

uses   POnCurv2d from Extrema,
       Pnt2d     from gp,
       Vec2d     from gp,
       HArray1OfPnt2d from TColgp

raises  DomainError  from Standard,
    	NotDone      from StdFail


    class LCCache2d instantiates CurveCache from Extrema (Curve1, Pnt2d from gp, HArray1OfPnt2d from TColgp);

    class ELCC2d    instantiates GenExtCC      from Extrema
        (Curve1,
         Tool1,
         Curve2,
         Tool2,
         LCCache2d,
         HArray1OfPnt2d from TColgp,
         POnCurv2d,
         Pnt2d,
         Vec2d);


    class LocECC2d    instantiates GenLocateExtCC      from Extrema
    	(Curve1,
	 Tool1,
	 Curve2,
	 Tool2,
         POnCurv2d,
         Pnt2d,
         Vec2d);


is
    Create (C1: Curve1; C2: Curve2; U0,V0: Real)
    	returns GLocateExtCC2d
    	---Purpose: Calculates the distance with a close point. The
    	--          close point is defined by a parameter value on each 
    	--          curve.
    	--          The function F(u,v)=distance(C1(u),C2(v)) has an 
    	--          extremun when gradient(f)=0. The algorithm searchs
    	--          the zero near the close point.
    	raises  DomainError;
    	    	-- if U0 and V0 are outside the definition ranges of the 
    	    	-- curves.
    
    IsDone (me) returns Boolean
    	---Purpose: Returns True if the distance is found.
    	is static;

    SquareDistance (me) returns Real
    	---Purpose: Returns the value of the extremum square distance.
	raises  NotDone from StdFail
	    	-- if IsDone(me)=False.
    	is static;

    Point (me; P1,P2: out POnCurv2d)
    	---Purpose: Returns the points of the extremum distance. 
    	--          P1 is on the first curve, P2 on the second one.
    	raises  NotDone from StdFail
    	    	-- if IsDone(me)=False.
    	is static;

fields
    myDone  : Boolean;
    mySqDist: Real;
    myPoint1: POnCurv2d;
    myPoint2: POnCurv2d;

end GLocateExtCC2d;
