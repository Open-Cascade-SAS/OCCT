-- Created on: 1993-08-26
-- Created by: Christian CAILLET
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



deferred class Modifier  from IFSelect  inherits GeneralModifier

    ---Purpose : This class gives a frame for Actions which can work globally
    --           on a File once completely defined (i.e. afterwards)
    --           
    --           Remark : if no Selection is set as criterium, the Modifier is
    --           set to work and should consider all the content of the Model
    --           produced.

uses CString, InterfaceModel, CopyTool, Protocol from Interface, ContextModif

is

    Initialize (maychangegraph : Boolean);
    ---Purpose : Calls inherited Initialize, transmits to it the information
    --           <maychangegraph>

    Perform (me; ctx  : in out ContextModif;
    	     target   : mutable InterfaceModel;
    	     protocol : Protocol from Interface;
    	     TC       : in out CopyTool) is deferred;
    ---Purpose : This deferred method defines the action specific to each class
    --           of Modifier. It is called by a ModelCopier, once the Model
    --           generated and filled. ModelCopier has already checked the
    --           criteria (Dispatch, Model Rank, Selection) before calling it.
    --           
    --           <ctx> detains informations about original data and selection.
    --           The result of copying, on which modifications are to be done,
    --           is <target>.
    --           <TC> allows to run additional copies as required
    --           
    --           In case of Error, use methods CCheck from the ContextModif
    --           to aknowledge an entity Check or a Global Check with messages

end Modifier;
