-- File:	QAAMINO.cdl
-- Created:	Thu Jul 18 16:58:18 2002
-- Author:	QA Admin
--		<qa@umnox.nnov.matra-dtv.fr>
---Copyright:	 Matra Datavision 2002

package QAAMINO
     uses Draw
is
    
    Commands(DI : in out Interpretor from Draw);
end;
