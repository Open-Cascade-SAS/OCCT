-- Created on: 1998-08-04
-- Created by: Christian CAILLET
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class AutoDesignReferencingItem from StepAP214 inherits SelectType from StepData

	-- <AutoDesignReferencingItem> is an EXPRESS Select Type construct translation.
	-- it gathers : 
--    (approval,
--    document_relationship,
--    externally_defined_representation,
--    mapped_item,
--    material_designation,
--    presentation_area,
--    presentation_view,
--    product_category,
--    product_definition,
--    product_definition_relationship,
--    property_definition,
--    representation,
--    representation_relationship,
--    shape_aspect);

uses

     Approval from StepBasic,
     DocumentRelationship from StepBasic,
     ExternallyDefinedRepresentation from StepRepr,
     MappedItem from StepRepr,
     MaterialDesignation from StepRepr,
     PresentationArea from StepVisual,
     PresentationView from StepVisual,
     ProductCategory from StepBasic,
     ProductDefinition from StepBasic,
     ProductDefinitionRelationship from StepBasic,
     PropertyDefinition from StepRepr,
     Representation from StepRepr,
     RepresentationRelationship from StepRepr,
     ShapeAspect from StepRepr

is

	Create returns AutoDesignReferencingItem;
	---Purpose : Returns a AutoDesignReferencingItem SelectType

	CaseNum (me; ent : Transient) returns Integer;
	---Purpose: Recognizes a AutoDesignReferencingItem Kind Entity that is :
	-- 1     Approval from StepBasic,
	-- 2     DocumentRelationship from StepBasic,
	-- 3     ExternallyDefinedRepresentation from StepRepr,
	-- 4     MappedItem from StepRepr,
	-- 5     MaterialDesignation from StepRepr,
	-- 6     PresentationArea from StepVisual,
	-- 7     PresentationView from StepVisual,
	-- 8     ProductCategory from StepBasic,
	-- 9     ProductDefinition from StepBasic,
	-- 10     ProductDefinitionRelationship from StepBasic,
	-- 11     PropertyDefinition from StepBasic,
	-- 12     Representation from StepRepr,
	-- 13     RepresentationRelationship from StepRepr,
	-- 14     ShapeAspect from StepRepr
	--        0 else


    Approval (me) returns Approval from StepBasic;
    DocumentRelationship (me) returns DocumentRelationship from StepBasic;
    ExternallyDefinedRepresentation (me) returns ExternallyDefinedRepresentation from StepRepr;
    MappedItem (me) returns MappedItem from StepRepr;
    MaterialDesignation (me) returns MaterialDesignation from StepRepr;
    PresentationArea (me) returns PresentationArea from StepVisual;
    PresentationView (me) returns PresentationView from StepVisual;
    ProductCategory (me) returns ProductCategory from StepBasic;
    ProductDefinition (me) returns ProductDefinition from StepBasic;
    ProductDefinitionRelationship (me) returns ProductDefinitionRelationship from StepBasic;
    PropertyDefinition (me) returns PropertyDefinition from StepRepr;
    Representation (me) returns Representation from StepRepr;
    RepresentationRelationship (me) returns RepresentationRelationship from StepRepr;
    ShapeAspect (me) returns ShapeAspect from StepRepr;

end AutoDesignReferencingItem;
