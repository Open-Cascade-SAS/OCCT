-- File:	MXCAFDoc_CentroidRetrievalDriver.cdl
-- Created:	Mon Sep 11 15:14:09 2000
-- Author:	data exchange team
--		<det@doomox>
---Copyright:	 Matra Datavision 2000


class CentroidRetrievalDriver from MXCAFDoc inherits  ARDriver from MDF 

	---Purpose: 

uses
    RRelocationTable from MDF,
    Attribute        from PDF,
    Attribute        from TDF,
    MessageDriver    from CDM

is
--    Create -- Version 0
--    returns mutable CentroidRetrievalDriver from MXCAFDoc;
    Create (theMsgDriver : MessageDriver from CDM)
    returns mutable CentroidRetrievalDriver from MXCAFDoc;
    
    VersionNumber(me) returns Integer from Standard;
    ---Purpose: Returns the version number from which the driver
    --          is available: 0.

    SourceType(me) returns Type from Standard;
    ---Purpose: Returns the type: XCAFDoc_Centroid

    NewEmpty (me)  returns mutable Attribute from TDF;

    Paste(me;
    	  Source     :         Attribute from PDF;
    	  Target     : mutable Attribute from TDF;
    	  RelocTable : RRelocationTable from MDF);

end CentroidRetrievalDriver;
