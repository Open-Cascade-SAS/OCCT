-- Created on: 1999-06-17
-- Created by: Vladislav ROMASHKO
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Function from PFunction inherits Attribute from PDF 

uses 
     
    Attribute from PDF, 
    GUID      from Standard 

is

    Create returns mutable Function from PFunction;
        
    SetDriverGUID(me : mutable; driverGUID : GUID from Standard);

    GetDriverGUID(me) returns GUID from Standard;

    GetFailure(me) returns Integer from Standard;
    
    SetFailure(me : mutable; mode : Integer from Standard);

fields

    myDriverGUID  : GUID     from Standard;
    myFailure     : Integer  from Standard;

end Function;
 
