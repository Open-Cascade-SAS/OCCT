-- Created on: 1993-03-23
-- Created by: BBL
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Modified:	02-06-98 : FMN ; Suppression appel Clear (deja fait dans ALienData)

class EuclidAlienImage from AlienImage inherits AlienUserImage from AlienImage

	---Version: 0.0

	---Purpose: This class defines an Euclid Alien image.
	---Keywords:
	---Warning:
	---References:

uses
	File 			from OSD,
	AsciiString 		from TCollection,
	ColorImage 		from Image,
	PseudoColorImage 	from Image,
	Image			from Image,
	EuclidAlienData 	from AlienImage

is
	Create returns mutable EuclidAlienImage from AlienImage;

	Clear( me : in out mutable) ;
	---Level: Public
	---Purpose: Frees memory allocated by EuclidAlienImage

	ToImage( me : in immutable ) 
	  returns mutable Image from Image ;
	---Level: Public
	---Purpose : Converts a EuclidAlienImage object to a Image object.

	FromImage( me : in out mutable ; anImage : in Image from Image ) ;
	---Level: Public
	---Purpose : converts a Image object to a EuclidAlienImage object.

	Read ( me : in out mutable; afile : in out File from OSD )
	  returns Boolean from Standard ;
	---Purpose: Reads content of a EuclidAlienImage object
	--          from a file .
	--          Returns True if file is a Euclid file .

	Write( me : in immutable; afile : in out File from OSD )
	  returns Boolean from Standard ;
	---Purpose: Writes content of a EuclidAlienImage object
	--          to a file .

fields
	myData : EuclidAlienData from AlienImage ;

end ;
 
