-- Created on: 1997-09-30
-- Created by: Roman BORISOV
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class CurveOnSurface from Approx 

	---Purpose: 
    ---Purpose: Approximation of   curve on surface

uses     
         Surface         from   Geom,
         HCurve2d          from   Adaptor2d, 
	 HSurface    from  Adaptor3d, 
         BSplineCurve    from   Geom,
         BSplineCurve    from   Geom2d,  
	 Shape  from  GeomAbs   
	  
raises  OutOfRange        from Standard,
        ConstructionError from Standard

is  

Create (C2D  :  HCurve2d    from  Adaptor2d;
	  Surf :  HSurface  from  Adaptor3d; 
	     First, 
	     Last, 		      
             Tol  :  Real; 
	     Continuity  :  Shape  from  GeomAbs; 
             MaxDegree  :  Integer  ; 
             MaxSegments  :  Integer; 
    	     Only3d, 
    	     Only2d : Boolean  from  Standard  =  Standard_False)   
    returns  CurveOnSurface   from  Approx  
    raises ConstructionError; 


    IsDone(me) returns Boolean from Standard;
    
    HasResult(me) returns  Boolean from Standard;
   
    Curve3d(me) 
    returns  BSplineCurve  from  Geom; 
     
    MaxError3d(me) returns  Real; 
    
    Curve2d(me)   
   
    ---Purpose: 
    returns  BSplineCurve  from  Geom2d; 
     
    MaxError2dU(me)  returns  Real; 
    MaxError2dV(me) returns Real;
    
    ---Purpose : returns the maximum errors relativly to the  U component or the V component of the  
    --                 2d Curve
    
fields   

    myCurve2d    : BSplineCurve  from  Geom2d; 
    myCurve3d    : BSplineCurve  from  Geom; 
    myIsDone     : Boolean       from  Standard;   
    myHasResult  : Boolean       from  Standard;
    myError3d    : Real          from  Standard; 
    myError2dU   : Real          from  Standard; 
    myError2dV   : Real          from  Standard;  
     
end CurveOnSurface;
