-- Created on: 1991-07-24
-- Created by: Christophe MARION
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package BRepPrim 

	---Purpose: this package implements the primitives of the 
	--          Primitives package with the BRep Topology
	--          
	--          Contains :
	--          a Builder implementing the Template from Primitives
	--          
	--          The instantiations of the algorithms :
	--                OneAxis
	--                Wedge
	--                
	--          The rotational primitives inherited from OneAxis
	--          
	--                Revolution
	--                   Cylinder
	--                   Cone
	--                   Sphere
	--                   Torus
	--                   
	--          The  class FaceBuilder is  a tool to  build a face
	--          from a Geom surface.

uses
    gp,
    Geom2d,
    Geom,
    Primitives,
    TopoDS,
    BRep

is
    class Builder;

    deferred class OneAxis instantiates OneAxis from Primitives(
    	Shell   from TopoDS,
	Face    from TopoDS,
	Wire    from TopoDS,
	Edge    from TopoDS,
	Vertex  from TopoDS,
	Builder from BRepPrim);
	
    class Revolution;
    
    class Cylinder;
    
    class Cone;
    
    class Sphere;
    
    class Torus;
    
    class GWedge instantiates Wedge from Primitives(
    	Shell   from TopoDS,
	Face    from TopoDS,
	Wire    from TopoDS,
	Edge    from TopoDS,
	Vertex  from TopoDS,
	Builder from BRepPrim);
	
    class Wedge;
	
    class FaceBuilder;
    
end BRepPrim;
