-- Created on: 1994-11-14
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Pave from TopOpeBRepBuild 
    inherits Loop from TopOpeBRepBuild

uses
    
    ShapeEnum from TopAbs,
    Shape from TopoDS, 
    --modified by NIZHNY-MZV  Mon Feb 21 14:29:26 2000
    Kind  from  TopOpeBRepDS
is

    Create(V : Shape from TopoDS; P : Real; bound : Boolean) returns Pave;
    ---Purpose: V = vertex, P = parameter of vertex <V>
    --          bound = True if <V> is an old vertex
    --          bound = False if <V> is a new vertex
    
    HasSameDomain(me : mutable; b : Boolean);
    SameDomain(me : mutable; VSD : Shape from TopoDS);

    HasSameDomain(me) returns Boolean from Standard;
    SameDomain(me) returns Shape from TopoDS;
    ---C++: return const &

    Vertex(me) returns Shape from TopoDS is static;
    ---C++: return const &

    ChangeVertex(me : mutable) returns Shape from TopoDS is static;
    ---C++: return &
    -- used only by PaveSet
    Parameter(me) returns Real from Standard is static;
 
    --modified by NIZHNY-MZV  Mon Feb 21 14:09:47 2000 
    Parameter(me:  mutable;  Par:  Real  from  Standard)  is static;
    --modified by NIZHNY-MZV  Mon Feb 21 14:25:58 2000 
    InterferenceType(me:  mutable)  returns  Kind  from  TopOpeBRepDS; 
    ---C++: return &
	  
    IsShape(me) returns Boolean from Standard is redefined;
    Shape(me) returns Shape from TopoDS is redefined;
    ---C++: return const &

    Dump(me) is redefined;
    
fields

    myVertex  : Shape from TopoDS;
    myParam   : Real from Standard;
    myIsShape : Boolean from Standard;
    myHasSameDomain : Boolean from Standard;
    mySameDomain : Shape from TopoDS;

    --modified by NIZHNY-MZV  Mon Feb 21 14:26:58 2000 
    myIntType  :  Kind  from  TopOpeBRepDS; 

end Pave from TopOpeBRepBuild;
