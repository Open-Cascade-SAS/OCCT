-- Created on: 2001-04-24
-- Created by: Christian CAILLET
-- Copyright (c) 2001-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

--		ckyd@photox.paris1.matra-dtv.fr>

class ToleranceValue  from StepShape    inherits TShared

    ---Purpose : Added for Dimensional Tolerances

uses
    MeasureWithUnit from StepBasic

is

    Create returns mutable ToleranceValue;

    Init (me : mutable; lower_bound, upper_bound : MeasureWithUnit from StepBasic);

    LowerBound (me) returns MeasureWithUnit from StepBasic;
    SetLowerBound (me : mutable; lower_bound : MeasureWithUnit from StepBasic);

    UpperBound (me) returns MeasureWithUnit from StepBasic;
    SetUpperBound (me : mutable; upper_bound : MeasureWithUnit from StepBasic);

fields

    theLowerBound : MeasureWithUnit from StepBasic;
    theUpperBound : MeasureWithUnit from StepBasic;

end ToleranceValue;
