-- Created on: 1991-09-18
-- Created by: Didier PIFFAULT
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



generic class ToolPolyhedron from Intf (Polyhedron as any)

    ---Purpose: Describes the signature  of  a polyedral surface with  only
    --          triangular facets and the information  necessary to compute
    --          the interferences.


uses    XYZ from gp,
    	Pnt from gp,
    	Box from Bnd,
	HArray1OfBox from Bnd


raises  OutOfRange from Standard


is  Bounding       (myclass; thePolyh : Polyhedron)
    	    	    returns Box from Bnd;
    ---Purpose: Returns the bounding box of the ToolPolyhedron.

    ComponentsBounding
       	    	   (myclass; thePolyh : Polyhedron)
    	    	    returns HArray1OfBox from Bnd;
    ---Purpose: Returns the array of boxes. The box <n> corresponding 
    --          to the triangle <n>.


    DeflectionOverEstimation
		   (myclass; thePolyh : Polyhedron)
    	    	    returns Real from Standard;
    ---Purpose: Returns the tolerance of the polygon.


-- Structure needings :

    NbTriangles	   (myclass; thePolyh : Polyhedron) 
    	    	    returns Integer from Standard;
    ---Purpose: Returns the number of triangles in this polyedron.


    Triangle	   (myclass; thePolyh : Polyhedron;
		    Index     : in Integer from Standard;
		    P1,P2,P3  : out Integer from Standard)
		    raises OutOfRange from Standard;
    ---Purpose: Returns the indices  of  the 3 points of  the triangle of
    --          address Index in the ToolPolyhedron.


    Point	   (myclass; thePolyh : Polyhedron;
		    Index : in Integer)
		    returns Pnt from gp
		    raises OutOfRange from Standard;
    ---Purpose: Returns the point of index i in the polyedron.


    TriConnex	   (myclass; thePolyh : Polyhedron;
		    Triang	 : in Integer;
		    Pivot,Pedge	 : in Integer;
		    TriCon	 : out Integer;
		    OtherPedge	 : out Integer)
		    returns Integer
		    raises OutOfRange from Standard;
    ---Purpose: Returns  the  triangle <Tricon> connected  to  the triangle
    --          <Triang> by  the edge <Pivot><Pedge>.   The  third point of
    --          the connected triangle is returned in <OtherPedge> (Used to
    --          turn  around a vertex).   When the edge  <Pivot><Pedge>  is
    --          free  (no  connected triangle) <Tricon> is  null.   In this
    --          case the function returns the triangle on the free bound of
    --          the polyhedron connected to <Triang> by vertex <Pivot>.



end ToolPolyhedron;
