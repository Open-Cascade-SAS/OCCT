-- Created on: 1993-02-22
-- Created by: Philippe DAUTRY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class Vector from PGeom inherits Geometry from PGeom

        ---Purpose :  Defines a vector in 3D space.
        --  It can be a Direction (unitary vector) or a vector
        --  with magnitude.
        --  
	---See Also : Vector from Geom.

uses Vec from gp

is


    Initialize;
	---Purpose: Initializes the field(s) with default value(s).
    	---Level: Internal 


    Initialize(aVec: Vec from gp);
	---Purpose: Initializes the field vec with <aVec>.
    	---Level: Internal 


  Vec (me: mutable; aVec: Vec from gp);
        ---Purpose : Set the field vec.
    	---Level: Internal 


  Vec (me)  returns Vec from gp;
        ---Purpose : Returns the value of the field vec.
    	---Level: Internal 


fields

  vec : Vec from gp is protected;

end;
