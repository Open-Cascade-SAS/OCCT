-- Created on: 1997-07-28
-- Created by: Pierre CHALAMET
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

deferred class TextureMap from Graphic3d

inherits TextureRoot from Graphic3d

  ---Purpose: This is an abstract class for managing texture applyable on polygons.

uses 

  TypeOfTexture from Graphic3d,
  TextureParams from Graphic3d,
  LevelOfTextureAnisotropy from Graphic3d,
  AsciiString   from TCollection

is

  Initialize (theFileName : AsciiString from TCollection;
              theType     : TypeOfTexture from Graphic3d);

  EnableSmooth (me : mutable);
  ---Level: public
  ---Purpose:
  -- enable texture smoothing

  IsSmoothed (me) returns Boolean from Standard;
  ---Level: public
  ---Purpose:
  -- Returns TRUE if the texture is smoothed.

  DisableSmooth (me : mutable);
  ---Level: public
  ---Purpose:
  -- disable texture smoothing

  EnableModulate (me : mutable);
  ---Level: public
  ---Purpose:
  -- enable texture modulate mode.
  -- the image is modulate with the shading of the surface.

  DisableModulate (me : mutable);
  ---Level: public
  ---Purpose:
  -- disable texture modulate mode.
  -- the image is directly decal on the surface.

  IsModulate (me) returns Boolean from Standard;
  ---Level: public
  ---Purpose:
  -- Returns TRUE if the texture is modulate.

  EnableRepeat (me : mutable);
  ---Level: public
  ---Purpose:
  -- use this methods if you want to enable
  -- texture repetition on your objects.

  DisableRepeat (me : mutable);
  ---Level: public
  ---Purpose:
  -- use this methods if you want to disable
  -- texture repetition on your objects.

  IsRepeat (me) returns Boolean from Standard;
  ---Level: public
  ---Purpose:
  -- Returns TRUE if the texture repeat is enable.

  AnisoFilter (me) returns LevelOfTextureAnisotropy from Graphic3d;
  ---Level   : public
  ---Purpose : @return level of anisontropy texture filter.
  -- Default value is Graphic3d_LOTA_OFF.

  SetAnisoFilter (me : mutable;
                  theLevel : LevelOfTextureAnisotropy from Graphic3d);
  ---Level   : public
  ---Purpose : @param theLevel level of anisontropy texture filter.

end TextureMap from Graphic3d;
