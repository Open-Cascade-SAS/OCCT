-- Created on: 1997-09-11
-- Created by: Roman BORISOV
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ApproxCurve from GeomConvert 
    	---Purpose: A framework to convert a 3D curve to a 3D BSpline.
    	-- This is done by approximation to a BSpline curve within a given tolerance.
	
uses 
    Curve          from  Geom, 
    BSplineCurve   from  Geom, 
    Shape          from  GeomAbs,
    OutOfRange     from  Standard          
    
raises  OutOfRange   from Standard, 
        ConstructionError  from  Standard

is
 
    Create  (Curve:  Curve  from  Geom; 
    	    Tol3d:  Real; 
    	    Order:  Shape  from  GeomAbs; 
    	    MaxSegments:  Integer; 
    	    MaxDegree:  Integer)  returns  ApproxCurve; 
        ---Purpose: Constructs a curve approximation framework defined by -
    	--   -      the conic Curve, 
    	--   -      the tolerance value Tol3d, 
    	--   -      the degree of continuity Order, 
    	--   -      the maximum number of segments
    	--     MaxSegments allowed in the resulting BSpline curve, and 
    	--   -      the highest degree MaxDeg which the
    	--     polynomial defining the BSpline curve may have.
        
    Curve(me)  returns  BSplineCurve  from  Geom; 
    	--- Purpose: Returns the BSpline curve resulting from the approximation algorithm.
        
    IsDone(me)  returns  Boolean  from  Standard; 
    	---Purpose:  returns  Standard_True  if  the  approximation  has   
    	-- been  done  within  requiered tolerance 
     
    HasResult(me) returns Boolean; 
    	---Purpose: Returns  Standard_True if the approximation did come out 
    	-- with a result that  is not NECESSARELY within the required tolerance

    MaxError(me)  returns  Real  from  Standard; 
    	---Purpose:  Returns the greatest distance between a point on the
    	-- source conic and the BSpline curve resulting from the
    	-- approximation. (>0 when an approximation 
    	--  has  been  done, 0  if  no  approximation) 
     
    Dump(me;  o:  in  out  OStream); 
    	---Purpose:  Print on the stream  o  information about the object

fields
    myCurve     : Curve           from  Geom;
    myIsDone    : Boolean         from  Standard; 
    myHasResult : Boolean         from  Standard;     
    myBSplCurve : BSplineCurve    from  Geom; 
    myMaxError  : Real            from  Standard; 
    
end ApproxCurve;
