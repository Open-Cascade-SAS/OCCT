--
-- File:	AlienImage_AidaAlienImage.cdl
-- Created:	23/03/93
-- Author:	BBL
-- Modified:	02-06-98 : FMN ; Suppression appel Clear (deja fait dans ALienData)
--
---Copyright:	Matravision 1993
--

class AidaAlienImage from AlienImage inherits AlienUserImage from AlienImage

	---Version: 0.0

	---Purpose: This class defines an Aida Alien image ( BYTEMAPS ).
	---Keywords:
	---Warning:
	---References:

uses
	File 			from OSD,
	ColorMap 		from Aspect,
	Image			from Image,
	DitheringMethod 	from Image,
	AidaAlienData 		from AlienImage

is
	Create returns mutable AidaAlienImage from AlienImage;

	Clear( me : in out mutable) ;
	---Level: Public
	---Purpose: Frees memory allocated by AidaAlienImage

	ToImage( me : in immutable ) 
	  returns mutable Image from Image ;
	---Level: Public
	  ---Purpose : convert a AidaAlienImage object to a Image object.

	FromImage( me : in out mutable ; anImage : in Image from Image ) ;
	---Level: Public
	  ---Purpose : convert a Image object to a AidaAlienImage object.

	Read ( me : in out mutable; afile : in out File from OSD )
	  returns Boolean from Standard ;
	---Level: Public
	  ---Purpose: Read content of a AidaAlienImage object from a file .
	  --          Returns True if file is a Aida file .

	Write( me : in immutable; afile : in out File from OSD )
	  returns Boolean from Standard ;
	---Level: Public
	  ---Purpose: Write content of a  AidaAlienImage object to a file .

	SetColorImageDitheringMethod( me : in out mutable ; 
				      aMethod : DitheringMethod from Image;
				      aColorMap : ColorMap from Aspect ) ;

	---Level: Public
	  ---Purpose: Set the ImageDitheringMethod and the ColorMap when
	  --          FromImage is called with a ColorImage .
	  --	      Aida BYTEMAPS file handle only PseudoColorImage .
	  --          Default value is DM_NearestColor,
	  --		ColorCubeColorMap( 40, 5,1, 8,6, 3,54 )

fields
	myData : AidaAlienData  from  AlienImage;

end ;
 
