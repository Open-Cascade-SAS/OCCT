-- Created on: 1991-10-10
-- Created by: Jean Claude VAUTHIER
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class ConeToBSplineSurface  from Convert

        --- Purpose :
        --  This algorithm converts a bounded Cone into a rational 
        --  B-spline  surface.
        --  The cone a Cone from package gp. Its parametrization is :
        --  P (U, V) =  Loc + V * Zdir +
        --              (R + V*Tan(Ang)) * (Cos(U)*Xdir + Sin(U)*Ydir)
        --  where Loc is the location point of the cone, Xdir, Ydir and Zdir
        --  are the normalized directions of the local cartesian coordinate
        --  system of the cone (Zdir is the direction of the Cone's axis) ,
        --  Ang is the cone semi-angle.  The U parametrization range is
        --  [0, 2PI].
        --- KeyWords :
        --  Convert, Cone, BSplineSurface.

inherits ElementarySurfaceToBSplineSurface

uses Cone from gp

raises DomainError from Standard

is

  Create (C : Cone; U1, U2, V1, V2 : Real)  returns ConeToBSplineSurface
       --- Purpose : 
       --  The equivalent B-spline surface as the same orientation as the 
       --  Cone in the U and V parametric directions.
     raises DomainError;
        --- Purpose :
        --  Raised if U1 = U2 or U1 = U2 + 2.0 * Pi
        --  Raised if V1 = V2.


  Create (C : Cone; V1, V2 : Real)          returns ConeToBSplineSurface
       --- Purpose : 
       --  The equivalent B-spline surface as the same orientation as the
       --  Cone in the U and V parametric directions.
     raises DomainError;
        --- Purpose :
        --  Raised if V1 = V2.



end ConeToBSplineSurface;



