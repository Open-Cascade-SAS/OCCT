-- Created on: 1997-03-26
-- Created by: Christian CAILLET
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ItemDefinedTransformation  from StepRepr    inherits TShared

    ---Purpose : Added from StepRepr Rev2 to Rev4

uses
     HAsciiString from TCollection,
     RepresentationItem from StepRepr

is

    Create returns mutable ItemDefinedTransformation;

    Init (me : mutable;
    	  aName : HAsciiString from TCollection;
	  aDescription : HAsciiString from TCollection;
	  aTransformItem1 : RepresentationItem from StepRepr;
	  aTransformItem2 : RepresentationItem from StepRepr);

    SetName (me : mutable; aName : HAsciiString from TCollection);
    Name    (me) returns HAsciiString from TCollection;

    SetDescription (me : mutable; aDescription : HAsciiString from TCollection);
    Description    (me) returns HAsciiString from TCollection;

    SetTransformItem1 (me : mutable; aItem : RepresentationItem from StepRepr);
    TransformItem1    (me) returns RepresentationItem;

    SetTransformItem2 (me : mutable; aItem : RepresentationItem from StepRepr);
    TransformItem2    (me) returns RepresentationItem;

fields

    theName : HAsciiString from TCollection;
    theDescription : HAsciiString from TCollection;
    theTransformItem1 : RepresentationItem from StepRepr;
    theTransformItem2 : RepresentationItem from StepRepr;

end ItemDefinedTransformation;
