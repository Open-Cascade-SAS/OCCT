-- Created on: 2002-12-18
-- Created by: data exchange team
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SelectArrReal from StepData inherits SelectNamed from StepData

    ---Purpose :


uses

    AsciiString from TCollection,
    HArray1OfReal from TColStd

is

    Create returns SelectArrReal;

--    HasName (me) returns Boolean  is redefined;

--    Name (me) returns CString  is redefined;

--    SetName (me : mutable; name : CString)  returns Boolean  is redefined;
    -- redefined to accept any name

    Kind(me) returns Integer  is redefined;
    --  fixed kind : ArrReal

    ArrReal(me) returns HArray1OfReal from TColStd;

    SetArrReal(me:mutable; arr : HArray1OfReal from TColStd);

fields

    theArr  : HArray1OfReal from TColStd;

end SelectArrReal;
