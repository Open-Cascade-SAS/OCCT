-- File:        PresentationStyleAssignment.cdl
-- Created:     Mon Dec  4 12:02:29 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWPresentationStyleAssignment from RWStepVisual

	---Purpose : Read & Write Module for PresentationStyleAssignment

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     PresentationStyleAssignment from StepVisual,
     EntityIterator from Interface

is

	Create returns RWPresentationStyleAssignment;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable PresentationStyleAssignment from StepVisual);

	WriteStep (me; SW : in out StepWriter; ent : PresentationStyleAssignment from StepVisual);

	Share(me; ent : PresentationStyleAssignment from StepVisual; iter : in out EntityIterator);

end RWPresentationStyleAssignment;
