-- Created on: 1994-02-24
-- Created by: Laurent BOURESCHE
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class CurveTool from BRepLProp

uses Vec   from gp,
     Pnt   from gp,
     Dir   from gp,
     Curve from BRepAdaptor

is

    Value(myclass; C : Curve from BRepAdaptor; U : Real; P : out Pnt);
    ---Purpose: Computes the point <P> of parameter <U> on the curve <C>.
     	
    D1   (myclass; C : Curve from BRepAdaptor; 
          U : Real; P : out Pnt; V1 : out Vec);
    ---Purpose: Computes the point <P> and first derivative <V1> of 
    --          parameter <U> on the curve <C>.

    D2   (myclass; C : Curve from BRepAdaptor; 
          U : Real; P : out Pnt; V1, V2 : out Vec);
    ---Purpose: Computes the point <P>, the first derivative <V1> and second
    --          derivative <V2> of parameter <U> on the curve <C>.
    
    D3   (myclass; C : Curve from BRepAdaptor; 
          U : Real; P : out Pnt; V1, V2, V3 : out Vec);
    ---Purpose: Computes the point <P>, the first derivative <V1>, the 
    --          second derivative <V2> and third derivative <V3> of 
    --          parameter <U> on the curve <C>.

     Continuity(myclass; C : Curve from BRepAdaptor) returns Integer;
     ---Purpose: returns the order of continuity of the curve <C>.
     --          returns 1 : first derivative only is computable
     --          returns 2 : first and second derivative only are computable.
     --          returns 3 : first, second and third are computable.

     FirstParameter(myclass; C : Curve from BRepAdaptor) returns Real;
     ---Purpose: returns the first parameter bound of the curve.
     --          
     
     LastParameter(myclass; C : Curve from BRepAdaptor) returns Real;
     ---Purpose: returns the last parameter bound of the curve.
     --          FirstParameter must be less than LastParamenter.

end CurveTool;


