-- File:	LoopPointTool.cdl
-- Created:	Mon Mar  9 16:55:09 1992
-- Author:	Isabelle GRIGNON
--		<isg@phobox>
---Copyright:	 Matra Datavision 1992

deferred generic class LoopPointTool from IntWalk 
    (LoopPoint as any)

	---Purpose: template class to describe the necessary ressources 
	--          for a point usedas a starting point for a marching 
	--          algorithm.
	--          The 'marching algorithm' determines the intersection 
	--          between an implicit surface and a parametrized surface.
	--          these point are inside the surface not on the boundaries.

uses Pnt from gp,
     Vec from gp,
     Dir2d from gp

is

    Value3d(myclass; PStart: LoopPoint)
    
      	---Purpose: Returns the 3d coordinates of the starting point.

    	returns Pnt from gp;


    Value2d(myclass; PStart: LoopPoint; U, V: out Real from Standard);
    
	---Purpose: Returns the <U,V> parameters which are associated 
	--          with <P>
	--          it's the parameters which start the marching algorithm


    Direction3d(myclass; PStart: LoopPoint)
    
        ---Purpose: returns the tangent at the intersectin in 3d space
        --          associated to <P>

    	returns Vec from gp;


    Direction2d(myclass; PStart: LoopPoint)
    
        ---Purpose: returns the tangent at the intersectin in the
        --          parametric space of the parametrized surface.This tangent
        --          is associated to the value2d

    	returns Dir2d from gp;


end LoopPointTool;
