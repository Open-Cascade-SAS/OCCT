-- Created on: 1993-03-09
-- Created by: Philippe DAUTRY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package TColGeom 

        ---Purpose : This package  is used to  instantiate of  several
        --         generic classes from  the package  TCollection with
        --         objects from the package Geom.

uses TCollection, Geom

is



    imported Array1OfCurve;
    imported Array1OfBezierCurve;
    imported Array1OfBSplineCurve;
    imported Array1OfSurface;

    imported transient class HArray1OfCurve;
    imported transient class HArray1OfBezierCurve;
    imported transient class HArray1OfBSplineCurve;
    imported transient class HArray1OfSurface;

    imported Array2OfSurface;
    imported Array2OfBezierSurface;

    imported transient class HArray2OfSurface;

    imported SequenceOfCurve;
    imported SequenceOfBoundedCurve;
    imported SequenceOfSurface;

    imported transient class HSequenceOfCurve;
    imported transient class HSequenceOfBoundedCurve;

end TColGeom;
