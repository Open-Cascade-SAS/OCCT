-- Created on: 1994-05-19
-- Created by: Yves FRICAUD
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


package Bisector 

    --- Purpose : This package provides the bisecting line between two
    --            geometric elements.

uses 
     MMgt,
     Standard,
     TCollection,
     TColStd,	
     TColgp,
     Geom2d,
     GeomAbs,
     gp,
     math,
     IntCurve,	
     GccInt,
     StdFail,
     IntRes2d
is

    deferred class Curve;
    
   	     class BisecAna;
    	     --- Purpose: This class provides the bisecting line between two
    	     --           geometric elements.The elements are Circles,Lines or
    	     --           Points. 

    	     class BisecPC;
	     ---Purpose: This class provides the bisecting line between a point
	     --          a Curve.
    
    	     class BisecCC;	
	     ---Purpose: This class provides the bisecting line between two
	     --          Curves. 

    class Bisec;
	---Purpose: This class provides the bisecting line between two
	--          geometris  elelements.  The   bisecting   line  is
	--          trimmed by a point, 
    
    class Inter;
    
    class PointOnBis;
    
    class PolyBis;
    
    private class FunctionH;
    
    private class FunctionInter;
    
    IsConvex (Cu : Curve from Geom2d; Sign : Real) 
    returns Boolean from Standard;
    
end Bisector;
