-- Created on: 1999-08-11
-- Created by: Roman LYGIN
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class TransferResultInfo from TransferBRep inherits TShared from MMgt 

    ---Purpose: Data structure for storing information on transfer result.
    --          At the moment it dispatches information for the following types:
    --          - result,
    --          - result + warning(s),
    --          - result + fail(s),
    --          - result + warning(s) + fail(s)
    --          - no result,
    --          - no result + warning(s),
    --          - no result + fail(s),
    --          - no result + warning(s) + fail(s),

is

    Create returns TransferResultInfo from TransferBRep;
    	---Purpose: Creates object with all fields nullified.
	
    Clear (me: mutable);
    	---Purpose: Resets all the fields.
	
    Result (me: mutable) returns Integer;
    	---C++: inline
    	---C++: return &
	
    ResultWarning (me: mutable) returns Integer;
    	---C++: inline
    	---C++: return &
	
    ResultFail (me: mutable) returns Integer;
    	---C++: inline
    	---C++: return &
	
    ResultWarningFail (me: mutable) returns Integer;
    	---C++: inline
    	---C++: return &
	
    NoResult (me: mutable) returns Integer;
    	---C++: inline
    	---C++: return &
	
    NoResultWarning (me: mutable) returns Integer;
    	---C++: inline
    	---C++: return &
	
    NoResultFail (me: mutable) returns Integer;
    	---C++: inline
    	---C++: return &
	
    NoResultWarningFail (me: mutable) returns Integer;
    	---C++: inline
    	---C++: return &
	
fields

    myR,  myRW,  myRF,  myRWF,
    myNR, myNRW, myNRF, myNRWF: Integer;
    
end TransferResultInfo;
