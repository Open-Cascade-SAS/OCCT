-- File:	Approx_Curve3d.cdl
-- Created:	Thu Aug 20 18:31:06 1998
-- Author:	Philippe MANGIN
--		<pmn@sgi29>
---Copyright:	 Matra Datavision 1998

class  Curve3d  from  Approx 

uses
    HCurve         from  Adaptor3d, 
    BSplineCurve   from  Geom, 
    Shape          from  GeomAbs,
    OutOfRange     from  Standard          
    
raises  OutOfRange   from Standard, 
        ConstructionError  from  Standard

is
 
    Create(Curve:  HCurve  from Adaptor3d; 
    	    Tol3d:  Real; 
    	    Order:  Shape  from  GeomAbs; 
    	    MaxSegments:  Integer; 
    	    MaxDegree:  Integer)  returns  Curve3d  from  Approx; 
        ---Purpose: Approximation  of  a  curve  with respect of the  
    --          requiered tolerance Tol3D. 
     
    Curve(me)  returns  BSplineCurve  from  Geom; 
     
    IsDone(me)  returns  Boolean  from  Standard; 
    ---Purpose:  returns  Standard_True  if  the  approximation  has   
    -- been  done  within  requiered tolerance 
     
    HasResult(me) returns Boolean; 
    ---Purpose: returns  Standard_True if the approximation did come out 
    -- with a result that  is not NECESSARELY within the required 
    -- tolerance

    MaxError(me)  returns  Real  from  Standard; 
    ---Purpose:  returns  the  Maximum  Error  (>0 when an approximation 
    --  has  been  done, 0  if  no  approximation) 
     
    Dump(me;  o:  in  out  OStream); 
    ---Purpose:  Print on the stream  o  information about the object

fields
    myIsDone    : Boolean         from  Standard; 
    myHasResult : Boolean         from  Standard;     
    myBSplCurve : BSplineCurve    from  Geom; 
    myMaxError  : Real            from  Standard; 
    
end Curve3d;
