-- Created on: 1993-01-13
-- Created by: CKY / Contract Toubro-Larsen ( Deepak PRABHU )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class GeneralLabel from IGESDimen  inherits IGESEntity

        ---Purpose: defines GeneralLabel, Type <210> Form <0>
        --          in package IGESDimen
        --          Used for general labeling with leaders

uses

        GeneralNote          from IGESDimen,
        LeaderArrow          from IGESDimen,
        HArray1OfLeaderArrow from IGESDimen

raises OutOfRange

is

        Create returns GeneralLabel;

        -- Specific Methods pertaining to the class

        Init (me          : mutable;
              aNote       : GeneralNote;
              someLeaders : HArray1OfLeaderArrow);
        ---Purpose : This method is used to set the fields of the class
        --           GeneralLabel
        --       - aNote       : General Note Entity
        --       - someLeaders : Associated Leader Entities

        Note (me) returns GeneralNote;
        ---Purpose : returns General Note Entity

        NbLeaders (me) returns Integer;
        ---Purpose : returns Number of Leaders

        Leader (me; Index : Integer) returns LeaderArrow
        raises OutOfRange;
        ---Purpose : returns Leader Entity
        -- raises exception if Index <= 0 or Index > NbLeaders()

fields

--
-- Class    : IGESDimen_GeneralLabel
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class GeneralLabel.
--
-- Reminder : A GeneralLabel instance is defined by :
--            - Note    : General Note Entity
--            - Leaders : Associated Leader Entities
-- An GeneralLabel Entity consists of a general note with one or more
-- associated leaders.

        theNote      : GeneralNote;
        theLeaders   : HArray1OfLeaderArrow;

end GeneralLabel;
