-- Created on: 1993-02-05
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package Contap

    ---Purpose: 

uses Standard,StdFail,MMgt, GeomAbs, TopAbs, TCollection, gp, TColgp,
     math, IntSurf, IntStart, IntWalk,
     Geom2d, TColStd, Geom, Adaptor3d,  Adaptor2d


is


    class Point;

    class Line;

    class SurfFunction;

    class ArcFunction;

    class SurfProps;

    class Contour;

    class TheSequenceOfPoint instantiates Sequence from TCollection (Point from Contap);

    class TheHSequenceOfPoint instantiates HSequence from TCollection
        (Point              from Contap,
         TheSequenceOfPoint from Contap);

    class TheSequenceOfLine instantiates Sequence from TCollection(Line from Contap);

    class TheSearch instantiates SearchOnBoundaries from IntStart
        (HVertex      from Adaptor3d,
         HCurve2d     from Adaptor2d,
         HCurve2dTool from Contap,
         HContTool    from Contap,
         TopolTool    from Adaptor3d,
         ArcFunction  from Contap);

    class TheIWalking instantiates IWalking from IntWalk
        (PathPoint               from IntSurf,
         PathPointTool           from IntSurf,
         SequenceOfPathPoint     from IntSurf,
         InteriorPoint           from IntSurf,
         InteriorPointTool       from IntSurf,
         SequenceOfInteriorPoint from IntSurf,
         HSurface                from Adaptor3d,
         HSurfaceTool            from Adaptor3d,
         SurfFunction            from Contap);

    class TheSearchInside instantiates SearchInside from IntStart
        (HSurface     from Adaptor3d,
         HSurfaceTool from Adaptor3d,
         TopolTool    from Adaptor3d,
         HContTool    from Contap,
         SurfFunction from Contap);

         
    class ContAna;

    enumeration TFunction is
        ContourStd,
        ContourPrs,
        DraftStd,
        DraftPrs
    end TFunction;

    enumeration IType is  -- a replacer dans IntSurf et fusionner avec IntPatch
    -- type of the line of contour
        Lin,       -- pour conflit avec deferred class Line
        Circle,
        Walking,
        Restriction
    end IType;

    class HContTool;
    
    class HCurve2dTool;

end Contap;
