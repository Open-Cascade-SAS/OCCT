-- Created on: 1997-02-21
-- Created by: Alexander BRIVIN
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ShadedShape from VrmlConverter  

   	---Purpose:  ShadedShape - computes  the  shading presentation of shapes
    	--           by triangulation algorithms, converts this one into VRML objects 
        --           and writes (adds) into anOStream.
        --           All requested properties of the representation including 
    	--           the maximal chordial deviation  are specify in aDrawer.  
        --           This  kind  of  the  presentation  is  converted  into
        --           IndexedFaceSet ( VRML ).

uses 
 
    Drawer       from  VrmlConverter, 
    Shape        from  TopoDS, 
    Face         from  TopoDS,
    Connect      from  Poly, 
    Array1OfDir  from  TColgp

is      
     
    Add(myclass; anOStream  : in out OStream from  Standard;
    	    	 aShape     :        Shape   from  TopoDS;
                 aDrawer    :        Drawer  from  VrmlConverter);

        
    ComputeNormal(myclass; aFace  :        Face        from TopoDS;
    	    	           pc     : in out Connect     from Poly;
		           Nor    : out    Array1OfDir from TColgp);

    
end ShadedShape  from  VrmlConverter;
