-- Created on: 1992-12-02
-- Created by: Isabelle GRIGNON
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SelGProps from GProp inherits GProps

    	    ---Purpose: 
    	    --          Computes the global properties of an elementary 
    	    --          surface (surface of the gp package)

uses  Cylinder from gp,
      Cone     from gp,
      Pnt      from gp,
      Sphere   from gp,
      Torus    from gp

is

  Create returns SelGProps;

  Create (S : Cylinder; Alpha1, Alpha2, Z1, Z2 : Real; SLocation : Pnt)   
     returns SelGProps;


  Create (S : Cone; Alpha1, Alpha2, Z1, Z2 : Real; SLocation : Pnt)   
     returns SelGProps;


  Create (S : Sphere from gp; Teta1, Teta2, Alpha1, Alpha2 : Real;
          SLocation : Pnt)   
     returns SelGProps;


  Create (S : Torus from gp; Teta1, Teta2, Alpha1, Alpha2 : Real;
          SLocation : Pnt)   
     returns SelGProps;

  SetLocation(me : in out ;SLocation :Pnt);

  Perform(me : in out;S : Cylinder; Alpha1, Alpha2, Z1, Z2 : Real);

  Perform(me : in out;S : Cone; Alpha1, Alpha2, Z1, Z2 : Real);

  Perform(me : in out;S : Sphere; Teta1, Teta2, Alpha1, Alpha2 : Real);

  Perform(me : in out;S : Torus; Teta1, Teta2, Alpha1, Alpha2 : Real);

end SelGProps;
