-- Created on: 2002-12-12
-- Created by: data exchange team
-- Copyright (c) 2002-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class RepresentedDefinition from StepRepr
inherits SelectType from StepData

    ---Purpose: Representation of STEP SELECT type RepresentedDefinition

uses
    GeneralProperty from StepBasic,
    PropertyDefinition from StepRepr,
    PropertyDefinitionRelationship from StepRepr,
    ShapeAspect from StepRepr,
    ShapeAspectRelationship from StepRepr

is
    Create returns RepresentedDefinition from StepRepr;
	---Purpose: Empty constructor

    CaseNum (me; ent: Transient) returns Integer;
	---Purpose: Recognizes a kind of RepresentedDefinition select type
	--          1 -> GeneralProperty from StepBasic
	--          2 -> PropertyDefinition from StepRepr
	--          3 -> PropertyDefinitionRelationship from StepRepr
	--          4 -> ShapeAspect from StepRepr
	--          5 -> ShapeAspectRelationship from StepRepr
	--          0 else

    GeneralProperty (me) returns GeneralProperty from StepBasic;
	---Purpose: Returns Value as GeneralProperty (or Null if another type)

    PropertyDefinition (me) returns PropertyDefinition from StepRepr;
	---Purpose: Returns Value as PropertyDefinition (or Null if another type)

    PropertyDefinitionRelationship (me) returns PropertyDefinitionRelationship from StepRepr;
	---Purpose: Returns Value as PropertyDefinitionRelationship (or Null if another type)

    ShapeAspect (me) returns ShapeAspect from StepRepr;
	---Purpose: Returns Value as ShapeAspect (or Null if another type)

    ShapeAspectRelationship (me) returns ShapeAspectRelationship from StepRepr;
	---Purpose: Returns Value as ShapeAspectRelationship (or Null if another type)

end RepresentedDefinition;
