-- File:        DocumentType.cdl
-- Created:     Mon Dec  4 12:02:29 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWDocumentType from RWStepBasic

	---Purpose : Read & Write Module for DocumentType

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     DocumentType from StepBasic,
     EntityIterator from Interface

is

	Create returns RWDocumentType;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable DocumentType from StepBasic);

	WriteStep (me; SW : in out StepWriter; ent : DocumentType from StepBasic);

	Share(me; ent : DocumentType from StepBasic; iter : in out EntityIterator);

end RWDocumentType;
