-- Created on: 1993-07-27
-- Created by: Jean Louis FRENKEL
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




deferred class Image from Image inherits TShared from MMgt

	---Purpose: This class defined the general behavior of an Image from
	--		Package Image .

uses

    PlaneAngle 		from Quantity,
    FlipType		from Image,
    Color 		from Quantity,
    Array1OfColor 	from Quantity,
    HArray1OfColor 	from Quantity,
    Pixel		from Aspect,
    PixelAddress 	from Image,
    TypeOfImage 	from Image,
    Type                from Standard
is
    Initialize( aPixelType : Type from Standard );
	---Level: Public
	---Purpose: Image constructor ,initialise the Image PixelType.

    Destroy( me : mutable )
	is virtual ;
	---C++: alias ~
	---Level: Public
	---Purpose: Image destructor.

    isSamePixel( me : immutable ; 
	X,Y    	     		: in Integer from Standard ;
	anotherImage 		: immutable like me ;
	anotherX,anotherY	: in Integer from Standard ) 
	returns Boolean from Standard is deferred ;
	---Level: Public
	---Purpose: Returns True if me->Pixel(X,Y) is equal to 
	--	    anotherImage->Pixel(anotherX,anotherY)

    PixelColor( me : immutable ; X,Y : in Integer from Standard )
    	returns Color from Quantity is deferred ;
	---C++: return const &
   	---Purpose: Returns the Color of an Image Pixel.

    RowColor  ( me : immutable ; Y : in Integer from Standard )
	returns HArray1OfColor from Quantity is virtual ;
	---Purpose: Returns the Color of an Image Pixel Row.

    RowColor  ( me       : immutable ; 
		Y        : in Integer from Standard ;
		aArray1  : in out Array1OfColor from Quantity )
	is virtual ;
	---Purpose: Stores the Color of an Image Pixel Row in aArray1.

    PixelType( me : immutable ) returns Type from Standard ;
	---Level: Public
	---Purpose: Returns the Image Pixel Type.

    Size    ( me : immutable )  returns Integer from Standard ;
	---Purpose: Returns the Image size in Pixel unit ( width*height) .

    InternalDup( me : mutable ; anImage : immutable like me ) 
	is deferred ;
	---Purpose : Duplicates an Image.

    -- ******************* Deferred method of Image ******************* 

    SetOrigin( me : mutable ; x,y : in Integer from Standard ) 
		is deferred ;
	---Purpose: Sets Image origin, for Rotation, copy between image ...
	--		Image origin is on the TOP LEFT . Y axis goes TOP to
	--		DOWN , X axis goes LEFT to RIGHT.

    LowerX  ( me : immutable )  returns Integer from Standard is deferred ;
	---Level: Public
	---Purpose: Returns the lower X Image coordinate ( X Origin ).

    UpperX  ( me : immutable )  returns Integer from Standard is deferred ;
	---Level: Public
	---Purpose: Returns the upper X Image coordinate 
	--		( X Origin + Image width - 1 ).

    Width   ( me : immutable )  returns Integer from Standard is deferred ;
	---Level: Public
	---Purpose: Returns the Image width.

    LowerY  ( me : immutable )  returns Integer from Standard is deferred ;
	---Level: Public
	---Purpose: Returns the lower Y Image coordinate ( Y Origin ).

    UpperY  ( me : immutable )  returns Integer from Standard is deferred ;
	---Level: Public
	---Purpose: Returns the upper Y Image coordinate 
	--		( Y Origin + Image height - 1 ).

    Height  ( me : immutable )  returns Integer from Standard is deferred ;
	---Level: Public
	---Purpose: Returns the Image height.
 
    Resize( me : mutable ;
	XOffset,XScale, YOffset,YScale : Real from Standard ) is deferred ;
	---Level: Public
	---Purpose: Resize an Image. Image Pixel are left unchanged at there
	--	      absolute positon. Resulting Image can be clipped.
	--	newLowerX = LowerX()*XScale + XOffset
	--	newLowerY = LowerY()*YScale + YOffset
	--	newUpperX = UpperX()*XScale + XOffset
	--	newUpperY = UpperY()*YScale + YOffset
	--	newWidth  = Width() *XScale
	--	newHeight = Height()*YScale

    Type    ( me : immutable )  returns TypeOfImage from Image is deferred ;
	---Level: Public
	---Purpose: Returns the ImageType TOI_ColorImage or TOI_PseudoColorImage

    Pixel   ( me : immutable ; 	X,Y    : in Integer from Standard ;
				aPixel : in out Pixel from Aspect ) 
	is deferred ;
	---Level: Public
	---Purpose: Get the Image Pixel Value at X,Y coordinate in aPixel.
	-- Warning: aPixel must have the same type than Image Pixel.

    SetPixel( me : mutable ; 	X,Y    : in Integer from Standard ;
				aPixel : in Pixel   from Aspect ) 
	is deferred ;
	---Level: Public
	---Purpose: Store aPixel in the Image  at X,Y coordinate .
	-- Warning: aPixel must have the same type than Image Pixel.

    Pixel   ( me : immutable ; 	X,Y    : in Integer from Standard ;
				aPixel : in out PixelAddress from Image ) 
	is deferred ;
	---Level: Public
	---Purpose: Get the Image Pixel Value at X,Y coordinate in aPixel.
	-- Warning: aPixel must have the same type than Image Pixel.

    SetPixel( me : mutable ; 	X,Y    : in Integer from Standard ;
				aPixel : in PixelAddress from Image ) 
	is deferred ;
	---Level: Public
	---Purpose: Store aPixel in the Image  at X,Y coordinate .
	-- Warning: aPixel must have the same type than Image Pixel.

    Transpose ( me : mutable ; aType : in FlipType from Image ) is deferred ;
	---Level: Public
	---Purpose: Transpose an Image( flipping across horizontal axis or 
	--		vertical axis, or across diagonal... )
	--	    This geometric transformation preserves all Image Pixels.
	--	    We don't need to interpolate pixels .
	--	    Warning : Image size change during Transpose.

    Clip      ( me : mutable ; X,Y,Width,Height:in Integer from Standard)
								is deferred ;
	---Level: Public
	---Purpose: Extract a SubImage starting at coordinate X,Y 
	--		to (X+Width-1),(Y+Height-1).
	--	    Warning : the Image size and origin change, new origin
	--	    is X,Y ; new size is Width,Height.

    Shift     ( me : mutable ; XShift,YShift  :in Integer from Standard)
								is deferred ;
	---Level: Public
	---Purpose: Translate an Image XShift pixel Right, YShift Down .
	--	    Shift parameter are Integer value.

    Fill      ( me : mutable ; SrcImage : immutable like me ) is deferred ;
	---Level: Public
	---Purpose: Fill me with SrcImage. SrcImage pixel are copied starting
	--	     at SrcImage->LowerX(),SrcImage->LowerY() in MyPixelField.
	--	     SrcImage Pixel are clipped outside <me>.

    Fill      ( me : mutable ; SrcImage : immutable like me ;
		SrcX, SrcY, SrcWidth, SrcHeight,
		X, Y : in Integer from Standard ) is deferred ;
	---Level: Public
	---Purpose: Fill me with a SubImage of SrcImage starting from 
	--	    SrcX, SrcY to (SrcX+SrcWidth-1),(SrcY+SrcHeight-1) in 
	--	    Src Image coordinate. SrcImage SubImage pixels are copied 
	--	    starting at X,Y in MyPixelField.
	--	    SrcImage Pixel are clipped outside <me>.

    Clear     ( me : mutable ) is deferred ;
	---Level: Public
	---Purpose: Fill the entire Image with the BackgroundPixel.

    Dup      ( me : immutable ) returns mutable Image from Image is deferred;
	---Level: Public
	---Purpose : Duplicate an Image.

    Dump( me : immutable ) is deferred ;
	---Level: Public
	---Purpose: Debug

fields
	myPixelType : Type from Standard ;

end Image from Image;
