-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Protocol from StepAP214 inherits Protocol from StepData
	---Purpose : Protocol for StepAP214 Entities
	--           It requires StepAP214 as a Resource

uses Protocol from Interface,
     CString from Standard

is
	Create returns mutable Protocol from StepAP214;
	TypeNumber (me; atype : any Type) returns Integer is redefined;
	---Purpose :Returns a Case Number for each of the StepAP214 Entities
	SchemaName(me) returns CString from Standard is redefined;
	-- was C++ : return const

    NbResources (me) returns Integer  is redefined;
    ---Purpose : Returns count of Protocol used as Resources (level one)

    Resource (me; num : Integer) returns Protocol from Interface  is redefined;
    ---Purpose : Returns a Resource, given its rank (between 1 and NbResources)

end Protocol;
