-- File:        DefinitionalRepresentation.cdl
-- Created:     Mon Dec  4 12:02:25 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWDefinitionalRepresentation from RWStepRepr

	---Purpose : Read & Write Module for DefinitionalRepresentation

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     DefinitionalRepresentation from StepRepr,
     EntityIterator from Interface

is

	Create returns RWDefinitionalRepresentation;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable DefinitionalRepresentation from StepRepr);

	WriteStep (me; SW : in out StepWriter; ent : DefinitionalRepresentation from StepRepr);

	Share(me; ent : DefinitionalRepresentation from StepRepr; iter : in out EntityIterator);

end RWDefinitionalRepresentation;
