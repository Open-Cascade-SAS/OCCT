-- Created on: 2018-03-15
-- Created by: Stephan GARNAUD (ARM)
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.








class Environment from OSD

   ---Purpose: Management of system environment variables
   --          An environment variable is composed of a variable name
   --          and its value.
   --
   --          To be portable among various systems, environment variables
   --          are local to a process.

uses Protection, Error, AsciiString from TCollection
raises ConstructionError, NullObject, OSDError

is
 Create returns Environment;
   ---Purpose: Creates the object Environment.
   ---Level: Public

 Create (Name : AsciiString) returns Environment
   ---Purpose: Creates an Environment variable initialized with value
   --          set to an empty AsciiString.
   ---Level: Public
   raises ConstructionError;

 Create (Name, Value : AsciiString) returns Environment
   ---Purpose: Creates an Environment variable initialized with Value.
   raises ConstructionError, NullObject;
   -- ConstructionError is raised when invalid character is encountered.
   ---Level: Public

 SetValue (me : in out; Value : AsciiString)
   ---Purpose: Changes environment variable value.
   --          Raises ConstructionError either if the string contains 
   --          characters not in range of ' '...'~' or if the string 
   --          contains the character '$' which is forbiden.
   ---Level: Public
   raises ConstructionError  is static;

 Value (me : in out) returns AsciiString is static ;
   ---Purpose: Gets the value of an environment variable
   ---Level: Public

 SetName (me : in out; name : AsciiString)
   ---Purpose: Changes environment variable name.
   --          Raises ConstructionError either if the string contains 
   --          characters not in range of ' '...'~' or if the string 
   --          contains the character '$' which is forbiden.
   ---Level: Public
   raises ConstructionError  is static;

 Name (me ) returns AsciiString  is static;
   ---Purpose: Gets the name of <me>.
   ---Level: Public

 Build (me : in out) is static ;
   ---Purpose: Sets the value of an environment variable
   --          into system (physically).
   ---Level: Public

 Remove(me : in out) is static ;
   ---Purpose: Removes (physically) an environment variable 
   ---Level: Public

 Failed (me) returns Boolean is static ;
   ---Purpose: Returns TRUE if an error occurs
   ---Level: Public

 Reset (me : in out) is static ;
   ---Purpose: Resets error counter to zero
   ---Level: Public
      
 Perror (me : in out)
   ---Purpose: Raises OSD_Error
   ---Level: Public
   raises OSDError is static ;

 Error (me) returns Integer is static ;
   ---Purpose: Returns error number if 'Failed' is TRUE.
   ---Level: Publi

fields
   myName  : AsciiString;  --- Name of the variable
   myValue : AsciiString;
   myError : Error;
end Environment from OSD;



