-- Created on: 1997-02-18
-- Created by: Stagiaire Francois DUMONT
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



package Hermit 

	---Purpose: This  is used to  reparameterize Rational  BSpline
	--           Curves so that we can   concatenate them later to
	--          build C1 Curves  It builds and 1D-reparameterizing
	--          function starting from an Hermite interpolation and
	--          adding knots and modifying poles of the 1D BSpline
	--          obtained that way. The goal is to build a(u) so that
	--          if we consider a BSpline curve 
	--                          N(u)
	--                 f(u) =  -----
        --                          D(u)
        --                          
        --          the function a(u)D(u) has value 1 at the umin and umax
        --          and has 0.0e0 derivative value a umin and umax.
        --          The details of the computation occuring in this package
        --          can be found by reading :
        --          " Etude sur la concatenation de NURBS en vue du 
        --            balayage de surfaces" PFE n S85 Ensam Lille
uses
    Geom,
    Geom2d,
    TColStd,
    TColgp
    
is			   					
            
    Solution( BS     :  BSplineCurve from Geom;
    	      TolPoles : in Real from Standard=0.000001;
	      TolKnots : in Real from Standard=0.000001)
      ---Purpose:returns the correct spline a(u) which will
      --                 be multiplicated with BS later.
    returns BSplineCurve from Geom2d;
    	    	
    Solution( BS     :  BSplineCurve from Geom2d;
    	      TolPoles : in Real from Standard=0.000001;
	      TolKnots : in Real from Standard=0.000001)
      ---Purpose:returns the correct spline a(u) which will
      --                 be multiplicated with BS later.
    returns BSplineCurve from Geom2d;
    
    Solutionbis( BS       :  BSplineCurve from Geom;
    	    	 Knotmin  : out Real from Standard;
		 Knotmax  : out Real from Standard;
    	         TolPoles : in Real from Standard=0.000001;
	         TolKnots : in Real from Standard=0.000001);
      ---Purpose:returns the knots to insert to a(u) to 
      --         stay with a constant sign and in the 
      --         tolerances. 
    
end Hermit;


