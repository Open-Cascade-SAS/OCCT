-- Created on: 1998-05-20
-- Created by: Christian CAILLET
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class SignText  from MoniTool    inherits TShared
 
        ---Purpose : Provides the basic service to get a text which identifies
        --           an object in a context
        --           It can be used for other classes (general signatures ...)
        --           It can also be used to build a message in which an object
        --           is to be identified
 
uses CString, Transient, AsciiString from TCollection
 
is
 
    Name (me) returns CString  is deferred;
    ---Purpose : Returns an identification of the Signature (a word), given at
    --           initialization time

    TextAlone (me; ent : any Transient)
    	returns AsciiString from TCollection  is virtual;
    ---Purpose : Gives a text as a signature for a transient object alone, i.e.
    --           without defined context.
    --           By default, calls Text with undefined context (Null Handle) and
    --           if empty, then returns DynamicType

    Text (me; ent : any Transient; context : any Transient)
    	returns AsciiString from TCollection  is deferred;
    ---Purpose : Gives a text as a signature for a transient object in a context
    --           If the context is senseless, it can be given as Null Handle
    --           empty result if nothing to give (at least the DynamicType could
    --           be sent ?)

end SignText;
