-- Created on: 1995-05-10
-- Created by: Denis PASCAL 
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- modified     Sergey Zaritchny



package PDataXtd 

	---Purpose: 


uses Standard,
     PDF,
     PTopoDS,
     PGeom,
     PNaming, 
     PDataStd,
     PCollection,
     PColStd,
     PTopLoc,
     PGeom, 
     TColStd,
     gp

is


    ---Purpose: General Data
    --          ============ 

    class Position;
    
    class Point;
    
    class Axis;
    
    class Plane;  

    class Geometry;  -- Point | Line ...etc..
    
    class Constraint;
    
    class Placement;
    
    class PatternStd;
    
    class Shape; 
     
 
end PDataXtd;
