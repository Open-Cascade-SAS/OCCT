-- Created on: 1993-04-30
-- Created by: Yves FRICAUD
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class BasicElt from MAT 

	---Purpose: A    BasicELt  is  associated   to  each  elemtary
	--          constituant of  the figure.

inherits 

    TShared from MMgt

uses
    Arc            from MAT,
    Side           from MAT,
    Address        from Standard
is
    
    Create (anInteger : Integer) 
    	--- Purpose : Constructor, <anInteger> is the <index> of <me>.
    returns mutable BasicElt from MAT;

    StartArc(me)  
    	--- Purpose : Return <startArcLeft> or <startArcRight> corresponding
    	--            to <aSide>.
    returns Arc is static;

    EndArc(me)  
    	--- Purpose : Return <endArcLeft> or <endArcRight> corresponding
    	--            to <aSide>.
    returns Arc is static;
     
    Index (me) 
    	--- Purpose : Return the <index> of <me> in Graph.TheBasicElts.
    returns Integer is static;

    GeomIndex(me) 
    	--- Purpose : Return the <GeomIndex> of <me>.
    returns Integer is static;
    
    SetStartArc (me : mutable ; anArc : Arc)
    is static;
    
    SetEndArc (me : mutable ; anArc : Arc)
    is static;
    
    SetIndex (me : mutable ; anInteger : Integer)
    is static;

    SetGeomIndex(me : mutable ; anInteger : Integer)
    is static;
    
fields
    startLeftArc  : Address from Standard;
    endLeftArc    : Address from Standard;
    index         : Integer;
    geomIndex     : Integer;
    
end BasicElt;






