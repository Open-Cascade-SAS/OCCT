-- Created on: 1997-05-14
-- Created by: Robert COUBLANC
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SensitiveTriangle from Select3D  
inherits SensitivePoly from Select3D

    ---Purpose: A framework to define selection of triangles in a view.
    -- This comes into play in the detection of meshing and triangulation in surfaces.
    -- In some cases this class can raise Standard_ConstructionError and 
    -- Standard_OutOfRange exceptions. For more details see Select3D_SensitivePoly.

uses
    EntityOwner      from SelectBasics,
    Projector        from Select3D,
    Lin              from gp,
    ListOfBox2d      from SelectBasics,
    PickArgs         from SelectBasics,
    Array1OfPnt2d    from TColgp,
    Box2d            from Bnd,
    XY               from gp,
    Pnt              from gp,
    TypeOfSensitivity from Select3D,
    Location          from TopLoc, 
    SensitiveEntity   from Select3D

raises
    ConstructionError from Standard,
    OutOfRange from Standard

is
    Create (OwnerId      : EntityOwner from SelectBasics;
            P1,P2,P3     : Pnt from gp;
            Sensitivity  : TypeOfSensitivity = Select3D_TOS_INTERIOR)
     returns SensitiveTriangle;
    ---Level: Public 
        ---Purpose: Constructs a sensitive triangle object defined by the
        -- owner OwnerId, the points P1, P2, P3, and the type of sensitivity Sensitivity. 

    Matches (me : mutable;
             thePickArgs : PickArgs from SelectBasics;
             theMatchDMin, theMatchDepth : out Real from Standard)
    returns Boolean is redefined static;
    ---Level: Public
    ---Purpose: Checks whether the sensitive entity matches the picking
    -- detection area (close to the picking line).
    -- For details please refer to base class declaration.

    Matches (me  :mutable; 
             XMin,YMin,XMax,YMax : Real from Standard;
             aTol: Real from Standard) 
    returns Boolean
    is redefined virtual;
        ---Level: Public 
     
    Matches (me  :mutable; 
             Polyline:Array1OfPnt2d from TColgp;
         aBox:Box2d from Bnd;
             aTol: Real from Standard) 
    returns Boolean
    is redefined virtual;
        ---Level: Public 
    
    
    ComputeDepth(me;EyeLine: Lin from gp) 
    returns Real from Standard;


    Points3D(me; P1,P2,P3 : out Pnt from gp) ;
        ---Purpose: Returns the 3D points P1, P2, P3 used at the time of construction.
    Center3D (me) returns Pnt from gp;
        ---Purpose: Returns the center point of the sensitive triangle created at construction time.
    Center2D (me) returns XY from gp;
        ---Purpose: WARNING : the returned Values are the original values
        --          without the stored  location (if there's one).
        --          To get the genuine value, One must apply this location
        --          (Method Location() )
    
    
    
    
    Status(me; 
             X,Y  : Real from Standard;
             aTol : Real from Standard ;
             Dmin : out Real from Standard)
    returns Integer from Standard;
    
    Status (myclass;
             p0,p1,p2: XY from gp ;
             aPoint  : XY from gp ;
             aTol    : Real from Standard;
             Dmin    : out Real from Standard) returns Integer from  Standard;
    ---Purpose: Dmin gives the distance between the cdg and aPoint return 

    Dump(me; S: in out OStream;FullDump : Boolean from Standard = Standard_True) is redefined virtual; 

    GetConnected(me: mutable; theLocation : Location from TopLoc) 
    returns SensitiveEntity from Select3D 
    is redefined virtual; 
        ---Level: Public 
        ---Purpose: Returns the copy of this


fields
    mytype  : TypeOfSensitivity from Select3D;
end SensitiveTriangle;
