-- Created on: 1991-07-23
-- Created by: Christophe MARION
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




package Primitives 

	---Purpose: This  package   describes   algorithms  to   build
	--          topological primitives.
	--          
	--          The algorithms  in  this package  are  generic. It
	--          contains :
	--          
	--           *   The Builder  signature   class. Describes the
	--           services    required  from    the  Topology  Data
	--           Structure to build the following primitives.
	--          
	--           * The  OneAxis generic class.  Algorithm  used to
	--           build rotational primitives.
	--               
	--           *  The  Wedge  generic  class. Algorithm to build
	--           boxes and wedges.

uses
    gp        -- gp provides all geometrical information

is


    enumeration Direction is 
	---Purpose: 
    	XMin, XMax, YMin, YMax, ZMin, ZMax
    end Direction;


    deferred generic class Builder;
    
    deferred generic class OneAxis;
    	
    generic class Wedge; 
    
end Primitives;
