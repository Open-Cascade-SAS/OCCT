-- File:	RWStepRepr_RWPropertyDefinition.cdl
-- Created:	Mon Jul  3 16:29:03 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class RWPropertyDefinition from RWStepRepr

    ---Purpose: Read & Write tool for PropertyDefinition

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    PropertyDefinition from StepRepr

is
    Create returns RWPropertyDefinition from RWStepRepr;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : PropertyDefinition from StepRepr);
	---Purpose: Reads PropertyDefinition

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: PropertyDefinition from StepRepr);
	---Purpose: Writes PropertyDefinition

    Share (me; ent : PropertyDefinition from StepRepr;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWPropertyDefinition;
