-- Created on: 1993-01-09
-- Created by: CKY / Contract Toubro-Larsen ( TCD )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class IntercharacterSpacing from IGESGraph  inherits IGESEntity

        ---Purpose: defines IGESIntercharacterSpacing, Type <406> Form <18>
        --          in package IGESGraph
        --
        --          Specifies the gap between letters when fixed-pitch
        --          spacing is used

uses  Integer, Real  -- no one specific type


is

        Create returns mutable IntercharacterSpacing;

        -- Specific Methods pertaining to the class

        Init (me       : mutable;
              nbProps  : Integer;
              anISpace : Real);
        ---Purpose : This method is used to set the fields of the class
        --           IntercharacterSpacing
        --       - nbProps  : Number of property values (NP = 1)
        --       - anISpace : Intercharacter spacing percentage

        NbPropertyValues (me) returns Integer;
        ---Purpose : returns the number of property values in <me>

        ISpace (me) returns Real;
        ---Purpose : returns the Intercharacter Space of <me> in percentage
        -- of the text height (Range = 0..100)

fields

--
-- Class    : IGESGraph_IntercharacterSpacing
--
-- Purpose  : Declaration of the variables specific to a
--            Intercharacter Spacing property.
--
-- Reminder : An Intercharacter spacing property is defined by :
--                  - Number of property values (NP=1)
--                  - ISpace
--

        theNbPropertyValues : Integer;

        theISpace           : Real;

end IntercharacterSpacing;
