-- File:	TPrsStd_PlaneDriver.cdl
-- Created:	Fri Aug  1 11:21:30 1997
-- Author:	SMO
---Copyright:	 Matra Datavision 1997


class PlaneDriver from TPrsStd inherits Driver from TPrsStd
---Purpose: An implementation of TPrsStd_Driver for planes.
uses

  GUID               from Standard,
  Label              from TDF,
  InteractiveObject  from AIS
is

    Create
    returns mutable PlaneDriver from TPrsStd;
---Purpose: Constructs an empty plane driver.
    Update (me : mutable ;
           aLabel      : Label from TDF;
	   anAISObject : in out InteractiveObject from AIS)
    returns Boolean from Standard
    is  redefined virtual;
    --- Purpose: Build the AISObject (if null) or update it.
    --           No compute is done.
    --           Returns <True> if informations was found
    --           and AISObject updated. 
	   

end PlaneDriver;

