-- Created on: 2001-12-13
-- Created by: Sergey KUUl
-- Copyright (c) 2001-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class TimerSentry from MoniTool

    ---Purpose: A tool to facilitate using MoniTool_Timer functionality
    --          by automatically ensuring consistency of start/stop actions
    --
    --          When instance of TimerSentry is created, a timer 
    --          with corresponding name is started
    --          When instance is deleted, timer stops

uses
    Timer from MoniTool
    
is

    Create (cname: CString from Standard) 
    returns TimerSentry from MoniTool;
        ---C++: inline
        ---Purpose: Constructor creates an instance and runs the corresponding timer
    
    Create (timer: Timer from MoniTool) 
    returns TimerSentry from MoniTool;
        ---C++: inline
        ---Purpose: Constructor creates an instance and runs the corresponding timer
    
    Destroy(me: in out);
        ---C++: inline
    	---Purpose: Destructor stops the associated timer
        ---C++: alias "Standard_EXPORT ~MoniTool_TimerSentry () { Destroy(); }"

    Timer (me) returns Timer from MoniTool;
        ---C++: inline

    Stop (me: in out);
        ---C++: inline
    	---Purpose: Manually stops the timer

fields

    myTimer: Timer from MoniTool;

end TimerSentry;
