-- Created on: 1997-02-12
-- Created by: Alexander BRIVIN
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class WWWInline from Vrml 

	---Purpose: defines a WWWInline node of VRML specifying group properties.
    	--  The  WWWInline  group  node  reads  its  children  from  anywhere  in  the   
    	--  World  Wide  Web.
	--  Exactly  when  its  children  are  read  is  not  defined; 
	--  reading  the  children  may  be  delayed  until  the  WWWInline  is  actually 
    	--  displayed. 
	--  WWWInline  with  an  empty  ("")  name  does  nothing. 
	--  WWWInline  behaves  like  a  Separator,  pushing  the  traversal  state 
	--  before  traversing  its  children  and  popping  it  afterwards.
    	--  By  defaults: 
	--    myName  ("")
	--    myBboxSize (0,0,0)
	--    myBboxCenter  (0,0,0)

uses
 
    AsciiString   from   TCollection,
    Vec           from   gp 

is
 
    Create returns  WWWInline from Vrml; 

    Create  ( aName        :   AsciiString from  TCollection; 
    	      aBboxSize    :   Vec         from  gp;
    	      aBboxCenter  :   Vec         from  gp )
    	returns  WWWInline from Vrml; 

    SetName ( me : in out; aName : AsciiString from TCollection );
    Name ( me )  returns  AsciiString from TCollection;

    SetBboxSize ( me : in out; aBboxSize  : Vec  from  gp);
    BboxSize ( me )  returns   Vec  from  gp;

    SetBboxCenter ( me : in out; aBboxCenter  : Vec  from  gp);
    BboxCenter ( me )  returns  Vec  from  gp;

    Print  ( me;  anOStream: in out OStream from Standard) returns OStream from Standard;
    ---C++:  return  & 

fields
 
    myName        :   AsciiString from TCollection;   -- URL name
    myBboxSize    :   Vec         from gp;            -- Size of 3D bounding box
    myBboxCenter  :   Vec         from gp;            -- Center of 3D bounding box
    
end WWWInline;

