-- File:	RWStepFEA_RWFeaGroup.cdl
-- Created:	Thu Dec 12 17:51:05 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWFeaGroup from RWStepFEA

    ---Purpose: Read & Write tool for FeaGroup

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    FeaGroup from StepFEA

is
    Create returns RWFeaGroup from RWStepFEA;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : FeaGroup from StepFEA);
	---Purpose: Reads FeaGroup

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: FeaGroup from StepFEA);
	---Purpose: Writes FeaGroup

    Share (me; ent : FeaGroup from StepFEA;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWFeaGroup;
