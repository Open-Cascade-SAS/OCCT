-- Created on: 2002-02-20
-- Created by: Andrey BETENEV
-- Copyright (c) 2002-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class ProgressScale from Message 

    ---Purpose: Internal data structure for scale in ProgressIndicator
    --
    --          Basically it defines three things:
    --          - name that can be used for generating user messages
    --          - limits and characteristics of the current scale,
    --            along with derived coefficients to map it into basic scale [0-1]
    --          - methods for conversion of values from current scale
    --            to basic one and back
    --
    --          NOTE: There is no special protection against bad input data
    --          like min > max etc. except cases when it can cause exception

uses
    HAsciiString from TCollection
is

    Create returns ProgressScale from Message;
    	---Purpose: Creates scale ranged from 0 to 100 with step 1

    ---Scope: Access to fields

    SetName(me : out; theName : CString);
    	---C++:inline
    SetName(me : out; theName : HAsciiString from TCollection);
    	---C++:inline
    	---Purpose: Sets scale name
    
    GetName(me) returns HAsciiString from TCollection;
    	---C++:inline
    	---Purpose: Gets scale name
	--          Name may be Null handle if not set

    SetMin(me : out; theMin : Real);
    	---C++:inline
    	---Purpose: Sets minimum value of scale
    
    GetMin(me) returns Real;
    	---C++:inline
    	---Purpose: Gets minimum value of scale

    SetMax(me : out; theMax : Real);
    	---C++:inline
    	---Purpose: Sets minimum value of scale
    
    GetMax(me) returns Real;
    	---C++:inline
    	---Purpose: Gets minimum value of scale

    SetRange (me: out; min, max: Real);
    	---C++: inline
    	---Purpose: Set both min and max
	
    SetStep(me : out; theStep : Real);
    	---C++:inline
    	---Purpose: Sets default step
    
    GetStep(me) returns Real;
    	---C++:inline
    	---Purpose: Gets default step

    SetInfinite(me : out; theInfinite : Boolean = Standard_True);
    	---C++:inline
    	---Purpose: Sets flag for infinite scale
    
    GetInfinite(me) returns Boolean;
    	---C++:inline
    	---Purpose: Gets flag for infinite scale

    SetScale (me: out; min, max, step: Real; theInfinite : Boolean = Standard_True);
    	---C++: inline
    	---Purpose: Set all scale parameters
	
    ---Scope: Mapping to base scale
    
    SetSpan (me: out; first, last: Real);
    	---C++: inline
    	---Purpose: Defines span occupied by the scale on the basis scale
	
    GetFirst (me) returns Real;
    	---C++: inline
    GetLast (me) returns Real;
    	---C++: inline
    	---Purpose: Return information on span occupied by the scale on the base scale
	
    LocalToBase (me; val: Real) returns Real;
    BaseToLocal (me; val: Real) returns Real;
    	---Purpose: Convert value from this scale to base one and back

fields
    
    myName: HAsciiString from TCollection; -- name
    
    myMin, myMax: Real;     -- range of a scale
    myStep : Real;          -- default step
    myInfinite: Boolean;    -- flag for infinite scale

    myFirst, myLast : Real; -- span on base scale

end ProgressScale;
