-- File:	StepFEA_FeaShellMembraneStiffness.cdl
-- Created:	Thu Dec 12 17:51:06 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class FeaShellMembraneStiffness from StepFEA
inherits FeaMaterialPropertyRepresentationItem from StepFEA

    ---Purpose: Representation of STEP entity FeaShellMembraneStiffness

uses
    HAsciiString from TCollection,
    SymmetricTensor42d from StepFEA

is
    Create returns FeaShellMembraneStiffness from StepFEA;
	---Purpose: Empty constructor

    Init (me: mutable; aRepresentationItem_Name: HAsciiString from TCollection;
                       aFeaConstants: SymmetricTensor42d from StepFEA);
	---Purpose: Initialize all fields (own and inherited)

    FeaConstants (me) returns SymmetricTensor42d from StepFEA;
	---Purpose: Returns field FeaConstants
    SetFeaConstants (me: mutable; FeaConstants: SymmetricTensor42d from StepFEA);
	---Purpose: Set field FeaConstants

fields
    theFeaConstants: SymmetricTensor42d from StepFEA;

end FeaShellMembraneStiffness;
