-- Created by: Peter KURNEV
-- Copyright (c) 2010-2014 OPEN CASCADE SAS
-- Copyright (c) 2007-2010 CEA/DEN, EDF R&D, OPEN CASCADE
-- Copyright (c) 2003-2007 OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN, CEDRAT,
--                         EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class FaceInfo from BOPDS 

	---Purpose: 
    	-- The class BOPDS_FaceInfo is to store  
    	-- handy information about state of face
uses     
    BaseAllocator from BOPCol,
    MapOfInteger from BOPCol,
    IndexedMapOfPaveBlock from BOPDS
   
--raises

is
    Create 
    	returns FaceInfo from BOPDS; 
    ---C++: inline 	 
    ---C++: alias "virtual ~BOPDS_FaceInfo();"  
      	---Purpose:  
    	--- Empty contructor  
    	---   
	 
    Create (theAllocator: BaseAllocator from BOPCol) 
    	returns FaceInfo from BOPDS;  
    ---C++: inline   
    	---Purpose:   
     	---  Contructor    
    	---  theAllocator - the allocator to manage the memory     
    	---    
	
    Clear(me:out); 
    	---Purpose:   
     	---  Clears the contents      
    
    SetIndex(me:out; 
    	    theI: Integer from Standard); 
    ---C++: inline 
     	---Purpose: 
    	--- Modifier   
	--- Sets the index of the face <theI> 
	
    Index(me) 
    	returns Integer from Standard; 
    ---C++: inline  
    	---Purpose: 
    	--- Selector   
	--- Returns the index of the face 
    --  
    -- In 
    --  
    PaveBlocksIn(me) 
	returns IndexedMapOfPaveBlock from BOPDS; 
    ---C++: return const &  
    ---C++: inline 
     	---Purpose: 
    	--- Selector   
	--- Returns the pave blocks of the face 
	--- that  have state In 
	 
    ChangePaveBlocksIn(me:out) 
    	returns IndexedMapOfPaveBlock from BOPDS;  
    ---C++: return &  
    ---C++: inline    
      	---Purpose: 
    	--- Selector/Modifier   
	--- Returns the pave blocks  
    	--  of the face 
	--- that  have state In 
	 
    VerticesIn(me) 
    	returns MapOfInteger from BOPCol;  
    ---C++: return const &  
    ---C++: inline  
     	---Purpose: 
    	--- Selector   
	--- Returns the list of indices for vertices  
    	--  of the face
	--- that have state In  
	
    ChangeVerticesIn(me:out) 
    	returns MapOfInteger from BOPCol;  
    ---C++: return &  
    ---C++: inline 
    	---Purpose: 
    	--- Selector/Modifier    
	--- Returns the list of indices for vertices  
    	--  of the face
	--- that have state In   
    --  
    -- On 
    --  
    PaveBlocksOn(me) 
	returns IndexedMapOfPaveBlock from BOPDS; 
    ---C++: return const &  
    ---C++: inline    
    	---Purpose: 
    	--- Selector   
	--- Returns the pave blocks of the face 
	--- that  have state On
     
    ChangePaveBlocksOn(me:out) 
    	returns IndexedMapOfPaveBlock from BOPDS;  
    ---C++: return &  
    ---C++: inline    
      	---Purpose: 
    	--- Selector/Modifier   
	--- Returns the pave blocks  
    	--  of the face 
	--- that  have state On 
    VerticesOn(me) 
    	returns MapOfInteger from BOPCol;  
    ---C++: return const &  
    ---C++: inline  
     	---Purpose: 
    	--- Selector   
	--- Returns the list of indices for vertices  
    	--  of the face
	--- that have state On 
	 
    ChangeVerticesOn(me:out) 
    	returns MapOfInteger from BOPCol;  
    ---C++: return &  
    ---C++: inline 
    	---Purpose: 
    	--- Selector/Modifier   
	--- Returns the list of indices for vertices  
    	--  of the face
	--- that have state On   
    --  
    -- Sections 
    --  
    PaveBlocksSc(me) 
	returns IndexedMapOfPaveBlock from BOPDS; 
    ---C++: return const &  
    ---C++: inline   
    	---Purpose: 
    	--- Selector   
	--- Returns the pave blocks of the face 
	--- that are  pave blocks of section edges  
     
    ChangePaveBlocksSc(me:out) 
    	returns IndexedMapOfPaveBlock from BOPDS;  
    ---C++: return &  
    ---C++: inline  
    	--- Selector/Modifier      
	--- Returns the pave blocks of the face 
	--- that are  pave blocks of section edges     
      
    VerticesSc(me) 
    	returns MapOfInteger from BOPCol;  
    ---C++: return const &  
    ---C++: inline  
    	---Purpose: 
    	--- Selector   
	--- Returns the list of indices for section  vertices  
    	--  of the face
     
    ChangeVerticesSc(me:out) 
    	returns MapOfInteger from BOPCol;  
    ---C++: return &  
    ---C++: inline 
    	---Purpose: 
    	--- Selector/Modifier   
	--- Returns the list of indices for section  vertices  
    	--  of the face 
    --  
    -- Others
    --    
    --Update(me:out) 
    --	is protected; 
     
fields 
    myAllocator   : BaseAllocator from BOPCol is protected; 
    myIndex       : Integer from Standard is protected; 
    myPaveBlocksIn: IndexedMapOfPaveBlock from BOPDS is protected;  
    myVerticesIn  : MapOfInteger from BOPCol is protected;  
    myPaveBlocksOn: IndexedMapOfPaveBlock from BOPDS is protected;  
    myVerticesOn  : MapOfInteger from BOPCol is protected;
    myPaveBlocksSc: IndexedMapOfPaveBlock from BOPDS is protected;  
    myVerticesSc  : MapOfInteger from BOPCol is protected;
 
end FaceInfo;
