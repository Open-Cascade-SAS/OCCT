-- Created on: 1996-10-21
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


package TestTopOpe

uses 
 
    Draw,
    TopOpeBRepBuild,
    TopOpeBRepDS,
    TopoDS
    
is

    AllCommands(I : in out Interpretor from Draw);
    ---Purpose: Defines all Top. Ope. test commands

    TOPOCommands(I : in out Interpretor from Draw);

    BOOPCommands(I : in out Interpretor from Draw);

    HDSCommands(I : in out Interpretor from Draw);
    ---Purpose: commands on a HDS involved in topological operations

    CurrentHB(HDS : HBuilder from TopOpeBRepBuild);
    ---Purpose : Defines the HBuilder on which BOOPCommands will operate.

    CurrentDS(HDS : HDataStructure from TopOpeBRepDS);
    ---Purpose : Defines the HDS on which HDSCommands/BOOPCommands will operate.

    Shapes(S1,S2 : Shape from TopoDS);
    ---Purpose: Defines current shapes of current topological operation

    MesureCommands(I : in out Interpretor from Draw);

    CORCommands(I : in out Interpretor from Draw);

    DSACommands(I : in out Interpretor from Draw);

    OtherCommands(I : in out Interpretor from Draw);

    Factory (theDI : out Interpretor from Draw);
    ---Purpose: Loads all Draw commands of TKDrawDEB. Used for plugin.

end TestTopOpe;
