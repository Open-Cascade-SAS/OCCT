-- Created on: 1993-01-26
-- Created by: Jean-Louis FRENKEL
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class ToolRFace from StdPrs 

	---Purpose: 
uses 
    Curve        from Geom2dAdaptor,
    Face         from TopoDS,
    HSurface     from BRepAdaptor,
    Curve2dPtr   from Adaptor2d,
    Orientation  from TopAbs,
    Explorer     from TopExp

is
    Create returns ToolRFace from StdPrs;    

    Create ( aSurface :HSurface from BRepAdaptor ) 
    returns ToolRFace from StdPrs;

    IsOriented (me) returns Boolean from Standard;

    Init(me: in out); 


    More(me) returns Boolean from Standard;

    Next(me: in out);

    Value(me) returns Curve2dPtr from Adaptor2d;

    Orientation(me) returns Orientation from TopAbs;    

fields
    myFace      : Face       from TopoDS;
    myExplorer  : Explorer   from TopExp;
    DummyCurve  : Curve      from Geom2dAdaptor;
    
end ToolRFace;


