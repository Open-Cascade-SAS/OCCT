-- Created on: 2002-12-12
-- Created by: data exchange team
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class PropertyDefinitionRepresentation from StepRepr
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity PropertyDefinitionRepresentation

uses
    RepresentedDefinition from StepRepr,
    Representation from StepRepr

is
    Create returns PropertyDefinitionRepresentation from StepRepr;
	---Purpose: Empty constructor

    Init (me: mutable; aDefinition: RepresentedDefinition from StepRepr;
                       aUsedRepresentation: Representation from StepRepr);
	---Purpose: Initialize all fields (own and inherited)

    Definition (me) returns RepresentedDefinition from StepRepr;
	---Purpose: Returns field Definition
    SetDefinition (me: mutable; Definition: RepresentedDefinition from StepRepr);
	---Purpose: Set field Definition

    UsedRepresentation (me) returns Representation from StepRepr;
	---Purpose: Returns field UsedRepresentation
    SetUsedRepresentation (me: mutable; UsedRepresentation: Representation from StepRepr);
	---Purpose: Set field UsedRepresentation

fields
    theDefinition: RepresentedDefinition from StepRepr;
    theUsedRepresentation: Representation from StepRepr;

end PropertyDefinitionRepresentation;
