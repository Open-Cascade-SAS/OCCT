-- File:	BRepTools_GTrsfModification.cdl
-- Created:	Mon Dec 30 15:58:53 1996
-- Author:	Stagiaire Mary FABIEN
--		<fbi@zozox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1996

class GTrsfModification from BRepTools inherits Modification from BRepTools

	---Purpose: Defines a modification of the  geometry by a  GTrsf
	--          from gp. All methods return True and transform the
	--          geometry.

uses Face     from TopoDS,
     Edge     from TopoDS,
     Vertex   from TopoDS,
     Location from TopLoc,
     Shape    from GeomAbs,
     
     Surface  from Geom,
     Curve    from Geom,
     Curve    from Geom2d,
     
     GTrsf     from gp,
     Pnt      from gp

is

    Create (T : GTrsf from gp) returns mutable GTrsfModification from BRepTools; 
    
    GTrsf(me: mutable)
	---Purpose: Gives an access on the GTrsf.
	---C++: return &
    	returns GTrsf from gp
	is static;


    NewSurface(me: mutable; F       :     Face     from TopoDS;
                            S       : out Surface  from Geom;
		            L       : out Location from TopLoc;
		            Tol     : out Real     from Standard;
                            RevWires : out Boolean from Standard;
                            RevFace  : out Boolean from Standard)
    
      	---Purpose: Returns Standard_True  if  the face  <F> has  been
      	--          modified.  In this  case, <S> is the new geometric
      	--          support of  the  face, <L> the  new location,<Tol>
      	--          the new  tolerance.<RevWires> has  to  be set   to
      	--          Standard_True   when the modification reverses the
      	--          normal of  the   surface.(the wires   have  to  be
      	--          reversed).   <RevFace>   has   to   be   set    to
      	--          Standard_True if  the orientation  of the modified
      	--          face changes in the  shells which contain  it.  --
      	--          Here, <RevFace>  will  return Standard_True if the
      	--          -- gp_Trsf is negative. 
    
    
    	returns Boolean from Standard
	;
	

    NewCurve(me: mutable; E  :     Edge     from TopoDS;
                          C  : out Curve    from Geom;
		          L  : out Location from TopLoc;
		          Tol: out Real     from Standard)
    
    	returns Boolean from Standard
	;
	
	---Purpose: Returns Standard_True  if  the edge  <E> has  been
	--          modified.  In this case,  <C> is the new geometric
	--          support of the  edge, <L> the  new location, <Tol>
	--          the         new    tolerance.   Otherwise, returns
	--          Standard_False,    and  <C>,  <L>,   <Tol> are not
	--          significant.
    

    NewPoint(me: mutable; V  :     Vertex   from TopoDS;
                          P  : out Pnt      from gp;
		          Tol: out Real     from Standard)
    
    	returns Boolean from Standard
	;
	
	---Purpose: Returns  Standard_True if the  vertex <V> has been
	--          modified.  In this  case, <P> is the new geometric
	--          support of the vertex,   <Tol> the new  tolerance.
	--          Otherwise, returns Standard_False, and <P>,  <Tol>
	--          are not significant.
    

    NewCurve2d(me: mutable;  E    :     Edge     from TopoDS;
                             F    :     Face     from TopoDS;
                             NewE :     Edge     from TopoDS;
                             NewF :     Face     from TopoDS;
                             C    : out Curve    from Geom2d;
		             Tol  : out Real     from Standard)
    
    	returns Boolean from Standard
	;
	
	---Purpose: Returns Standard_True if  the edge  <E> has a  new
	--          curve on surface on the face <F>.In this case, <C>
	--          is the new geometric support of  the edge, <L> the
	--          new location, <Tol> the new tolerance.
	--          Otherwise, returns  Standard_False, and <C>,  <L>,
	--          <Tol> are not significant.
    

    NewParameter(me: mutable; V  :     Vertex   from TopoDS;
                              E  :     Edge     from TopoDS;
                              P  : out Real     from Standard;
  		              Tol: out Real     from Standard)
    
    	returns Boolean from Standard
	;
	
	---Purpose: Returns Standard_True if the Vertex  <V> has a new
	--          parameter on the  edge <E>. In  this case,  <P> is
	--          the parameter,    <Tol>  the     new    tolerance.
	--          Otherwise, returns Standard_False, and <P>,  <Tol>
	--          are not significant.
    


    

    Continuity(me: mutable; E          : Edge from TopoDS;
    	                    F1,F2      : Face from TopoDS;
			    NewE       : Edge from TopoDS;
			    NewF1,NewF2: Face from TopoDS)
    
    	returns Shape from GeomAbs
	
	---Purpose: Returns the  continuity of  <NewE> between <NewF1>
	--          and <NewF2>.
	--          
	--          <NewE> is the new  edge created from <E>.  <NewF1>
	--          (resp. <NewF2>) is the new  face created from <F1>
	--          (resp. <F2>).

    	;



fields

    myGTrsf : GTrsf from gp;
    myGScale: Real;

end GTrsfModification;
