-- Created on: 1993-03-26
-- Created by: Christian CAILLET
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DefaultGeneral  from StepData    inherits GeneralModule  from StepData

    ---Purpose : DefaultGeneral defines a GeneralModule which processes
    --           Unknown Entity from StepData  only

uses OStream, Transient ,
     EntityIterator , CopyTool, Check, ShareTool

is

    Create returns DefaultGeneral;
    ---Purpose : Creates a Default General Module

    	--  Reconduction because limitation cdl  --

    FillSharedCase (me; casenum : Integer; ent : Transient;
    	iter : in out EntityIterator);
    ---Purpose : Specific filling of the list of Entities shared by an Entity
    --           <ent>, which is an UnknownEntity from StepData.

    CheckCase (me; casenum : Integer; ent : Transient; shares : ShareTool;
    	       ach : in out Check);
    ---Purpose : Specific Checking of an Entity <ent>

    NewVoid (me; CN : Integer; entto : out Transient)
    	returns Boolean;
    ---Purpose : Specific creation of a new void entity

    CopyCase (me; casenum : Integer;
    	      entfrom : Transient; entto : Transient;
    	      TC : in out CopyTool);
    ---Purpose : Specific Copy ("Deep") from <entfrom> to <entto> (same type)
    --           by using a CopyTool which provides its working Map.
    --           Use method Transferred from TransferControl to work


end DefaultGeneral;
