-- Created on: 1991-10-04
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.





class BSplineSurfaceKnotSplitting   from GeomConvert

        --- Purpose : An algorithm to determine isoparametric curves along
    	-- which a BSpline surface should be split in order to
    	-- obtain patches of the same continuity.
        --  For a B-spline surface the discontinuities are localised at
        --  the knot values. Between two knots values the B-spline is
        --  infinitely continuously differentiable.  For each parametric 
        --  direction at a knot of range index the continuity in this
        --  direction is equal to :  Degree - Mult (Index)   where  Degree
        --  is the degree of the basis B-spline functions and Mult the
        --  multiplicity of the knot of range Index in the given direction.
        --  If for your computation you need to have B-spline surface with a 
        --  minima of continuity it can be interesting to know between which
        --  knot values, a B-spline patch, has a continuity of given order.
        --  This algorithm computes the indexes of the knots where you should
        --  split the surface, to obtain patches with a constant continuity
        --  given at the construction time. If you just want to compute the
        --  local derivatives on the surface you don't need to create the
        --  BSpline patches, you can use the functions LocalD1, LocalD2, 
        --  LocalD3, LocalDN of the class BSplineSurface from package Geom.




uses  BSplineSurface       from Geom,
      Array1OfInteger      from TColStd,
      HArray1OfInteger      from TColStd

raises  DimensionError  from Standard,
        RangeError      from Standard
  
is


  Create (BasisSurface : BSplineSurface; 
          UContinuityRange, VContinuityRange : Integer)
     returns BSplineSurfaceKnotSplitting;
    	--- Purpose : Determines the u- and v-isoparametric curves
    	--  along which the BSpline surface BasisSurface
    	-- should be split in order to obtain patches with a
    	-- degree of continuity equal to UContinuityRange in
    	-- the u parametric direction, and to
    	-- VContinuityRange in the v parametric direction.
    	-- These isoparametric curves are defined by
    	-- parameters, which are BasisSurface knot values in
    	-- the u or v parametric direction. They are identified
    	-- by indices in the BasisSurface knots table in the
    	-- corresponding parametric direction.
    	-- Use the available interrogation functions to access
    	-- computed values, followed by the global function
    	-- SplitBSplineSurface (provided by the package
    	-- GeomConvert) to split the surface.
    	-- Exceptions
    	-- Standard_RangeError if UContinuityRange or
    	-- VContinuityRange is less than zero.

  NbUSplits (me)   returns Integer  is static;
        --- Purpose : Returns the number of u-isoparametric curves
    	-- along which the analysed BSpline surface should be
    	-- split in order to obtain patches with the continuity
    	-- required by this framework.
    	-- The parameters which define these curves are knot
    	-- values in the corresponding parametric direction.
    	-- Note that the four curves which bound the surface are
    	-- counted among these splitting curves.
        
  NbVSplits (me)  returns Integer   is static;
       	--- Purpose : Returns the number of v-isoparametric curves
    	-- along which the analysed BSpline surface should be
    	-- split in order to obtain patches with the continuity
    	-- required by this framework.
    	-- The parameters which define these curves are knot
    	-- values in the corresponding parametric direction.
    	-- Note that the four curves which bound the surface are
    	-- counted among these splitting curves.


  Splitting (me; USplit, VSplit : in out Array1OfInteger)
        --- Purpose: Loads the USplit and VSplit tables with the split
    	-- knots values computed in this framework. Each value
    	-- in these tables is an index in the knots table
    	-- corresponding to the u or v parametric direction of
    	-- the BSpline surface analysed by this algorithm.
    	-- The USplit and VSplit values are given in ascending
    	-- order and comprise the indices of the knots which
    	-- give the first and last isoparametric curves of the
    	-- surface in the corresponding parametric direction.
    	-- Use two consecutive values from the USplit table and
    	-- two consecutive values from the VSplit table as
    	-- arguments of the global function
    	-- SplitBSplineSurface (provided by the package
    	-- GeomConvert) to split the surface.
    	-- Exceptions
    	-- Standard_DimensionError if:
    	-- -   the array USplit was not created with the following bounds:
    	--   -   1 , and
    	--   -   the number of split knots in the u parametric
    	--    direction computed in this framework (as given
    	--    by the function NbUSplits); or
    	-- -   the array VSplit was not created with the following bounds:
    	--   -   1 , and
    	--   -   the number of split knots in the v parametric
    	--    direction computed in this framework (as given
    	--    by the function NbVSplits).
        raises DimensionError
            is static;
           

  USplitValue (me; UIndex : Integer)   returns Integer
        --- Purpose : Returns the split knot of index UIndex
    	-- to the split knots table for the u  parametric direction
    	-- computed in this framework. The returned value is
    	-- an index in the knots table relative to the u
    	--  parametric direction of the BSpline surface analysed by this algorithm.
    	-- Note: If UIndex is equal to 1, or to the number of split knots for the u
    	--  parametric direction computed in
    	-- this framework, the corresponding knot gives the
    	-- parameter of one of the bounding curves of the surface.
    	-- Exceptions
    	-- Standard_RangeError if UIndex  is less than 1 or greater than the number
    	-- of split knots for the u parametric direction computed in this framework.
     raises RangeError
     is static;


  VSplitValue (me; VIndex : Integer)   returns Integer
        --- Purpose :  Returns the split knot of index VIndex
    	-- to the split knots table for the v  parametric direction
    	-- computed in this framework. The returned value is
    	-- an index in the knots table relative to the v
    	--  parametric direction of the BSpline surface analysed by this algorithm.
    	-- Note: If UIndex is equal to 1, or to the number of split knots for the v
    	--  parametric direction computed in
    	-- this framework, the corresponding knot gives the
    	-- parameter of one of the bounding curves of the surface.
    	-- Exceptions
    	-- Standard_RangeError if VIndex  is less than 1 or greater than the number
    	-- of split knots for the v parametric direction computed in this framework.
            raises RangeError
     is static;

       
              
fields  

  usplitIndexes : HArray1OfInteger;
  vsplitIndexes : HArray1OfInteger;
  
end BSplineSurfaceKnotSplitting;
