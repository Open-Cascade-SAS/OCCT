-- Created on: 1994-06-01
-- Created by: Christian CAILLET
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class SetVersion5  from IGESSelect  inherits ModelModifier from IGESSelect

    ---Purpose : Sets IGES Version (coded in global parameter 23) to be at least
    --           IGES 5.1 . If it is older, it is set to IGES 5.1, and
    --           LastChangeDate (new Global n0 25) is added (current time)
    --           Else, it does nothing (i.e. changes neither IGES Version nor
    --           LastChangeDate)

uses AsciiString from TCollection,
     IGESModel, CopyTool, ContextModif

is

    Create returns mutable SetVersion5;
    ---Purpose : Creates an SetVersion5, which uses the system Date for Last
    --           Change Date

    Performing (me; ctx : in out ContextModif;
    	        target  : mutable IGESModel;
                TC      : in out CopyTool);
    ---Purpose : Specific action : only <target> is used : IGES Version (coded)
    --           is upgraded to 5.1 if it is older, and it this case the new
    --           global parameter 25 (LastChangeDate) is set to current time

    Label (me) returns AsciiString from TCollection;
    ---Purpose : Returns a text which is
    --           "Update IGES Version to 5.1"

end SetVersion5;
