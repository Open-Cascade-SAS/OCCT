-- Created on: 1993-04-06
-- Created by: Philippe DAUTRY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



package PGeom2d 

        ---Purpose :  This  package contains   the definition   of the
        --         geometric persistent objects such as point, vector,
        --         axis placement, curves, surfaces.
        --  
        --  All these entities are defined in 2D space.
        --  This package gives the possibility :
        --    . to create geometric objects with given or default field values,
        --    . to set field values,
        --    . to get field values.


uses PColStd, gp, PColgp, GeomAbs

is


  class Transformation from PGeom2d;


  deferred class Geometry from PGeom2d;


     deferred class Point from PGeom2d;
              class  CartesianPoint from PGeom2d;


     deferred class Vector from PGeom2d;
              class Direction from PGeom2d;
              class VectorWithMagnitude from PGeom2d;
     

     class AxisPlacement from PGeom2d;


     deferred class Curve from PGeom2d;

              class Line from PGeom2d;

              deferred class Conic from PGeom2d;
                       class Circle from PGeom2d;
                       class Ellipse from PGeom2d;
                       class Hyperbola from PGeom2d;
                       class Parabola from PGeom2d;

              deferred class BoundedCurve from PGeom2d;
                       class BezierCurve from PGeom2d;
                       class BSplineCurve from PGeom2d;
                       class TrimmedCurve from PGeom2d;

              class  OffsetCurve from PGeom2d;

end PGeom2d;
