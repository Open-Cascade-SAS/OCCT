-- Created on: 1994-12-09
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class NurbsConvert from BRepBuilderAPI inherits ModifyShape from BRepBuilderAPI

	---Purpose: Conversion of the complete geometry of a shape into
    	-- NURBS geometry. For example, all curves supporting
    	-- edges of the basis shape are converted into BSpline
    	-- curves, and all surfaces supporting its faces are
    	-- converted into BSpline surfaces.

uses 

    Shape             from TopoDS,
    Face              from TopoDS,
    ShapeModification from BRepBuilderAPI,
    ListOfShape       from TopTools
     
is

    Create returns NurbsConvert from BRepBuilderAPI;
    	---Purpose: Constructs a framework for converting the geometry of a
    	-- shape into NURBS geometry. Use the function Perform
    	-- to define the shape to convert.
    Create(S: Shape from TopoDS; 
           Copy: Boolean from Standard  =  Standard_False)

    	returns NurbsConvert from BRepBuilderAPI;
	---Purpose:  Builds a new shape by converting the geometry of the
    	-- shape S into NURBS geometry. Specifically, all curves
    	-- supporting edges of S are converted into BSpline
    	-- curves, and all surfaces supporting its faces are
    	-- converted into BSpline surfaces.
    	-- Use the function Shape to access the new shape.
    	-- Note: the constructed framework can be reused to
    	-- convert other shapes. You specify these with the
    	-- function Perform.

    Perform(me: in out; S   : Shape   from TopoDS; 
                        Copy: Boolean from Standard  =  Standard_False)

	---Purpose: Builds a new shape by converting the geometry of the
    	-- shape S into NURBS geometry.
    	-- Specifically, all curves supporting edges of S are
    	-- converted into BSpline curves, and all surfaces
    	-- supporting its faces are converted into BSpline surfaces.
    	-- Use the function Shape to access the new shape.
    	-- Note: this framework can be reused to convert other
    	-- shapes: you specify them by calling the function Perform again.
    	is static;

end NurbsConvert;
