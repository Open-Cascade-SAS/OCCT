-- Created on: 2004-06-24
-- Created by: STV
-- Copyright (c) 2004-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


private class ColorScale from V3d inherits ColorScale from Aspect

    ---Purpose: A colorscale class
uses

       --View           from V3d,
       LayerMgr         from V3d,
       LayerMgrPointer  from V3d,
       --Layer          from Visual3d,
       Color          from Quantity,
       ExtendedString from TCollection

is

       ---Category: Public

       Create(aMgr : LayerMgr from V3d)
       returns ColorScale from V3d;
       ---Purpose: Returns returns ColorScale from V3d.
    
       --View(me)
       --returns View from V3d;
       ---Purpose: Returns View from V3d.
    
       Display(me : mutable);

       Erase(me : mutable);

       IsDisplayed(me)
       returns Boolean from Standard;

       ---Category: Protected

       UpdateColorScale(me : mutable)
       is redefined protected;

       --BeginPaint(me : mutable)
       --returns Boolean from Standard
       --is redefined protected;

       --EndPaint(me : mutable)
       --returns Boolean from Standard
       --is redefined protected;

       PaintRect(me : mutable; X, Y, W, H : Integer from Standard;
                               aColor     : Color from Quantity;
                               aFilled    : Boolean from Standard = Standard_False)
       is redefined;

       PaintText(me : mutable; aText  : ExtendedString from TCollection;
                               X, Y   : Integer from Standard;
                               aColor : Color from Quantity)
       is redefined;

       TextWidth(me; aText : ExtendedString from TCollection)
       returns Integer from Standard
       is redefined;

       TextHeight(me; aText : ExtendedString from TCollection)
       returns Integer from Standard
       is redefined;

       TextSize( me;
                AText    : ExtendedString from TCollection;
                AHeight  : Integer from Standard;
                AWidth   : in out Integer from Standard;
                AnAscent : in out Integer from Standard;
                ADescent : in out Integer from Standard );

       DrawScale(me : mutable);

    ---Category: Private

       --Overlay(me)
       --returns Layer from Visual3d
       --is private;

fields

       --myView     : View from V3d;
       myLayerMgr : LayerMgrPointer from V3d;
       --myOverlay  : Layer from Visual3d;
       myDisplay  : Boolean from Standard;

end ColorScale;
