-- Created on: 1997-04-09
-- Created by: VAUTHIER Jean-Claude
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Real from PDataStd inherits Attribute from PDF

	---Purpose: 

uses Real from Standard

is

    Create returns mutable Real from PDataStd;

    
    Create (Value     : Real from Standard;
            Dimension : Integer from Standard)
    returns mutable Real from PDataStd;
    
    Get (me) returns Real from Standard;

    Set (me : mutable; V : Real from Standard);
    
    SetDimension (me : mutable; DIM : Integer from Standard);
    
    GetDimension (me)
    returns Integer from Standard;

fields

    myValue     : Real    from Standard;
    myDimension : Integer from Standard;

end Real;
