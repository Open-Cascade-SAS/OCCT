-- Created on: 1997-01-08
-- Created by: Robert COUBLANC
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ConnectedInteractive from AIS inherits InteractiveObject from AIS

	---Purpose: Defines an Interactive Object through a connection to
    	-- another Interactive   Object, which serves as a
    	-- reference, and which is located elsewhere in the viewer.
    	-- This allows you to use the Connected Interactive
    	-- Object without having to recalculate presentation,
    	-- selection or graphic structure. These are deduced
    	-- from your reference object.
    	-- The relation between the connected interactive object
    	-- and its source is generally one of geometric transformation. 
        -- AIS_ConnectedInteractive class doesn't support selection
        -- modes different from 0. Descendants should redefine ComputeSelection()
        -- method in order to handle other selection modes and generate connected
        -- sensitive entities properly. Refer to AIS_ConnectedShape class
        -- for exisiting implementation of a connected interactive object
        -- for AIS_Shape that supports all standard sub-shape selection modes.
    	-- Warning
    	-- An Interactive entity which is view (or projector)
    	-- dependent requires recalculation of views in hidden
    	-- parts mode depending on the position of the
    	-- projector in each view. You should derive the entity's
    	-- inheritance from ConnectedInteractive and redefine
    	-- its compute method to enable this type of calculation.

uses
    Location              from TopLoc,
    Transformation        from Geom,
    PresentationManager3d from PrsMgr,
    Presentation          from Prs3d,
    TypeOfPresentation3d  from PrsMgr,
    Selection             from SelectMgr,
    Projector             from Prs3d,
    KindOfInteractive     from AIS
raises
    NotImplemented from Standard

is

    Create (aTypeOfPresentation3d: TypeOfPresentation3d from PrsMgr = PrsMgr_TOP_AllView) 
    returns  mutable  ConnectedInteractive  from  AIS;
    	---Purpose:
    	-- Disconnects the previous view and sets highlight
    	-- mode to 0. This highlights the wireframe presentation
    	-- aTypeOfPresentation3d.
    	-- Top_AllView deactivates hidden line removal.
    
    Type(me) returns KindOfInteractive from AIS 
    is redefined virtual;
  	---Purpose: Returns KOI_Object

    Signature(me) returns Integer from Standard
    is redefined virtual;
	---Purpose: Returns 1


    Connect(me          : mutable; 
    	    anotherIObj : InteractiveObject from AIS) is virtual;
    	---Purpose: Establishes the connection between the Connected
    	-- Interactive Object, anotherIobj, and its reference
    	-- entity. If a previous connection with an Interactive
    	-- Object already exists, it is removed by Disconnect.
    	-- The second syntax also initiates the location of the
    	-- Connected Interactive Object.

    Connect(me:mutable;
    	    anotherIobj: InteractiveObject from AIS;
	    aLocation : Location from TopLoc) is virtual;
        ---Purpose: 
	    

    HasConnection(me) returns Boolean from Standard;
        ---C++: inline
    	---Purpose:
    	-- Returns true if there is a connection established
    	-- between the presentation and its source reference.
	
    ConnectedTo(me) returns any InteractiveObject from AIS;
     	---C++: inline
	---C++: return const&
    	---Purpose:
    	-- Returns the connection with the reference Interactive Object.

	    
    Disconnect(me:mutable);
	---Purpose: Clears the connection with a source reference. The
    	-- presentation will no longer be displayed.
    	-- Warning Must be done before deleting the presentation.

    Compute(me                   : mutable;
            aPresentationManager : PresentationManager3d from PrsMgr;
            aPresentation        : mutable Presentation from Prs3d;
            aMode                : Integer from Standard = 0)
	---Level: Public 
	---Purpose: Calculates the view aPresentation and its updates.
    	-- The latter are managed by aPresentationManager.
    	-- The display mode aMode is 0 by default.
    	--    this method is redefined virtual;
	--          when the instance is connected to another
    	--          InteractiveObject,this method doesn't
    	--          compute anything, but just uses the 
	--          presentation of this last object, with
	--          a transformation if there's one stored. 
    is redefined virtual private;

    Compute(me            : mutable;
    	    aProjector    : Projector from Prs3d;
    	    aTrsf         : Transformation from Geom;
	    aPresentation : mutable Presentation from Prs3d)
    is redefined;
	---Purpose: Computes the presentation according to a point of view
	--          given by <aProjector>. 
	--          To be Used when the associated degenerated Presentations 
	--          have been transformed by <aTrsf> which is not a Pure
	--          Translation. The HLR Prs can't be deducted automatically
	--          WARNING :<aTrsf> must be applied
	--           to the object to display before computation  !!!


    Compute(me:mutable;
    	        aProjector: Projector from Prs3d;
                aPresentation: mutable Presentation from Prs3d)
    is redefined;     
    
    ComputeSelection(me:mutable; aSelection :mutable Selection from SelectMgr;
                                 aMode      : Integer) is redefined virtual private;
	---Level: Public 
	---Purpose: Generates sensitive entities by copying 
        -- them from myReference selection, creates and sets an entity 
        -- owner for this entities and adds them to aSelection

    AcceptShapeDecomposition(me) returns Boolean from Standard is 
    redefined virtual;
	---C++: inline


    UpdateLocation(me:mutable) is redefined virtual;

    UpdateLocation(me:mutable;aSel:Selection from SelectMgr) is redefined virtual;
	---Purpose: For this class, the  location effect is treated in the
	--           compute   &     computeSelection  methods.  So     the
	--        UpdateLocation Methods are redefined to do nothing else

--   UpdateLocation(me:mutable;P : mutable Presentation from Prs3d) is redefined virtual;
    
fields

    myReference    : InteractiveObject from AIS is protected;
        ---Purpose: To have the time to Disconnect below, the old is kept for a while. 
    myOldReference : InteractiveObject from AIS is protected; 

end ConnectedInteractive;


