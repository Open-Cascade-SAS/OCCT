-- Created on: 1992-11-13
-- Created by: GG
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Package:     V3d.cdl
-- Modified:    stt:25-02-98; S3558: ajout ViewStdAdapter
--              ZOV - Mars 30 1998
--              stt:08-04-98; suppr. ViewStdAdapter
--              16-09-98 ; BGN : Ajout TypeOfTriedronEcho,
--                               TypeOfTriedronPosition.
--              22-09-98; BGN: S3989 (anciennement S3819): report
--                             dans Aspect des TypeOfTriedron*
-- Purpose:     Specifications provisoires

package V3d

        ---Purpose: This package contains the set of commands and services
        --          of the 3D Viewer. It provides a set of high level commands
        --          to control the views and viewing modes. This package is
        --          complementary to the Visual3D graphic package.
        --    Warning
        -- The CSF_WALKTHROUGH variable enables you to
        -- manage the perspective of the view in the viewer by
        -- defining setenv CSF_WALKTHROUGH "Yes".
        -- If you use the syntax unsetenv
        -- CSF_WALKTHROUGH, you undefine the variable
        -- (you make sure that the variable is deactivated). In
        -- this case, the eye is located outside the 3D bounding
        -- box of the view. This is the default behavior for
        -- managing the view perspective.


uses
        TColStd,
        Graphic3d,
        Visual3d,
        MMgt,
        TCollection,
        Quantity,
        Aspect,
        Image,
        gp,
        OSD,
        Font

is

        ------------------------------
        ---Category:  The extern types
        ------------------------------

        alias Coordinate is Length from Quantity;
        ---Purpose: User-defined coordinate in the reference plane of
        --          view (Projection or Mapping).


        alias Parameter is Parameter from Quantity;

        --------------------------
        --Category: The Exceptions
        --------------------------

        exception BadValue inherits OutOfRange;
        exception UnMapped inherits DomainError;

        -----------------------------
        ---Category: The Enumerations
        -----------------------------

        enumeration TypeOfView is ORTHOGRAPHIC,PERSPECTIVE
        end TypeOfView ;
        ---Purpose: Defines the type of projection of the view.

        enumeration TypeOfShadingModel is COLOR,MULTICOLOR,FLAT,GOURAUD,HIDDEN
              end TypeOfShadingModel ;
        ---Purpose:
        -- Defines the type of shading for the graphic object:
        -- -   V3d_COLOR: simple surface color,
        -- -   V3d_MULTICOLOR: interpolated colors,
        -- -   V3d_FLAT: flat shading,
        -- -   V3d_GOURAUD: Gouraud shading,
        -- -   V3d_HIDDEN: hidden line removal.

        enumeration  TypeOfSurfaceDetail  is  TEX_NONE, TEX_ENVIRONMENT, TEX_ALL
               end TypeOfSurfaceDetail;
        ---Purpose: Modes of visualization for objects in a view
        -- -   V3d_TEX_NONE: no texture mapping,
        -- -   V3d_TEX_ENVIRONMENT: environment mapping only,
        -- -   V3d_TEX_ALL: environment and texture mapping.

       enumeration TypeOfVisualization is      WIREFRAME,ZBUFFER
               end TypeOfVisualization ;
        ---Purpose: Determines the type of visualization in the view, either
        -- WIREFRAME or ZBUFFER (shading).

        enumeration TypeOfZclipping is     OFF,BACK,FRONT,SLICE
        --          Type "BACK"    Remove rear part
        --          Type "FRONT"   Remove front part
        --               "SLICE"   Keep the slice between the front plane
        --                         plane depth + half the thickness
        --                         and the rear plane
        --                         plane depth - half the thickness.
        --               "OFF"     ZClipping deactivated.
        end TypeOfZclipping ;
        ---Purpose: The available options are
        -- -   V3d_OFF: Zclipping (clipping executed in the
        --   depth of the view) is deactivated,
        -- -   V3d_BACK: back Zclipping is activated,
        -- -   V3d_FRONT: front Zclipping is activated,
        -- -   V3d_SLICE: both front and back Zclippings are activated.

        enumeration TypeOfLight is AMBIENT,DIRECTIONAL,POSITIONAL,SPOT
        end TypeOfLight ;
        ---Purpose: Determines the type of light.

        enumeration TypeOfUpdate is ASAP,WAIT
        end TypeOfUpdate ;
        ---Purpose: Determines the type of update of the view
        -- -   V3d_ASAP: as soon as possible. The view is updated immediately after a modification.
        -- -   V3d_WAIT: deferred. The view is updated when the Update function is called.

        enumeration TypeOfAxe is X,Y,Z
        end TypeOfAxe ;
        ---Purpose: Determines the axis type through the coordinates X, Y, Z.

        enumeration TypeOfOrientation is Xpos,Ypos,Zpos,Xneg,Yneg,Zneg,
            XposYpos,XposZpos,YposZpos,XnegYneg,XnegYpos,XnegZneg,
            XnegZpos,YnegZneg,YnegZpos,XposYneg,XposZneg,YposZneg,
            XposYposZpos,XposYnegZpos,XposYposZneg,XnegYposZpos,
            XposYnegZneg,XnegYposZneg,XnegYnegZpos,XnegYnegZneg
        end TypeOfOrientation ;
        ---Purpose: Determines the type of orientation.

        enumeration TypeOfRepresentation is SIMPLE,COMPLETE,PARTIAL,SAMELAST
        end TypeOfRepresentation;


        enumeration TypeOfPickLight is POSITIONLIGHT,SPACELIGHT,
            RADIUSTEXTLIGHT,ExtRADIUSLIGHT,IntRADIUSLIGHT,
            NOTHING
        end TypeOfPickLight;

        enumeration TypeOfPickCamera is POSITIONCAMERA,SPACECAMERA,
            RADIUSTEXTCAMERA,ExtRADIUSCAMERA,IntRADIUSCAMERA,
            NOTHINGCAMERA
        end TypeOfPickCamera;

    enumeration TypeOfProjectionModel is
        TPM_SCREEN,TPM_WALKTHROUGH
    end TypeOfProjectionModel;

        enumeration TypeOfBackfacingModel is
            TOBM_AUTOMATIC, TOBM_ALWAYS_DISPLAYED, TOBM_NEVER_DISPLAYED
        end TypeOfBackfacingModel;
        ---Purpose  : Modes of display of back faces in the view
        --
        --            TOBM_AUTOMATIC graphic's structure setting is in use
        --            TOBM_ALWAYS_DISPLAYED     force display of back faces
        --            TOBM_NEVER_DISPLAYED      disable display of back faces

        ------------------------
        ---Category: The classes
        ------------------------

        class Viewer;
        ---Purpose: Provides the services of a 3D viewer.

        class View;
        ---Purpose: Provides a set of services common to all types of view.

        class OrthographicView;
        ---Purpose: Services of an orthogonal view.

        class PerspectiveView;
        ---Purpose: Services of a perspective view.

        class LayerMgr;
        ---Purpose: Services of layer management.

        deferred class Light;
        ---Purpose: Provides services common to all types of luminous source.
        --          (base class for AmbientLight and PositionLight)


        class AmbientLight;
        ---Purpose: Services of ambient light sources.

        deferred class PositionLight;
        ---Purpose: Provides services common to Positional,Directional,Spot Lights.

        class PositionalLight;
        ---Purpose: Services of positional light sources.

        class DirectionalLight;
        ---Purpose: Services of directional light sources.

        class SpotLight;
        ---Purpose: Services of spot light sources.

        ---------------------------------
        ---Category: Instantiated classes
        ---------------------------------

        private class ListOfTransient;

        pointer ViewerPointer to Viewer from V3d;
        pointer ViewPointer to View from V3d;
        pointer LayerMgrPointer to LayerMgr from V3d;

        private class RectangularGrid;
        private class CircularGrid;

        private class ColorScale;
    private class ColorScaleLayerItem;

        ---------------------------------
        ---Category: Methodes de package
        ---------------------------------

        GetProjAxis( Orientation : TypeOfOrientation )
                                returns Vector from Graphic3d ;
        ---Purpose: Determines the orientation vector corresponding
        --          to the predefined orientation type.

        ArrowOfRadius ( garrow   : mutable Group from Graphic3d;
                        X0,Y0,Z0 : Coordinate;
                        DX,DY,DZ : Parameter;
                        Alpha    : PlaneAngle from Quantity;
                        Lng      : Parameter ) is protected;
        ---Level: Advanced
        ---Purpose: Compute the graphic structure of arrow.
        --          X0,Y0,Z0 : coordinate of the arrow.
        --          DX,DY,DZ : Direction of the arrow.
        --          Alpha    : Angle of arrow.
        --          Lng      : Length of arrow.

        CircleInPlane ( gcircle  : mutable Group from Graphic3d;
                        X0,Y0,Z0 : Coordinate;
                        VX,VY,VZ : Parameter;
                        Radius   : Parameter ) is protected;
        ---Level: Advanced
        ---Purpose: Compute the graphic structure of circle.
        --          X0,Y0,Z0 : Center of circle.
        --          VX,VY,VZ : Axis of circle.
        --          Radius   : Radius of circle.

        SwitchViewsinWindow(aPreviousView: View from V3d;
                            aNextView: View from V3d);


        DrawSphere(aViewer: Viewer from V3d; aRadius: Length from Quantity =1000);
        ---Purpose: test.

        PickGrid(aViewer: Viewer from V3d; aRadius: Length from Quantity =1000);
        ---Purpose: test.

        SetPlane(aViewer: Viewer from V3d; x1,y1,z1,x2,y2,z2: Length from Quantity);
        ---Purpose: test.

end V3d;

