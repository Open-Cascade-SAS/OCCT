-- Created on: 1996-12-05
-- Created by: Jean-Pierre COMBE/Odile Olivier
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PerpendicularRelation from AIS inherits Relation from AIS
    	---Purpose: A framework to display constraints of perpendicularity
    	-- between two or more interactive datums. These
    	-- datums can be edges or faces.
uses Shape                 from TopoDS,
     Presentation          from Prs3d,
     PresentationManager3d from PrsMgr,
     Selection             from SelectMgr,
     Pnt                   from gp,
     Dir                   from gp,
     Projector             from Prs3d,
     Transformation        from Geom,
     Plane                 from Geom

is
    Create (aFShape     : Shape          from TopoDS;
    	    aSShape     : Shape          from TopoDS;
	    aPlane      : Plane          from Geom)
	---Purpose:  Constructs an object to display constraints of
    	-- perpendicularity on shapes.
    	-- This object is defined by a first shape aFShape, a
    	-- second shape aSShape, and a plane aPlane.
    	-- aPlane is the plane of reference to show and test the
    	-- perpendicular relation between two shapes, at least
    	-- one of which has a revolved surface.
    returns mutable PerpendicularRelation from AIS;

    Create (aFShape     : Shape          from TopoDS;
    	    aSShape     : Shape          from TopoDS)
	---Purpose:  Constructs an object to display constraints of
    	-- perpendicularity on shapes.
    	-- This object is defined by a first shape aFShape and a
    	-- second shape aSShape.
    returns mutable PerpendicularRelation from AIS;

-- -- Methods from PresentableObject

    Compute(me            : mutable;
    	    aPresentationManager: PresentationManager3d from PrsMgr;
    	    aPresentation : mutable Presentation from Prs3d;
    	    aMode         : Integer from Standard= 0) 
    is redefined static private;
    
    Compute(me:mutable;
    	        aProjector: Projector from Prs3d;
                aPresentation: mutable Presentation from Prs3d)
    is redefined static private;     

    Compute(me            : mutable;
    	    aProjector    : Projector from Prs3d;
    	    aTrsf         : Transformation from Geom;
	    aPresentation : mutable Presentation from Prs3d)
    is redefined;
    	---Purpose: computes the presentation according to a point of view
    	--          given by <aProjector>. 
    	--          To be Used when the associated degenerated Presentations 
    	--          have been transformed by <aTrsf> which is not a Pure
    	--          Translation. The HLR Prs can't be deducted automatically
    	--          WARNING :<aTrsf> must be applied
    	--           to the object to display before computation  !!!

-- Methods from SelectableObject

    ComputeSelection(me         : mutable;
    	    	     aSelection : mutable Selection from SelectMgr;
    	    	     aMode      : Integer from Standard)is private;


--
--     Computation private methods
--

    ComputeTwoFacesPerpendicular(me: mutable;
    	    	    	         aPresentation : mutable Presentation from Prs3d)
    is private;
    
    ComputeTwoEdgesPerpendicular(me: mutable;
    	    	    	         aPresentation : mutable Presentation from Prs3d)
    is private;
    

fields

    myFAttach     : Pnt from gp;
    mySAttach     : Pnt from gp;
    
end PerpendicularRelation;


