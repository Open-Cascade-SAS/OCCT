-- Created on: 1995-10-06
-- Created by: Jing Cheng MEI
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class ShapeDirPresentation from DsgPrs

	---Purpose: A framework to define display of the normal to the
    	-- surface of a shape.

uses
    Shape  from TopoDS,
    Presentation from Prs3d,
    Drawer from Prs3d
    
is

    Add(myclass; prs: Presentation from Prs3d;
                 aDrawer: Drawer from Prs3d;
    	    	 shape: Shape from TopoDS; 
                 mode: Integer from Standard);
    	---Purpose: Adds the shape shape and the mode mode to the
    	-- presentation object prs.
    	-- The display attributes of the normal are defined by the
    	-- attribute manager aDrawer.
    	-- mode determines whether the first or the last point of
    	-- the normal is given to the presentation object. If the
    	-- first point: 0; if the last point, 1.
        
end ShapeDirPresentation;
