-- Created on: 1996-05-28
-- Created by: Denis PASCAL
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Angle from DrawDim inherits Dimension from DrawDim

	---Purpose: 

uses Face    from TopoDS,
     Display from Draw

is

    Create (plane1 : Face from TopoDS; 
            plane2 : Face from TopoDS)
    returns mutable Angle from DrawDim;
    
    Plane1 (me) returns Face from TopoDS;
	---C++: return const&

    Plane1 (me : mutable; plane : Face from TopoDS);

    Plane2  (me) returns Face from TopoDS;
	---C++: return const&

    Plane2 (me : mutable; plane : Face from TopoDS);    

    DrawOn (me; dis : in out Display);
    
fields

    myPlane1 : Face from TopoDS;
    myPlane2 : Face from TopoDS;
    
end Angle;

