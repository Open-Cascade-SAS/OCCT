-- Created on: 1995-03-13
-- Created by: Christian CAILLET
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



package XSControl

    ---Purpose : This package provides complements to IFSelect & Co for
    --           control of a session

uses Standard , MMgt, TCollection , TColStd, Dico,
     Interface, Transfer, IFSelect, Message,
     TopoDS,    TopTools, TopAbs ,   Geom, Geom2d, gp

is

    deferred class Controller;
    class TransferReader;
    class TransferWriter;

    class WorkSession;
    class SelectForTransfer;
    class SignTransferStatus;
    class ConnectedShapes;

    class Reader;
    class Writer;

    class Functions;
    class FuncShape;
    class Utils;
    class Vars;

    Session (pilot : SessionPilot from IFSelect) returns WorkSession from XSControl;
    ---Purpose : Returns the WorkSession of a SessionPilot, but casts it as
    --           from XSControl : it then gives access to Control & Transfers

    Vars    (pilot : SessionPilot from IFSelect) returns Vars from XSControl;
    ---Purpose : Returns the Vars of a SessionPilot, it is brought by Session
    --           it provides access to external variables

end XSControl;
