-- Created on: 1992-11-17
-- Created by: Christian CAILLET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class DispPerOne  from IFSelect  inherits Dispatch

    ---Purpose : A DispPerOne gathers all the input Entities into as many
    --           Packets as there Root Entities from the Final Selection,
    --           that is, one Packet per Entity

uses AsciiString from TCollection, Graph, SubPartsIterator

is

    Create returns mutable DispPerOne;
    ---Purpose : Creates a DispPerOne

    Label (me) returns AsciiString from TCollection;
    ---Purpose : Returns as Label, "One File per Input Entity"

    	--  --    Evaluation    --  --

    LimitedMax (me; nbent : Integer; max : out Integer) returns Boolean
    	is redefined;
    ---Purpose : Returns True, maximum limit is given as <nbent>

    PacketsCount (me; G : Graph; count : out Integer) returns Boolean
    	is redefined;
    ---Purpose : Returns True (count is easy to know) and count is the length
    --           of the input list (RootResult from FinalSelection)

    Packets (me; G : Graph; packs : in out SubPartsIterator);
    ---Purpose : Returns the list of produced Packets. It defines one Packet
    --           per Entity given by RootResult from the Final Selection.

end DispPerOne;
