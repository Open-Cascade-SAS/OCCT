-- Created on: 1993-01-11
-- Created by: CKY / Contract Toubro-Larsen ( Anand NATRAJAN )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class PartNumber from IGESAppli  inherits IGESEntity

        ---Purpose: defines PartNumber, Type <406> Form <9>
        --          in package IGESAppli
        --          Attaches a set of text strings that define the common
        --          part numbers to an entity being used to represent a
        --          physical component

uses

        HAsciiString from TCollection

is

        Create returns mutable PartNumber;

        -- Specific Methods pertaining to the class

        Init (me        : mutable; 
              nbPropVal : Integer;
              aGenName  : HAsciiString;
              aMilName  : HAsciiString;
              aVendName : HAsciiString;
              anIntName : HAsciiString);
        ---Purpose : This method is used to set the fields of the class
        --           PartNumber
        --       - nbPropVal : number of property values, always = 4
        --       - aGenName  : Generic part number or name
        --       - aMilName  : Military Standard (MIL-STD) part number
        --       - aVendName : Vendor part number or name
        --       - anIntName : Internal part number

        NbPropertyValues (me) returns Integer;
        ---Purpose : returns number of property values, always = 4

        GenericNumber (me) returns HAsciiString from TCollection;
        ---Purpose : returns Generic part number or name

        MilitaryNumber (me) returns HAsciiString from TCollection;
        ---Purpose : returns Military Standard (MIL-STD) part number

        VendorNumber (me) returns HAsciiString from TCollection;
        ---Purpose : returns Vendor part number or name

        InternalNumber (me) returns HAsciiString from TCollection;
        ---Purpose : returns Internal part number

fields

--
-- Class    : IGESAppli_PartNumber
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class PartNumber.
--
-- Reminder : A PartNumber instance is defined by :
--            - number of property values, always = 4
--            - Generic part number or name
--            - Military Standard (MIL-STD) part number
--            - Vendor part number or name
--            - Internal part number

        theNbPropertyValues : Integer;
        theGenericNumber    : HAsciiString;
        theMilitaryNumber   : HAsciiString;
        theVendorNumber     : HAsciiString;
        theInternalNumber   : HAsciiString;

end PartNumber;
