-- Created on: 1998-04-17
-- Created by: Andre LIEUTIER
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class  HPG0Constraint  from  NLPlate  inherits  HGPPConstraint from  NLPlate 
---Purpose: define a PinPoint G0  Constraint  used to load a Non Linear
--          Plate
uses
     XY from gp,
     XYZ from gp
     
is
    Create(UV : XY; Value : XYZ) returns mutable HPG0Constraint;
    -- create a G0 Constraint
    -- 

    SetUVFreeSliding(me: mutable; UVFree : Boolean) 
    is  redefined;
    -- If True, allow the UV value to  be modified during optimization
    --  this  is meaningless (has  no  effect) on   non G0 Constraints
    -- default is False
    -- 
    -- 

    SetIncrementalLoadAllowed(me: mutable; ILA : Boolean) 
    is  redefined;
    -- If True, allow the Constraint to be loaded incrementally during optimization
    -- default is False
    -- 


    UVFreeSliding(me)  returns  Boolean 
    is  redefined;
    -- If True, allow the UV value to be modified during optimization
    -- default is False
    -- 

    IncrementalLoadAllowed(me)  returns  Boolean 
    is redefined;
    -- If True, allow the Constraint to be loaded incrementally during optimization
    -- default is False
    -- 

    ActiveOrder(me)  returns  Integer 
    is   redefined; 
    --  returns the constraint active  order, i.e. the maximum between
    --  -- the initial constraint i.e 0 (for G0 Constraints)
    --  
    -- 

    IsG0(me) returns Boolean 
    is  redefined;

    G0Target(me) returns XYZ 
    ---C++: return const &
    is   redefined; 

fields
    myXYZTarget : XYZ from gp;
    UVIsFree : Boolean;
    IncrementalLoadingAllowed : Boolean;
end;
