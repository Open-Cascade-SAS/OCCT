-- Created on: 1998-10-15
-- Created by: Christian CAILLET
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class GraphCounter  from IFSelect    inherits SignCounter  from IFSelect

    ---Purpose : A GraphCounter computes values to be sorted with the help of
    --           a Graph. I.E. not from a Signature
    --           
    --           The default GraphCounter works with an Applied Selection (a
    --           SelectDeduct), the value is the count of selected entities
    --           from each input entities)

uses HSequenceOfTransient from TColStd,
     Graph from Interface, SelectDeduct from IFSelect

is

    Create (withmap  : Boolean = Standard_True;
            withlist : Boolean = Standard_False) returns GraphCounter;
    ---Purpose : Creates a GraphCounter, without applied selection

    Applied (me) returns SelectDeduct;
    ---Purpose : Returns the applied selection

    SetApplied (me : mutable; sel : SelectDeduct);
    ---Purpose : Sets a new applied selection

    AddWithGraph (me : mutable; list : HSequenceOfTransient; graph : Graph)
        is redefined virtual;
    ---Purpose : Adds a list of entities in the context given by the graph
    --           Default takes the count of entities selected by the applied
    --           selection, when it is given each entity of the list
    --           Can be redefined

fields

    theapplied : SelectDeduct;

end GraphCounter;
