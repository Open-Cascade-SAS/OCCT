-- Created on: 1995-12-04
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.





package RWStepVisual 

uses

	StepData, Interface, TCollection, TColStd, StepVisual

is


--class ReadWriteModule;

--class GeneralModule;

-- Removed from Rev2 to Rev4 : class RWAnnotationCurveOccurrence;
-- Removed from Rev2 to Rev4 : class RWAnnotationFillArea;
-- Removed from Rev2 to Rev4 : class RWAnnotationFillAreaOccurrence;
-- Removed from Rev2 to Rev4 : class RWAnnotationOccurrence;
-- Removed from Rev2 to Rev4 : class RWAnnotationSubfigureOccurrence;
-- Removed from Rev2 to Rev4 : class RWAnnotationSymbol;
-- Removed from Rev2 to Rev4 : class RWAnnotationSymbolOccurrence;
-- Removed from Rev2 to Rev4 : class RWAnnotationText;
-- Removed from Rev2 to Rev4 : class RWAnnotationTextOccurrence;
class RWAreaInSet;
class RWBackgroundColour;
class RWCameraImage;
class RWCameraModel;
class RWCameraModelD2;
class RWCameraModelD3;
class RWCameraUsage;
class RWColour;
class RWColourRgb;
class RWColourSpecification;
class RWContextDependentInvisibility;
class RWContextDependentOverRidingStyledItem;
-- Removed from CC1-Rev2 to CC1-Rev4, re-added CC2-Rev4 :
class RWCompositeText;
-- Removed from Rev2 to Rev4 : class RWCompositeTextWithAssociatedCurves;
-- Removed from Rev2 to Rev4 : class RWCompositeTextWithBlankingBox;
-- Removed from CC1-Rev2 to CC1-Rev4, re-added CC2-Rev4 :
class RWCompositeTextWithExtent;

class RWCurveStyle;
class RWCurveStyleFont;
class RWCurveStyleFontPattern;
-- Removed from Rev2 to Rev4 : class RWDefinedSymbol;
-- Removed from Rev2 to Rev4 : class RWDimensionCurve;
-- Removed from Rev2 to Rev4 : class RWDimensionCurveTerminator;
-- Removed from Rev2 to Rev4 : class RWDraughtingAnnotationOccurrence;
-- Removed from Rev2 to Rev4 : class RWDraughtingCallout;
class RWDraughtingModel; -- added for CAX-IF TR3
class RWDraughtingPreDefinedColour;
class RWDraughtingPreDefinedCurveFont;
-- Removed from Rev2 to Rev4 : class RWDraughtingSubfigureRepresentation;
-- Removed from Rev2 to Rev4 : class RWDraughtingSymbolRepresentation;
-- Removed from Rev2 to Rev4 : class RWDraughtingTextLiteralWithDelineation;
-- Removed from Rev2 to Rev4 : class RWDrawingDefinition;
-- Removed from Rev2 to Rev4 : class RWDrawingRevision;
--moved to RWStepBasic: class RWExternalSource;
class RWExternallyDefinedCurveFont;
-- Removed from Rev2 to Rev4 : class RWExternallyDefinedHatchStyle;
--moved to RWStepBasic: class RWExternallyDefinedItem;
-- Removed from Rev2 to Rev4 : class RWExternallyDefinedSymbol;
-- Removed from Rev2 to Rev4 : class RWExternallyDefinedTextFont;
-- Removed from Rev2 to Rev4 : class RWExternallyDefinedTileStyle;
class RWFillAreaStyle;
class RWFillAreaStyleColour;
-- Removed from Rev2 to Rev4 : class RWFillAreaStyleHatching;
-- Removed from Rev2 to Rev4 : class RWFillAreaStyleTileSymbolWithStyle;
-- Removed from Rev2 to Rev4 : class RWFillAreaStyleTiles;
class RWInvisibility;
class RWMechanicalDesignGeometricPresentationArea;
class RWMechanicalDesignGeometricPresentationRepresentation;
-- Removed from Rev2 to Rev4 : class RWMechanicalDesignPresentationArea;
class RWOverRidingStyledItem;
class RWPlanarBox;
class RWPlanarExtent;
class RWPointStyle;
class RWPreDefinedColour;
class RWPreDefinedCurveFont;
class RWPreDefinedItem;
-- Removed from Rev2 to Rev4 : class RWPreDefinedSymbol;
-- Removed from Rev2 to Rev4 : class RWPreDefinedTextFont;
class RWPresentationArea;
class RWPresentationLayerAssignment;
class RWPresentationRepresentation;
class RWPresentationSet;
class RWPresentationSize;
class RWPresentationStyleAssignment;
class RWPresentationStyleByContext;
class RWPresentationView;
-- Removed from Rev2 to Rev4 : class RWProductDataRepresentationView;
class RWStyledItem;
class RWSurfaceSideStyle;
class RWSurfaceStyleBoundary;
class RWSurfaceStyleControlGrid;
class RWSurfaceStyleFillArea;
class RWSurfaceStyleParameterLine;
class RWSurfaceStyleSegmentationCurve;
class RWSurfaceStyleSilhouette;
class RWSurfaceStyleUsage;
-- Removed from Rev2 to Rev4 : class RWSymbolColour;
-- Removed from Rev2 to Rev4 : class RWSymbolRepresentation;
-- Removed from Rev2 to Rev4 : class RWSymbolRepresentationMap;
-- Removed from Rev2 to Rev4 : class RWSymbolStyle;
-- Removed from Rev2 to Rev4 : class RWSymbolTarget;
class RWTemplate;
class RWTemplateInstance;
-- Removed from Rev2 to Rev4 : class RWTerminatorSymbol;
-- Removed from CC1-Rev2 to CC1-Rev4, re-added CC2-Rev4 :
class RWTextLiteral;
-- Removed from Rev2 to Rev4 : class RWTextLiteralWithAssociatedCurves;
-- Removed from Rev2 to Rev4 : class RWTextLiteralWithBlankingBox;
-- Removed from Rev2 to Rev4 : class RWTextLiteralWithDelineation;
-- Removed from Rev2 to Rev4 : class RWTextLiteralWithExtent;
-- Removed from CC1-Rev2 to CC1-Rev4, re-added CC2-Rev4 :
class RWTextStyle;
class RWTextStyleForDefinedFont;
class RWTextStyleWithBoxCharacteristics;
-- Removed from Rev2 to Rev4 : class RWTextStyleWithMirror;
class RWViewVolume;

    -- Added from Rev2 to Rev4
class RWPresentedItemRepresentation;
class RWPresentationLayerUsage;


	---Package Method ---

--	Init;
	---Purpose: enforced the initialisation of the  libraries

end RWStepVisual;
