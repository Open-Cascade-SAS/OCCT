-- Created on: 2001-08-28
-- Created by: data exchange team
-- Copyright (c) 2001-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Curve from ShapeCustom 

	---Purpose: Converts BSpline curve to periodic

uses

    Curve from Geom

is

    Create returns Curve from ShapeCustom;
    
    Create (C: Curve from Geom) returns Curve from ShapeCustom;
    
    Init (me: in out; C: Curve from Geom);
    
    ConvertToPeriodic (me: in out; substitute: Boolean; preci: Real = -1)
    returns Curve from Geom;
        ---Purpose: Tries to convert the Curve to the Periodic form
    	--          Returns the resulting curve
    	--          Works only if the Curve is BSpline and is closed with 
        --          Precision::Confusion()
    	--          Else, or in case of failure, returns a Null Handle
fields

    myCurve: Curve from Geom;

end Curve;
