--
-- File      :  ExternalReferenceFile.cdl
-- Created   :  Sat 9 Jan 1993
-- Author    : CKY / Contract Toubro-Larsen ( Anand NATRAJAN )
--
---Copyright : MATRA-DATAVISION  1993
--

class ExternalReferenceFile from IGESBasic  inherits IGESEntity

        ---Purpose: defines ExternalReferenceFile, Type <406> Form <12>
        --          in package IGESBasic
        --          References definitions residing in another file

uses

        HAsciiString from TCollection,
        HArray1OfHAsciiString from Interface

raises OutOfRange

is

        Create returns mutable ExternalReferenceFile;

        -- Specific Methods pertaining to the class

        Init (me : mutable; aNameArray : HArray1OfHAsciiString);
        ---Purpose : This method is used to set the fields of the class
        --           ExternalReferenceFile
        --       - aNameArray : External Reference File Names

        NbListEntries (me) returns Integer;
        ---Purpose : returns number of External Reference File Names

        Name (me; Index : Integer) returns HAsciiString from TCollection
        raises OutOfRange;
        ---Purpose : returns External Reference File Name
        -- raises exception if Index <= 0 or Index > NbListEntries()

fields

--
-- Class    : IGESBasic_ExternalReferenceFile
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class ExternalReferenceFile.
--
-- Reminder : A ExternalReferenceFile instance is defined by :
--            - External Reference File Names

        theNames : HArray1OfHAsciiString;

end ExternalReferenceFile;
