-- Created on: 1997-02-10
-- Created by: Robert COUBLANC
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class GraphicTool from AIS 

	---Purpose: 

uses
    Drawer          from Prs3d,
    TypeOfAttribute from AIS,
    NameOfColor     from Quantity,
    Color     	    from Quantity,
    TypeOfLine      from Aspect,
    MaterialAspect  from Graphic3d


is

    GetLineColor(myclass; aDrawer : Drawer from Prs3d; TheTypeOfAttributes :  TypeOfAttribute  from  AIS) 
    returns NameOfColor from Quantity; 
    
    GetLineColor(myclass; aDrawer : Drawer from Prs3d; 
		TheTypeOfAttributes :  TypeOfAttribute  from  AIS;
		TheLineColor: out Color from Quantity);
    
    GetLineWidth(myclass; aDrawer : Drawer from Prs3d; TheTypeOfAttributes :  TypeOfAttribute  from  AIS)
    returns Real from Standard;
    
    
    GetLineType (myclass; aDrawer : Drawer from Prs3d; TheTypeOfAttributes :  TypeOfAttribute  from  AIS)  
    returns TypeOfLine from Aspect;
    
    
    GetLineAtt(myclass;
    	       aDrawer : Drawer from Prs3d;
    	       TheTypeOfAttributes :  TypeOfAttribute  from  AIS; 
    	       aCol   : in out NameOfColor from Quantity;
	       aWidth : in out Real from Standard;
	       aTyp   : in out TypeOfLine from Aspect);
	       
	       
    GetInteriorColor(myclass;
    	    	    aDrawer : Drawer from Prs3d) 
    returns NameOfColor from  Quantity;

    GetInteriorColor(myclass;
    	    	    aDrawer : Drawer from Prs3d;
		    aColor: out Color from Quantity);

    GetMaterial(myclass; aDrawer:Drawer from Prs3d)
    returns MaterialAspect from Graphic3d;
	       
end GraphicTool;

