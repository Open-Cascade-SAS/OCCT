-- File:	StepRepr_RepresentationRelationshipWithTransformation.cdl
-- Created:	Tue Jun 30 18:09:19 1998
-- Author:	Christian CAILLET
--		<cky@heliox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1998


class RepresentationRelationshipWithTransformation  from StepRepr
    inherits ShapeRepresentationRelationship

    -- in principle, inherits RepresentationRelationship
    -- But <Shape>... only adds a constraint on a field, this allows to
    -- simplify the multiple inheritance between ShapeRR and RRWithTransf...

uses
     HAsciiString from TCollection,
     Representation from StepRepr,
     Transformation from StepRepr

is

    Create returns mutable RepresentationRelationshipWithTransformation;

    Init (me : mutable;
              aName : mutable HAsciiString from TCollection;
              aDescription : mutable HAsciiString from TCollection;
              aRep1 : mutable Representation from StepRepr;
              aRep2 : mutable Representation from StepRepr;
	      aTransf : Transformation);

    TransformationOperator (me) returns Transformation;
    SetTransformationOperator (me : mutable; aTrans : Transformation);

fields

    theTrans : Transformation;

end RepresentationRelationshipWithTransformation;
