-- Created on: 1992-03-27
-- Created by: Isabelle GRIGNON
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




generic class ZerParFunc from IntImp
    (ThePSurface     as any;
     ThePSurfaceTool as any)  -- as PSurfaceTool from IntImp (ThePSurface)


inherits FunctionSetWithDerivatives from math			       

	---Purpose: this function is associated to IWalking
	--          it's the definition of the line F(x,y,z)=0 
	--          where x=X(u,v),y=Y(u,v),z=Z(u,v)

uses Pnt                from gp,
     Dir                from gp,
     Vec                from gp,
     Dir2d              from gp,
     ConstIsoparametric from IntImp,
     Array1OfReal       from TColStd,
     Vector             from math,
     Matrix             from math

raises UndefinedDerivative from StdFail,     
       ConstructionError   from Standard
is

    Create 
    	---Purpose: Raises Construction Error
    	--          
    	returns ZerParFunc from IntImp;

    Create( S1,S2 : ThePSurface )

    	returns ZerParFunc from IntImp;


    NbVariables(me)

    	returns Integer from Standard

    	is static;


    NbEquations(me)

    	returns Integer from Standard

    	is static;


    Value(me : in out;X : in  Vector from math;
                      F : out Vector from math)

    	returns Boolean from Standard
    	is static;


    Derivatives(me : in out;X : in  Vector from math;
                            D : out Matrix from math)

    	returns Boolean from Standard
    	is static;


    Values(me : in out;
           X: in  Vector from math;
           F: out Vector from math; D: out Matrix from math)

    	returns Boolean from Standard
    	is static;

    
    ComputeParameters(me : in out; 
                      ChoixIso: ConstIsoparametric from IntImp; 
                      Param: Array1OfReal from TColStd;
                      UVap,BornInf,BornSup,Tolerance : out Vector from math)
    is static;

    
    Root(me)

    	---Purpose: returns somme des fi*fi

    	returns Real from Standard
	---C++: inline

    	is static;
    

    Point(me)

    	returns Pnt from gp
	---C++: inline

    	is static;
    

    IsTangent(me : in out; UVap : Vector from math;
    	    	    	   Param : out Array1OfReal from TColStd;
    	    	    	   BestChoix :  out ConstIsoparametric from IntImp)

    	returns Boolean from Standard
    	is static;
    

    Direction(me)

    	returns Dir from gp
	---C++: inline

    	raises UndefinedDerivative from StdFail
    	is static;
    

    DirectionOnS1(me)

    	returns Dir2d from gp
	---C++: inline

    	raises UndefinedDerivative from StdFail
    	is static;


    DirectionOnS2(me)

    	returns Dir2d from gp
	---C++: inline

    	raises UndefinedDerivative from StdFail
    	is static;
    

    AuxillarSurface1(me)

    	returns ThePSurface
	---C++: return const&
	---C++: inline

    	is static;


    AuxillarSurface2(me)

    	returns ThePSurface
	---C++: return const&
	---C++: inline

    	is static;

    
fields

    surf1      : Address from Standard; --- ThePSurface;
    surf2      : Address from Standard; --- ThePSurface;
    pntsol1    : Pnt     from gp; --point solution=milieu(pntsol1,pntsol2)
    pntsol2    : Pnt     from gp;
    f          : Real    from Standard[3];  -- equations
    compute    : Boolean from Standard;     --indicateur si tangence calculee
    tangent    : Boolean from Standard;     --indicateur si tangente
    tgduv      : Real    from Standard[4] ; --composante en u,en v de la
                   -- tangente ds plan tg du 1 ier et 2ieme caro
    dpuv       : Vec     from gp[4];        -- dp/du,dp/dv  sur 1ier et 2 ieme
                                            -- caro
    chxIso     : ConstIsoparametric from IntImp; -- indicateur sur l'iso 
                                                 -- constante
    paramConst : Real from Standard; -- parametre de l iso

    ua0,va0,ua1,va1 : Real from Standard; -- surf1 
    ub0,vb0,ub1,vb1 : Real from Standard; -- surf2  
    ures1,ures2,vres1,vres2 : Real from Standard; -- U et V Resolution
    
end ZerParFunc;

