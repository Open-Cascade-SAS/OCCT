-- Created on: 1993-03-23
-- Created by: BBL
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class ColorMapEntry from Aspect inherits Storable from Standard

	---Version: 0.0

	---Purpose: This class defines a colormap entry.
	--	    A colormap entry is an association between
	--	    a RGB object and a index in the colormap.
	---Keywords:
	---Warning:
	---References:

uses
	Color from Quantity

raises
	OutOfRange 	from Standard,
	BadAccess 	from Aspect

is
	Create
	returns ColorMapEntry from Aspect;
	---Level: Public
	---Purpose: Creates an unallocated colormap entry
	
	Create ( index : in Integer from Standard;
		 rgb : in Color from Quantity)
 	returns ColorMapEntry;
	---Level: Public
	---Purpose: Creates an allocated colormap entry

	Create ( entry : in ColorMapEntry from Aspect )
 	returns ColorMapEntry
	---Level: Public
	---Purpose: Creates an allocated colormap entry.
	--  Warning: Raises error if the colormap entry <entry>
	--	    is unallocated.
	raises BadAccess from Aspect;

	SetValue ( me: in out; index : in Integer from Standard;
			rgb : in Color from Quantity );
	---Level: Public
 	---Purpose: Sets colormap entry value and allocates it.
 
	SetValue ( me: in out; entry : in ColorMapEntry from Aspect);
	---Level: Public
 	---Purpose: Sets colormap entry value and allocates it.
	---C++: alias operator =
 
	SetColor ( me: in out; rgb : in Color from Quantity );
	---Level: Public
 	---Purpose: Sets color <rgb> of colormap entry.

	Color ( me : in ) returns Color from Quantity
	---Warning: Raises error if the colormap entry is unallocated .
	raises BadAccess from Aspect;
	---C++: return const & 

	SetIndex ( me: in out; index : in Integer from Standard);
	---Level: Public
 	---Purpose: Sets index value of a colormap entry.

	Index ( me : in ) returns Integer from Standard 
	---Warning: Raises error if the colormap entry is unallocated .
	raises BadAccess from Aspect;

	Free ( me : in out );
	---Level: Public
	---Purpose: Unallocates the colormap entry.

	IsAllocated ( me : in )
	returns Boolean from Standard;
	---Level: Public
	---Purpose: Returns True if the colormap entry is allocated.
	--  Warning: A colormap entry is allocated when the color and
	--	    the index is defined.

        Dump( me : in ) ;
	---Level: Internal

fields
	allocated 	: Boolean from Standard;
	mycolor		: Color from Quantity;
	myindex 	: Integer from Standard;
	myColorIsDef	: Boolean from Standard;
	myIndexIsDef	: Boolean from Standard;

end ColorMapEntry from Aspect;
