-- Created on: 1993-01-27
-- Created by: Philippe DAUTRY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class NumLinearRegularSweep from BRepSweep

	---Purpose: This  a generic  class  is  used   to build Sweept
	--          primitives   with    a  generating  "shape"  and a
	--          directing "line".
    	--          
    	--          The indexation and type analysis services required
    	--          for the generatrix are given by <Tool from BRepSweep>.
    	--          
    	--          The indexation and type analysis services required
    	--          for the directrix are given by <NumShapeTool from Sweep>.
    	--          
    	--          The iteration services required for the generatrix
    	--          are given by <Iterator from BRepSweep>.
    	--          
    	--          The iteration services required  for the directrix
    	--          are given by <NumShapeIterator from Sweep>.
	--          
	--          The topology is like a grid of shapes.  Each shape
	--          of the grid  must be addressable without confusion
	--          by one  or  two objects   from  the generating  or
	--          directing   shapes.  Here are  exemples of correct
	--          associations to address:
	--          
	--          - a vertex : GenVertex - DirVertex
	--          - an edge  : GenVertex - DirEdge
	--          -          : GenEdge   - DirVertex
	--          - a face   : GenEdge   - DirEdge
	--                       GenFace   - DirVertex
	--                       ...
    	--          
    	--          "GenObject" is used to identify an object from the
    	--          Generating     Shape,  and  "DirObject"  from  the
    	--          Directing Shape.  So may they   be  from different
    	--          types.
    	--          
    	--          The method Has... is given because in some special
    	--          cases, a vertex,    an  edge or   a   face may  be
    	--          geometricaly nonexistant or not usefull.

uses

    Orientation from TopAbs,
    Array2OfBoolean from TColStd,
    Shape from TopoDS,
    NumShape from Sweep,
    Builder from BRepSweep,
    Tool from BRepSweep,
    NumShapeTool from Sweep,
    Iterator from BRepSweep,
    NumShapeIterator from Sweep,
    Array2OfShape from TopTools,
    SequenceOfShape from TopTools

raises

    NoMoreObject from Standard,
    NoSuchObject from Standard,
    RangeError from Standard,
    DomainError from Standard


is


    -- """""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""

    Initialize(aBuilder  : Builder from BRepSweep;
	       aGenShape : Shape from TopoDS;
	       aDirWire  : NumShape from Sweep);
	---Purpose: Creates a NumLinearRegularSweep.    <aBuilder>  gives
	--          basic topological services.

    -- """""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""
    --  Deferred Methods supporting the creation of the geometric part.

    -- """""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""
    
    MakeEmptyVertex(me : in out; aGenV: Shape from TopoDS; aDirV: NumShape from Sweep)
    returns Shape from TopoDS is deferred;
	---Purpose: Builds the vertex addressed by [aGenV,aDirV], with its
	--          geometric part, but without subcomponents.
    ---C++ : alias "  Standard_EXPORT virtual ~BRepSweep_NumLinearRegularSweep();"
    
    MakeEmptyDirectingEdge(me: in out; aGenV: Shape from TopoDS; aDirE: NumShape from Sweep)
    returns Shape from TopoDS
	---Purpose: Builds the edge addressed by [aGenV,aDirE], with its
	--          geometric part, but without subcomponents.
    is deferred;
    
    MakeEmptyGeneratingEdge(me: in out; aGenE: Shape from TopoDS; aDirV: NumShape from Sweep)
    returns Shape from TopoDS
	---Purpose: Builds the edge addressed by [aGenE,aDirV], with its
	--          geometric part, but without subcomponents.
    is deferred;
    
    SetParameters(me         : in out; 
    	    	  aNewFace   : Shape from TopoDS; 
    	      	  aNewVertex : in out Shape from TopoDS;
    	    	  aGenF      : Shape from TopoDS; 
    	    	  aGenV      : Shape from TopoDS;
    	    	  aDirV      : NumShape from Sweep)
	---Purpose: Sets the  parameters of the new  vertex  on the new
	--          face. The new face and  new vertex where generated
	--          from aGenF, aGenV and aDirV .
    is deferred;
    
    SetDirectingParameter(me         : in out; 
    	    	          aNewEdge   : Shape from TopoDS; 
    	    	    	  aNewVertex : in out Shape from TopoDS;
    	    	          aGenV      : Shape from TopoDS;
    	    	          aDirE      : NumShape from Sweep; 
    	    	    	  aDirV      : NumShape from Sweep)
	---Purpose: Sets the  parameter of the new  vertex  on the new
	--          edge. The new edge and  new vertex where generated
	--          from aGenV aDirE, and aDirV.
    is deferred;

    SetGeneratingParameter(me         : in out; 
    	    	    	   aNewEdge   : Shape from TopoDS; 
                           aNewVertex : in out Shape from TopoDS;
    	    	    	   aGenE      : Shape from TopoDS; 
                           aGenV      : Shape from TopoDS;
    	    	    	   aDirV      : NumShape from Sweep)
	---Purpose: Sets the  parameter of the new  vertex  on the new
	--          edge. The new edge and  new vertex where generated
	--          from aGenE, aGenV and aDirV .
    is deferred;

    MakeEmptyFace(me       : in out; 
    	    	  aGenS    : Shape from TopoDS; 
    	    	  aDirS    : NumShape from Sweep)
    returns Shape from TopoDS
	---Purpose: Builds the face  addressed by  [aGenS,aDirS], with
	--          its geometric part, but without subcomponents. The
	--          couple aGenS, aDirS  can be a "generating face and
	--          a directing vertex"   or "a generating  edge and a
	--          directing  edge".
    is deferred;
    
    SetPCurve(me       : in out;
 	      aNewFace : Shape from TopoDS; 
              aNewEdge : in out Shape from TopoDS;
	      aGenF    : Shape from TopoDS; 
              aGenE    : Shape from TopoDS;
	      aDirV    : NumShape from Sweep;
    	      orien    : Orientation from TopAbs)
	 ---Purpose: Sets the PCurve for a new edge on a new face. The
	 --          new edge and  the  new face were generated  using
	 --          aGenF, aGenE and aDirV.
    is deferred;
    
    SetGeneratingPCurve(me       : in out;
    	    	    	aNewFace : Shape from TopoDS; 
                        aNewEdge : in out Shape from TopoDS;
			aGenE    : Shape from TopoDS; 
                        aDirE    : NumShape from Sweep;
			aDirV    : NumShape from Sweep;
   	                orien    : Orientation from TopAbs)

	 ---Purpose: Sets the PCurve for a new edge on a new face. The
	 --          new edge and  the  new face were generated  using
	 --          aGenE, aDirE and aDirV.
    is deferred;
    	    
    SetDirectingPCurve(me       : in out;
    	    	       aNewFace : Shape from TopoDS; 
                       aNewEdge : in out Shape from TopoDS;
		       aGenE    : Shape from TopoDS; 
		       aGenV    : Shape from TopoDS; 
                       aDirE    : NumShape from Sweep;
 	               orien    : Orientation from TopAbs)
		       
	 ---Purpose: Sets the PCurve for a new edge on a new face. The
	 --          new edge and  the  new face were generated  using
	 --          aGenE, aDirE and aGenV.
    is deferred;
    
    DirectSolid(me       : in out; 
    	    	aGenS    : Shape from TopoDS; 
    	    	aDirS    : NumShape from Sweep)
    returns Orientation from TopAbs
	---Purpose: Returns the Orientation of the  shell in the solid
	--          generated by the face aGenS  with  the edge aDirS.
	--          It is  REVERSED  if the surface is  swept  in  the
	--          direction of the normal.
    is deferred;
    
    GGDShapeIsToAdd (me;
    	    	     aNewShape    : Shape from TopoDS;
    	    	     aNewSubShape : Shape from TopoDS;
      	    	     aGenS        : Shape from TopoDS;
		     aSubGenS     : Shape from TopoDS;
    	    	     aDirS        : NumShape from Sweep)
    returns Boolean from Standard
	---Purpose: Returns   true   if  aNewSubShape    (addressed by
	--          aSubGenS  and aDirS)  must  be added  in aNewShape
	--          (addressed by aGenS and aDirS).
    is deferred;
    
    GDDShapeIsToAdd (me;
    	    	     aNewShape    : Shape from TopoDS;
    	    	     aNewSubShape : Shape from TopoDS;
      	    	     aGenS        : Shape from TopoDS;
    	    	     aDirS        : NumShape from Sweep;
   	    	     aSubDirS     : NumShape from Sweep)
    returns Boolean from Standard
	---Purpose: Returns   true   if  aNewSubShape    (addressed by
	--          aGenS  and aSubDirS)  must  be added  in aNewShape
	--          (addressed by aGenS and aDirS).
    is deferred;
    
    
    SeparatedWires (me;
    	    	     aNewShape    : Shape from TopoDS;
    	    	     aNewSubShape : Shape from TopoDS;
      	    	     aGenS        : Shape from TopoDS;
		     aSubGenS     : Shape from TopoDS;
    	    	     aDirS        : NumShape from Sweep)
    returns Boolean from Standard
	---Purpose: In  some  particular  cases  the   topology  of  a
	--          generated  face must be  composed  of  independant
	--          closed wires,  in this case  this function returns
	--          true.
    is deferred;
    

    SplitShell (me; aNewShape    : Shape from TopoDS)
    returns Shape from TopoDS
	---Purpose: In  some  particular  cases  the   topology  of  a
	--          generated  Shell must be  composed  of  independant
	--          closed Shells,  in this case  this function returns
	--          a Compound of independant Shells.
    is virtual;
    

    -- """"""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""
    --  Method coding the continuities on the edges between 2 faces
    -- """"""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""
    SetContinuity(me : in out; aGenS : Shape from TopoDS; aDirS : NumShape from Sweep)
       ---Purpose: Called to propagate the continuity of  every vertex
       --          between two edges of the  generating wire  aGenS on
       --          the generated edge and faces.
    is deferred;

        
    -- """""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""
    --  User end methods.
    --
    -- """""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""
    
    -- Shapes
    -- """"""

    HasShape(me; aGenS : Shape from TopoDS; aDirS : NumShape from Sweep) 
    	  returns Boolean from Standard
	---Purpose: Returns true   if aDirS   and aGenS  addresses   a
	--          resulting Shape. In some  specific cases the shape
	--          can  be    geometrically   inexsistant,  then this
	--          function returns false.
    is deferred;

    Shape(me: in out; aGenS : Shape from TopoDS; aDirS : NumShape from Sweep) 
    	  returns Shape from TopoDS
	---Purpose: Returns the resulting  Shape indexed by aDirS  and
	--          aGenS.
    is static;


    Shape(me: in out; aGenS : Shape from TopoDS) 
    	  returns Shape from TopoDS
	---Purpose: Returns  the resulting Shape  indexed by myDirWire
	--          and aGenS.
    is static;

    Shape(me: in out) 
    	  returns Shape from TopoDS
	---Purpose: Returns the resulting  Shape indexed by  myDirWire
	--          and myGenShape.
    is static;

    FirstShape(me: in out) 
    	  returns Shape from TopoDS
	---Purpose: Returns the resulting Shape  indexed by the  first
	--          Vertex  of myDirWire and myGenShape.
    is static;

    LastShape(me: in out) 
    	  returns Shape from TopoDS
	---Purpose: Returns the  resulting Shape  indexed by the  last
	--          Vertex of myDirWire and myGenShape.
    is static;
    

    FirstShape(me: in out; aGenS : Shape from TopoDS) 
    	  returns Shape from TopoDS
	---Purpose: Returns the resulting Shape  indexed by the  first
	--          Vertex  of myDirWire and aGenS.
    is static;

    LastShape(me: in out; aGenS : Shape from TopoDS) 
    	  returns Shape from TopoDS
	---Purpose: Returns the  resulting Shape  indexed by the  last
	--          Vertex of myDirWire and aGenS.
    is static;
    
    
    Closed(me) returns Boolean from Standard is static;

fields

    -- Topology builder.

    myBuilder  : Builder from BRepSweep is protected;  

    -- Generating shape
    
    myGenShape : Shape from TopoDS is protected;

    -- Directing line
    
    myDirWire  : NumShape from Sweep is protected;

    -- shape tools.

    myGenShapeTool   : Tool from BRepSweep is protected;
    myDirShapeTool   : NumShapeTool from Sweep is protected;

    -- Array of built objects (NbGShapes,NbDShapes).
    myShapes       : Array2OfShape from TopTools is protected;

    -- Array of built objects flags (NbGShapes,NbDShapes).
    myBuiltShapes : Array2OfBoolean from TColStd is protected;
    	    	
end NumLinearRegularSweep;
