-- Created on: 1991-03-29
-- Created by: Remi GILET
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

generic class Circ2d2TanOn from GccGeo (
    TheCurve         as any; --
    TheTool          as any; --
    TheQCurve        as any; -- as QualifiedCurve from GccEnt
    	    	             --                  (TheCurve)
    TheParGenCurve   as any; -- as ParGenCurve from GccGeo 
    	    	    	     --               (TheCurve)
    TheHParGenCurve  as Transient;
    TheCurvePGTool   as any; -- as CurvePGTool from GccGeo 
    	    	    	     --               (Thecurve,
    	    	       	     --                TheTool,
    	    	       	     --                TheParGenCurve)
    TheIntConicCurve as any) -- as TheIntConicCurveOfGOffsetInter from IntCurve
    	    	    	     --                            (TheParGenCurve,
    	    	    	     --                             TheCurvePGTool)


	---Purpose: This class implements the algorithms used to 
	--          create 2d circles TANgent to 2 entities and 
	--          having the center ON a curve.
	--          The order of the tangency argument is always
	--          QualifiedCirc, QualifiedLin, QualifiedCurv, Pnt2d. 
	--          the arguments are :
	--            - The two tangency arguments (lines, circles or points).
	--            - The center line (a curve).
	--            - The parameter for each tangency argument which 
	--            is a curve.
	--            - The tolerance.

-- inherits Entity from Standard

uses Pnt2d            from gp,
     Lin2d            from gp,
     Circ2d           from gp,  
     QualifiedCirc    from GccEnt,
     QualifiedLin     from GccEnt,
     Array1OfCirc2d   from TColgp,
     Array1OfPnt2d    from TColgp,
     Array1OfInteger  from TColStd,
     Array1OfReal     from TColStd,
     Position         from GccEnt,
     Array1OfPosition from GccEnt
     
raises NotDone      from StdFail,
       BadQualifier from GccEnt,
       OutOfRange   from Standard

is

Create(Qualified1 :        QualifiedCirc from GccEnt  ;
       Qualified2 :        QualifiedCirc from GccEnt  ;
       OnCurv     :        TheCurve                   ;
       Tolerance  :        Real          from Standard) returns Circ2d2TanOn
    ---Purpose: This method implements the algorithms used to 
    --          create 2d circles TANgent to two 2d circles and 
    --          having the center ON a curve.
raises BadQualifier from GccEnt;

Create(Qualified1 :        QualifiedCirc from GccEnt  ;
       Qualified2 :        QualifiedLin  from GccEnt  ;
       OnCurv     :        TheCurve                   ;
       Tolerance  :        Real          from Standard) returns Circ2d2TanOn
    ---Purpose: This method implements the algorithms used to 
    --          create 2d circles TANgent to a 2d circle and a 2d line
    --          having the center ON a curve.
raises BadQualifier from GccEnt;

Create(Qualified1 :        QualifiedCirc from GccEnt  ;
       Point2     :        Pnt2d         from gp      ;
       OnCurv     :        TheCurve                   ;
       Tolerance  :        Real          from Standard) returns Circ2d2TanOn
    ---Purpose: This method implements the algorithms used to 
    --          create 2d circles TANgent to a 2d circle and a point
    --          having the center ON a curve.
raises BadQualifier from GccEnt;

Create(Qualified1 :        QualifiedLin  from GccEnt  ;
       Qualified2 :        QualifiedLin  from GccEnt  ;
       OnCurv     :        TheCurve                   ;
       Tolerance  :        Real          from Standard) returns Circ2d2TanOn
    ---Purpose: This method implements the algorithms used to 
    --          create 2d circles TANgent to two 2d lines
    --          having the center ON a curve.
raises BadQualifier from GccEnt;

Create(Qualified1 :        QualifiedLin  from GccEnt  ;
       Qualified2 :        Pnt2d         from gp      ;
       OnCurv     :        TheCurve                   ;
       Tolerance  :        Real          from Standard) returns Circ2d2TanOn
    ---Purpose: This method implements the algorithms used to 
    --          create 2d circles TANgent to a 2d line and a point
    --          having the center ON a 2d line.
raises BadQualifier from GccEnt;

Create(Point1     :        Pnt2d         from gp      ;
       Point2     :        Pnt2d         from gp      ;
       OnCurv     :        TheCurve                   ;
       Tolerance  :        Real          from Standard) returns Circ2d2TanOn ;
    ---Purpose: This method implements the algorithms used to 
    --          create 2d circles TANgent to two points
    --          having the center ON a 2d line.

-- ....................................................................

IsDone(me) returns Boolean from Standard
is static;
    ---Purpose: This method returns True if the construction 
    --          algorithm succeeded.

NbSolutions(me) returns Integer from Standard
    ---Purpose: This method returns the number of solutions.
raises NotDone
is static;
    ---Purpose: It raises NotDone if the construction algorithm 
    --          didn't succeed.

ThisSolution(me ; Index : Integer) returns Circ2d from gp 
    ---Purpose: Returns the solution number Index and raises OutOfRange 
    --  	exception if Index is greater than the number of solutions.
    --          Be careful: the Index is only a way to get all the 
    --          solutions, but is not associated to those outside the 
    --          context of the algorithm-object.
raises OutOfRange, NotDone
is static;
    ---Purpose: It raises NotDone if the construction algorithm 
    --          didn't succeed.
    --          It raises OutOfRange if Index is greater than the 
    --          number of solutions.

WhichQualifier(me                                  ;
    	       Index   :     Integer  from Standard;
	       Qualif1 : out Position from GccEnt  ;
	       Qualif2 : out Position from GccEnt  )
raises OutOfRange, NotDone
is static;
    ---Purpose: It returns the informations about the qualifiers of 
    --          the tangency 
    --          arguments concerning the solution number Index.
    --          It returns the real qualifiers (the qualifiers given to the 
    --          constructor method in case of enclosed, enclosing and outside 
    --          and the qualifiers computedin case of unqualified).

Tangency1(me                                     ;
          Index         : Integer   from Standard;
          ParSol,ParArg : out Real  from Standard;
          PntSol        : out Pnt2d from gp      )
    ---Purpose: Returns informations about the tangency point between the 
    --          result number Index and the first argument.
    --          ParSol is the intrinsic parameter of the point on the 
    --          solution curv.
    --          ParArg is the intrinsic parameter of the point on the 
    --          argument curv.
    --          PntSol is the tangency point on the solution curv.
    --          PntArg is the tangency point on the argument curv.
raises OutOfRange, NotDone
is static;
    ---Purpose: It raises NotDone if the construction algorithm 
    --          didn't succeed.
    --          It raises OutOfRange if Index is greater than the 
    --          number of solutions.

Tangency2(me                                     ;
          Index         : Integer   from Standard;
          ParSol,ParArg : out Real  from Standard;
          PntSol        : out Pnt2d from gp      )
    ---Purpose: Returns informations about the tangency point between the 
    --          result number Index and the second argument.
    --          ParSol is the intrinsic parameter of the point on the 
    --          solution curv.
    --          ParArg is the intrinsic parameter of the point on the 
    --          argument curv.
    --          PntSol is the tangency point on the solution curv.
    --          PntArg is the tangency point on the argument curv.
raises OutOfRange, NotDone
is static;
    ---Purpose: It raises NotDone if the construction algorithm 
    --          didn't succeed.
    --          It raises OutOfRange if Index is greater than the 
    --          number of solutions.

CenterOn3 (me                                     ;
           Index         : Integer   from Standard;
           ParArg        : out Real  from Standard;
           PntSol        : out Pnt2d from gp      )
    ---Purpose: Returns informations about the center (on the curv) 
    --          of the result.
    --          ParArg is the intrinsic parameter of the point on 
    --          the argument curv.
    --          PntSol is the center point of the solution curv.
raises OutOfRange, NotDone
is static;
    ---Purpose: It raises NotDone if the construction algorithm 
    --          didn't succeed.
    --          It raises OutOfRange if Index is greater than the 
    --          number of solutions.

IsTheSame1(me                           ;
           Index : Integer from Standard) returns Boolean from Standard
    ---Purpose: Returns True if the solution number Index is equal to 
    --          the first argument and False in the other cases.
raises OutOfRange, NotDone
is static;
    ---Purpose: It raises NotDone if the construction algorithm 
    --          didn't succeed.
    --          It raises OutOfRange if Index is greater than the 
    --          number of solutions.

IsTheSame2(me                           ;
           Index : Integer from Standard) returns Boolean from Standard
    ---Purpose: Returns True if the solution number Index is equal to 
    --          the second argument and False in the other cases.
raises OutOfRange, NotDone
is static;
    ---Purpose: It raises NotDone if the construction algorithm 
    --          didn't succeed.
    --          It raises OutOfRange if Index is greater than the 
    --          number of solutions.

fields

    WellDone : Boolean from Standard;
    ---Purpose: True if the algorithm succeeded.

    NbrSol   : Integer from Standard;
    ---Purpose: Number of solutions.

    cirsol   : Array1OfCirc2d from TColgp;
    ---Purpose: The solutions.

    qualifier1 : Array1OfPosition from GccEnt;
    ---Purpose: The qualifiers of the first argument.

    qualifier2 : Array1OfPosition from GccEnt;
    ---Purpose: The qualifiers of the second argument.

    TheSame1 : Array1OfInteger from TColStd;
    ---Purpose: 1 if the solution and the first argument are the same 
    --          (2 circles).
    --          If R1 is the radius of the first argument and Rsol the radius 
    --          of the solution and dist the distance between the two centers,
    --          we consider the two circles are identical if R1+dist-Rsol is 
    --          less than Tolerance.
    --          0 in the other cases.

    TheSame2 : Array1OfInteger from TColStd;
    ---Purpose: 1 if the solution and the second argument are the same 
    --          (2 circles).
    --          If R2 is the radius of the second argument and Rsol the radius 
    --          of the solution and dist the distance between the two centers,
    --          we consider the two circles are identical if R2+dist-Rsol is 
    --          less than Tolerance.
    --          0 in the other cases.

    pnttg1sol   : Array1OfPnt2d from TColgp;
    ---Purpose: The tangency point between the solution and the first 
    --          argument on the solution.

    pnttg2sol   : Array1OfPnt2d from TColgp;
    ---Purpose: The tangency point between the solution and the second 
    --          argument on the solution.

    pntcen   : Array1OfPnt2d from TColgp;
    ---Purpose: The center point of the solution on the third argument.

    par1sol   : Array1OfReal from TColStd;
    ---Purpose: The parameter of the tangency point between the solution 
    --          and the first argument on the solution.

    par2sol   : Array1OfReal from TColStd;
    ---Purpose: The parameter of the tangency point between the solution 
    --          and the second argument on the solution.

    pararg1   : Array1OfReal from TColStd;
    ---Purpose: The parameter of the tangency point between the solution 
    --          and the first argument on the first argument.

    pararg2   : Array1OfReal from TColStd;
    ---Purpose: The parameter of the tangency point between the solution 
    --          and the second argument on the second argument.

    parcen3   : Array1OfReal from TColStd;
    ---Purpose: The parameter of the center point of the solution on the 
    --          second argument.

end Circ2d2TanOn;
