-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class OrientedFace from StepShape 

inherits Face from StepShape 

uses

	Boolean from Standard, 
	HArray1OfFaceBound from StepShape, 
	FaceBound from StepShape, 
	HAsciiString from TCollection
is

	Create returns OrientedFace;
	---Purpose: Returns a OrientedFace


	Init (me : mutable;
	      aName : HAsciiString from TCollection;
	      aBounds : HArray1OfFaceBound from StepShape) is redefined;

	Init (me : mutable;
	      aName : HAsciiString from TCollection;
	      aFaceElement : Face from StepShape;
	      aOrientation : Boolean from Standard) is virtual;

	-- Specific Methods for Field Data Access --

	SetFaceElement(me : mutable; aFaceElement : Face);
	FaceElement (me) returns Face;
	SetOrientation(me : mutable; aOrientation : Boolean);
	Orientation (me) returns Boolean;
	SetBounds(me : mutable; aBounds : HArray1OfFaceBound) is redefined;
	Bounds (me) returns HArray1OfFaceBound is redefined;
	BoundsValue (me; num : Integer) returns FaceBound is redefined;
	NbBounds (me) returns Integer is redefined;

fields

	faceElement : Face from StepShape;
	orientation : Boolean from Standard;

 -- 
 -- NB : field <bounds> inherited from classe <face> is redeclared.
 --      it shall appears in a physical file as a *.
 --

end OrientedFace;
