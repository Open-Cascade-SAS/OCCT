-- Created on: 1990-12-11
-- Created by: Remi Lequette
-- Copyright (c) 1990-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Update:      Frederic Maupas


class HShape from PTopoDS inherits ExternShareable from ObjMgt

    ---Purpose: The PTopoDS_HShape is the Persistent view of a TopoDS_Shape.
  -- This can be a vertex, an edge, a wire, a face, a shell, a solid and so on.
 -- It can be shared by other objects.
    --  a  HShape contains :
    --          
    --          - a reference to a TShape.
    --          
    --          - a Location  to put the TShape in  a local coordinate
    --          system.
    --          
    --          - an Orientation.
    --          
    --          It inherits from ExternShareable, so that it can be shared
    --          by other objects located outside the container.
    
uses

    Orientation   from TopAbs,
    TShape        from PTopoDS,
    Location      from PTopLoc
    
is
    Create returns mutable HShape from PTopoDS;
    ---Level: Internal 

    TShape(me) returns any TShape from PTopoDS
    ---Level: Internal 
    is static;

    TShape(me : mutable; T : TShape from PTopoDS)
    ---Level: Internal 
    is static;

    Location(me) returns Location from PTopLoc
    ---Level: Internal 
    is static;
	
    Location(me : mutable; L : Location from PTopLoc)
    ---Level: Internal 
    is static;
	
    Orientation(me) returns Orientation from TopAbs
    ---Level: Internal 
    is static;

    Orientation(me: mutable; O : Orientation from TopAbs)
    ---Level: Internal 
    is static;
    
fields
    myTShape   : TShape      from PTopoDS;
    myLocation : Location    from PTopLoc;
    myOrient   : Orientation from TopAbs;

end HShape;
