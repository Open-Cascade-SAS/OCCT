-- Created on: 1998-06-03
-- Created by: data exchange team
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



package ShapeUpgrade 

    	---Purpose:  This package provides tools
    	-- for splitting and converting shapes by some criteria. It
    	-- provides modifications of the kind when one topological
    	-- object can be converted or splitted to several ones. In
    	-- particular this package contains high level API classes which perform: 
    	--      converting geometry of shapes up to given continuity, 
    	--      splitting revolutions by U to segments less than given value, 
    	--      converting to beziers, 
    	--      splitting closed faces. 
    
uses
    gp,
    Geom,
    Geom2d,
    GeomAbs,
    Adaptor3d,
    GeomAdaptor,
    Geom2dAPI,
    TopLoc,
    TColStd,
    TColGeom,
    TColGeom2d,
    TCollection,
    TopoDS,
    TopTools,
    TopAbs,
    ShapeExtend,
    ShapeBuild,
    ShapeAnalysis,
    BRepBuilderAPI

is

    --- Instanciation of generic classes (tools)
    
    private class Tool;
    
    	class EdgeDivide;
	
	    class ClosedEdgeDivide;
	    
    	class WireDivide;
    
    	class FaceDivide;
    
    	    class ClosedFaceDivide;
	    class FaceDivideArea;
    
    class ShapeDivide;
    	class ShapeDivideArea;
    
    class ShapeDivideContinuity;    
    	---Purpose: API Tool for converting shapes with C0 geometry into C1 ones
    
    class ShapeDivideAngle;
    	---Purpose: API Class for splitting revolutions to segments less than 90

    class ShapeConvertToBezier;
    	---Purpose: API Class for convering curves to beziers.
	
    class ShapeDivideClosed;
    	---Purpose:
	
    class ShapeDivideClosedEdges;
    	---Purpose:
	
    class SplitCurve;
	class SplitCurve2d;
    	    class SplitCurve2dContinuity;
	    class ConvertCurve2dToBezier;
    	class SplitCurve3d;
    	    class SplitCurve3dContinuity;
	    class ConvertCurve3dToBezier;
	
    class SplitSurface;
    	class SplitSurfaceContinuity;
	class SplitSurfaceAngle;
	class ConvertSurfaceToBezierBasis;
	class SplitSurfaceArea;
	
    class ShellSewing;
    	---Purpose: Provides access to a sewing algorithms from BRepOffsetAPI
    class FixSmallCurves;
    ---Purpose:
    class FixSmallBezierCurves;
    ---Purpose:
    
    class RemoveLocations;
    ---Purpose: Removes all locations sub-shapes of specified shape
    
    class RemoveInternalWires;
    ---Purpose: Removes all internal wires having area less than specified min area
    
    C0BSplineToSequenceOfC1BSplineCurve (BS   : BSplineCurve from Geom;
    	    	    	    	         seqBS: out HSequenceOfBoundedCurve from TColGeom)
    returns Boolean;
				      
    C0BSplineToSequenceOfC1BSplineCurve (BS   : BSplineCurve from Geom2d;
    	    	    	    	         seqBS: out HSequenceOfBoundedCurve from TColGeom2d)
    returns Boolean;
    --- Purpose: Converts C0 B-Spline curve into sequence of C1 B-Spline curves.
    --           This method splits B-Spline at the knots with multiplicities
    --           equal to degree, i.e. unlike method
    --           GeomConvert::C0BSplineToArrayOfC1BSplineCurve this one does not
    --           use any tolerance and therefore does not change the geometry of
    --           B-Spline.
    --           Returns True if C0 B-Spline was successfully splitted, else
    --           returns False (if BS is C1 B-Spline).

end ShapeUpgrade;
