-- Created on: 1997-03-16
-- Created by: SMO
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



package TPrsStd 

	---Purpose: The visualization attribute implements the
    	-- Application Interactive Services in the context
    	-- of Open CASCADE Application Framework.


    ---Category: GUID 
    --           04fb4d05-5690-11d1-8940-080009dc3333   TPrsStd_AISViewer
    --           04fb4d00-5690-11d1-8940-080009dc3333	TPrsStd_AISPresentation
   
uses
    Standard,
    TCollection,
    TColStd,
    MMgt,
    Quantity,
    Graphic3d,
    AIS,
    V3d,    
    TDF,
    TDataXtd,
    Geom,
    TopoDS,
    gp
    
    
is


    ---Category: Attributes 
    --           ==========
    
    class AISViewer;
    
    class AISPresentation;  

    ---Category : Drivers to build and/or update AIS objects
    --            ==========================================

    deferred class Driver;
      class PointDriver ;         -- to display Point
      class AxisDriver ;          -- to display Axis
      class PlaneDriver ;         -- to display Plane
      class GeometryDriver;       -- to display Geometry
      class ConstraintDriver;     -- to display Constraint
      class NamedShapeDriver;     -- to display NamedShape
    
    class DriverTable ;               
    
    ---Category: Tools
    --           =====

    class ConstraintTools;

    class DataMapOfGUIDDriver
    instantiates DataMap from TCollection(GUID      from Standard, 
	    	 		       	  Driver from TPrsStd, 
				          GUID      from Standard); 
end TPrsStd;

