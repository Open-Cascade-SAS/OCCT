-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package PColStd 

uses PCollection,
     TCollection,
     TColStd

is


--                             Instantiations de PCollection          --
--                             *****************************          --
------------------------------------------------------------------------

--
--       Instantiations HSequence (Integer,Real,Persistent,
--                                 HAsciiString,
--                                 HExtendedString)
--       **************************************************
--       
class HSequenceOfInteger instantiates 
           HSequence from PCollection(Integer);
class HSequenceOfReal instantiates 
           HSequence from PCollection(Real);
class HSequenceOfPersistent instantiates 
           HSequence from PCollection(Persistent);
class HSequenceOfHAsciiString instantiates 
           HSequence from PCollection(HAsciiString from PCollection);
class HSequenceOfHExtendedString instantiates 
           HSequence from PCollection(HExtendedString from PCollection);
--
--       Instantiations HSingleList (Integer,Real,Persistent)
--       *****************************************************
--       
class HSingleListOfInteger instantiates 
           HSingleList from PCollection(Integer);
class HSingleListOfReal instantiates 
           HSingleList from PCollection(Real);
class HSingleListOfPersistent instantiates 
           HSingleList from PCollection(Persistent);
--       Instantiations HDoubleList (Integer,Real,Persistent)
--       *********************************************
--       
class HDoubleListOfInteger instantiates 
           HDoubleList from PCollection(Integer);
class HDoubleListOfReal instantiates 
           HDoubleList from PCollection(Real);
class HDoubleListOfPersistent instantiates 
           HDoubleList from PCollection(Persistent);
--
--       Instantiations HArray1 (Integer,Real,Persistent)
--       ****************************************************
--       
    class HArray1OfInteger instantiates 
                        HArray1 from PCollection(Integer);

    class HArray1OfReal instantiates 
                        HArray1 from PCollection(Real);

    class HArray1OfExtendedString instantiates 
                        HArray1 from PCollection(HExtendedString from PCollection);

    class HArray1OfPersistent instantiates 
                        HArray1 from PCollection(Persistent);
--
--       Instantiations HArray2 (Integer,Real,Persistent)
--       ****************************************************
--       
    class HArray2OfInteger instantiates
                        HArray2 from PCollection(Integer);
    class HArray2OfReal instantiates 
                        HArray2 from PCollection(Real);
    class HArray2OfPersistent instantiates 
                        HArray2 from PCollection(Persistent);

--       Instantiations Hash (Integer)
--       *****************************
--
class HOfInteger instantiates Hash from PCollection(Integer);
class HOfReal instantiates Hash from PCollection(Real);
class HOfAsciiString instantiates Hash from PCollection(HAsciiString from PCollection);
---Purpose: Hash on the Handle.
class HashAsciiString;
---Purpose: Hash on the string.
class HOfExtendedString instantiates Hash from PCollection(HExtendedString from PCollection); 
---Purpose: Hash on the Handle
class HashExtendedString;
---Purpose: Hash on the string.

end PColStd;


