-- Created on: 2001-07-25
-- Created by: Julia DOROVSKIKH
-- Copyright (c) 2001-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package XmlDrivers

uses
    Standard,
    TDF,
    TDocStd,
    TCollection,
    TColStd,
    CDM,
    PCDM,
    XmlObjMgt,
    XmlMDF,
    XmlLDrivers

is
    class DocumentStorageDriver;
    class DocumentRetrievalDriver;

    Factory (theGUID : GUID from Standard) returns Transient from Standard;

    AttributeDrivers (theMsgDriver: MessageDriver from CDM)
        returns ADriverTable from XmlMDF;

end XmlDrivers;
