-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Person from StepBasic 

inherits TShared from MMgt

uses

	HAsciiString from TCollection, 
	HArray1OfHAsciiString from Interface, 
	Boolean from Standard
is

	Create returns Person;
	---Purpose: Returns a Person

	Init (me : mutable;
	      aId : HAsciiString from TCollection;
	      hasAlastName : Boolean from Standard;
	      aLastName : HAsciiString from TCollection;
	      hasAfirstName : Boolean from Standard;
	      aFirstName : HAsciiString from TCollection;
	      hasAmiddleNames : Boolean from Standard;
	      aMiddleNames : HArray1OfHAsciiString from Interface;
	      hasAprefixTitles : Boolean from Standard;
	      aPrefixTitles : HArray1OfHAsciiString from Interface;
	      hasAsuffixTitles : Boolean from Standard;
	      aSuffixTitles : HArray1OfHAsciiString from Interface) is virtual;

	-- Specific Methods for Field Data Access --

	SetId(me : mutable; aId : HAsciiString);
	Id (me) returns HAsciiString;
	SetLastName(me : mutable; aLastName : HAsciiString);
	UnSetLastName (me:mutable);
	LastName (me) returns HAsciiString;
	HasLastName (me) returns Boolean;
	SetFirstName(me : mutable; aFirstName : HAsciiString);
	UnSetFirstName (me:mutable);
	FirstName (me) returns HAsciiString;
	HasFirstName (me) returns Boolean;
	SetMiddleNames(me : mutable; aMiddleNames : HArray1OfHAsciiString);
	UnSetMiddleNames (me:mutable);
	MiddleNames (me) returns HArray1OfHAsciiString;
	HasMiddleNames (me) returns Boolean;
	MiddleNamesValue (me; num : Integer) returns HAsciiString;
	NbMiddleNames (me) returns Integer;
	SetPrefixTitles(me : mutable; aPrefixTitles : HArray1OfHAsciiString);
	UnSetPrefixTitles (me:mutable);
	PrefixTitles (me) returns HArray1OfHAsciiString;
	HasPrefixTitles (me) returns Boolean;
	PrefixTitlesValue (me; num : Integer) returns HAsciiString;
	NbPrefixTitles (me) returns Integer;
	SetSuffixTitles(me : mutable; aSuffixTitles : HArray1OfHAsciiString);
	UnSetSuffixTitles (me:mutable);
	SuffixTitles (me) returns HArray1OfHAsciiString;
	HasSuffixTitles (me) returns Boolean;
	SuffixTitlesValue (me; num : Integer) returns HAsciiString;
	NbSuffixTitles (me) returns Integer;

fields

	id : HAsciiString from TCollection;
	lastName : HAsciiString from TCollection;   -- OPTIONAL can be NULL
	firstName : HAsciiString from TCollection;   -- OPTIONAL can be NULL
	middleNames : HArray1OfHAsciiString from Interface;   -- OPTIONAL can be NULL
	prefixTitles : HArray1OfHAsciiString from Interface;   -- OPTIONAL can be NULL
	suffixTitles : HArray1OfHAsciiString from Interface;   -- OPTIONAL can be NULL
	hasLastName : Boolean from Standard;
	hasFirstName : Boolean from Standard;
	hasMiddleNames : Boolean from Standard;
	hasPrefixTitles : Boolean from Standard;
	hasSuffixTitles : Boolean from Standard;

end Person;
