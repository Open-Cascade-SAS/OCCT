-- Created on: 1993-01-11
-- Created by: CKY / Contract Toubro-Larsen ( Anand NATRAJAN )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class LevelToPWBLayerMap from IGESAppli  inherits IGESEntity

        ---Purpose: defines LevelToPWBLayerMap, Type <406> Form <24>
        --          in package IGESAppli
        --          Used to correlate an exchange file level number with
        --          its corresponding native level identifier, physical PWB
        --          layer number and predefined functional level
        --          identification

uses

        HAsciiString           from TCollection,
        HArray1OfInteger       from TColStd,
        HArray1OfHAsciiString  from Interface

raises DimensionMismatch, OutOfRange

is

        Create returns mutable LevelToPWBLayerMap;

        -- Specific Methods pertaining to the class

        Init (me              : mutable;
              nbPropVal       : Integer;
              allExchLevels   : HArray1OfInteger;
              allNativeLevels : HArray1OfHAsciiString;
              allPhysLevels   : HArray1OfInteger;
              allExchIdents   : HArray1OfHAsciiString)
        raises DimensionMismatch;
        ---Purpose : This method is used to set the fields of the class
        --           LevelToPWBLayerMap
        --       - nbPropVal       : Number of property values
        --       - allExchLevels   : Exchange File Level Numbers
        --       - allNativeLevels : Native Level Identifications
        --       - allPhysLevels   : Physical Layer Numbers
        --       - allExchIdents   : Exchange File Level Identifications
        -- raises exception if allExchLevels, allNativeLevels, allPhysLevels
        -- and all ExchIdents are not of same dimensions

        NbPropertyValues (me) returns Integer;
        ---Purpose : returns number of property values

        NbLevelToLayerDefs (me) returns Integer;
        ---Purpose : returns number of level to layer definitions

        ExchangeFileLevelNumber (me; Index : Integer) returns Integer
        raises OutOfRange;
        ---Purpose : returns Exchange File Level Number
        -- raises exception if Index <= 0 or Index > NbLevelToLayerDefs

        NativeLevel (me; Index : Integer) returns HAsciiString from TCollection
        raises OutOfRange;
        ---Purpose : returns Native Level Identification
        -- raises exception if Index <= 0 or Index > NbLevelToLayerDefs

        PhysicalLayerNumber (me; Index : Integer) returns Integer
        raises OutOfRange;
        ---Purpose : returns Physical Layer Number
        -- raises exception if Index <= 0 or Index > NbLevelToLayerDefs

        ExchangeFileLevelIdent (me; Index : Integer)
                    returns HAsciiString from TCollection
        raises OutOfRange;
        -- returns Exchange File Level Identification
        -- raises exception if Index <= 0 or Index > NbLevelToLayerDefs

fields

--
-- Class    : IGESAppli_LevelToPWBLayerMap
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class LevelToPWBLayerMap.
--
-- Reminder : A LevelToPWBLayerMap instance is defined by :
--            - Number of property values
--            - Exchange File Level Numbers
--            - Native Level Identifications
--            - Physical Layer Numbers
--            - Exchange File Level Identifications

        theNbPropertyValues        : Integer;
        theExchangeFileLevelNumber : HArray1OfInteger;
        theNativeLevel             : HArray1OfHAsciiString;
        thePhysicalLayerNumber     : HArray1OfInteger;
        theExchangeFileLevelIdent  : HArray1OfHAsciiString;

end LevelToPWBLayerMap;
