-- File:	StepVisual_DraughtingModel.cdl
-- Created:	Thu Jan 13 10:08:42 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0
-- Copyright:	Matra Datavision 1999

class DraughtingModel from StepVisual
inherits Representation from StepRepr

    ---Purpose: Representation of STEP entity DraughtingModel

uses
    HAsciiString from TCollection,
    HArray1OfRepresentationItem from StepRepr,
    RepresentationContext from StepRepr

is
    Create returns DraughtingModel from StepVisual;
	---Purpose: Empty constructor

end DraughtingModel;
