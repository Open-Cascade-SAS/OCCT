-- Created on: 1997-10-02
-- Created by: Denis PASCAL
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package DPrsStd 

        ---Purpose:  commands for presentation based on AIS
        --           ======================================


uses Draw


is    

    ---Purpose: Presentation commands
    --          =====================

    AllCommands (I : in out Interpretor from Draw);
    ---Purpose: to load all sketch commands   


    AISPresentationCommands (I : in out Interpretor from Draw);
    ---Purpose: to display....etc... ais presentation

    AISViewerCommands (I : in out Interpretor from Draw);
    ---Purpose: to repaint...etc... ais viewer

    BasicCommands (I : in out Interpretor from Draw);
    ---Purpose: set/get position attribute

    Factory (theDI : out Interpretor from Draw);
    ---Purpose: Loads all Draw commands of  TKDCAF. Used for plugin. 
    
end DPrsStd;




