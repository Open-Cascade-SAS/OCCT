-- Created on: 1997-03-26
-- Created by: Christian CAILLET
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class AutoDesignPresentedItemSelect from StepAP214 inherits SelectType from StepData

	-- <AutoDesignPresentedItemSelect> is an EXPRESS Select Type construct translation.
	-- it gathers : ProductDefinition, ProductDefinitionShape, RepresentationRelationship, ShapeAspect

uses
     ProductDefinition from StepBasic,
     ProductDefinitionRelationship from StepBasic,
     ProductDefinitionShape from StepRepr,
     RepresentationRelationship from StepRepr,
     ShapeAspect from StepRepr,
     DocumentRelationship from StepBasic

is

	Create returns AutoDesignPresentedItemSelect;
	---Purpose : Returns a AutoDesignPresentedItemSelect SelectType

	CaseNum (me; ent : Transient) returns Integer;
	---Purpose: Recognizes a AutoDesignPresentedItemSelect Kind Entity that is :
	--  1 -> ProductDefinition,
	--  2 -> ProductDefinitionRelationship,
	--  3 -> ProductDefinitionShape
	--  4 -> RepresentationRelationship
	--  5 -> ShapeAspect
	--  6 -> DocumentRelationship,
	--        0 else

    ProductDefinitionRelationship (me) returns any ProductDefinitionRelationship;
    ---Purpose : returns Value as a ProductDefinitionRelationship (Null if another type)

    ProductDefinition (me) returns any ProductDefinition;
    ---Purpose : returns Value as a ProductDefinition (Null if another type)

    ProductDefinitionShape (me) returns any ProductDefinitionShape;
    ---Purpose : returns Value as a ProductDefinitionShape (Null if another type)

    RepresentationRelationship (me) returns any RepresentationRelationship;
    ---Purpose : returns Value as a RepresentationRelationship (Null if another type)

    ShapeAspect (me) returns any ShapeAspect;
    ---Purpose : returns Value as a ShapeAspect (Null if another type)

    DocumentRelationship (me) returns any DocumentRelationship;
    ---Purpose : returns Value as a DocumentRelationship (Null if another type)

end AutoDesignPresentedItemSelect;
