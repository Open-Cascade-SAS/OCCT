-- File:	RWStepDimTol_RWGeometricTolerance.cdl
-- Created:	Wed Jun  4 13:34:35 2003 
-- Author:	Galina KULIKOVA
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWGeometricTolerance from RWStepDimTol

    ---Purpose: Read & Write tool for GeometricTolerance

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    GeometricTolerance from StepDimTol

is
    Create returns RWGeometricTolerance from RWStepDimTol;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : GeometricTolerance from StepDimTol);
	---Purpose: Reads GeometricTolerance

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: GeometricTolerance from StepDimTol);
	---Purpose: Writes GeometricTolerance

    Share (me; ent : GeometricTolerance from StepDimTol;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWGeometricTolerance;
