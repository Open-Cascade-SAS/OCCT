-- Created on: 1991-09-02
-- Created by: Mireille MERCIEN
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

generic class HStack from PCollection (Item as Storable) 
inherits Persistent

    ---Purpose: A stack is a list of items in which items are
    -- added and removed from the same end, called the 
    -- top of the stack.

raises   NoSuchObject from Standard


    class StackNode instantiates HSingleList from PCollection(Item);

    class StackIterator from PCollection 
    	    	    	    	    	   
        ---Purpose: Iterator of the Stack class.

    raises NoMoreObject from Standard,
           NoSuchObject from Standard
    is     
 
     	Create(S : HStack from PCollection) 
    	returns StackIterator from PCollection;
        ---Purpose: Creates an iterator on the stack S.
        -- Set the iterator at the beginning of the stack S.

     	More(me) returns Boolean from Standard;
        ---Level: Public
        ---Purpose: Returns True if there are other items.

     	Next(me: in out) raises NoMoreObject from Standard;
        ---Level: Public
	---Purpose: Sets the iterator to the next item.
	    
	Value(me) returns any Item raises NoSuchObject from Standard;
        ---Level: Public
	---Purpose: Returns the item value corresponding to 
	-- the current position of the iterator.

    fields
    	 TheIterator : StackNode;
    end;


is
     Create returns mutable HStack from PCollection;
       ---Purpose: Creates an empty stack.

     Depth(me) returns Integer from Standard;
       ---Level: Public
       ---Purpose: Returns the number of items in the stack.
       ---Example: if me = (A B C) 
       -- returns 3

     IsEmpty(me) returns Boolean from Standard;
       ---Level: Public
       ---Purpose: Returns True if the stack contains no item.

     Top(me) returns any Item 
       ---Level: Public
       ---Purpose: Returns the item on the top of the stack.
       -- Raises an exception if the stack is empty.
       ---Example: before
       --   me = (A B C) 
       -- after
       --   me = (A B C)
       -- returns 
       --   C
      raises NoSuchObject from Standard;

     FTop(me) returns StackNode; 
       ---Level: Public
       ---Purpose: Returns the field TheTop (the top of the stack).

     Push(me : mutable; T : Item);
       ---Level: Public
       ---Purpose: Inserts an item on the top of the stack.
       ---Example: before
       --   me = (A B) , T = C
       -- after
       --   me = (A B C)

     Pop(me : mutable) raises NoSuchObject from Standard;
       ---Level: Public
       ---Purpose: Removes an item from the top of the stack.
       -- Raises an exception if the stack is empty.
       ---Example: before
       --   me = (A B C) 
       -- after    
       --   me = (A B)
       -- returns
       --   C

     Clear(me : mutable);
       ---Level: Public
       ---Purpose: Removes all the items from the stack.
       ---Example: before
       --   me = (A B C) 
       -- after
       --   me = ()
 
     ChangeTop(me:mutable; T : Item) raises NoSuchObject from Standard;
       ---Level: Public
       ---Purpose: Replaces the top of the stack with T.
       -- Raises an exception if the stack is empty.
       ---Example: before
       --   me = (A B C) , T = D
       -- after
       --   me = (A B D)


     ShallowCopy(me) 
        returns mutable like me 
        is redefined;
        ---Level: Advanced
	---C++: function call


     ShallowDump (me; s: in out OStream) 
        is redefined;
        ---Level: Advanced
    	---C++: function call



fields
     TheTop   : StackNode;
     TheDepth : Integer from Standard;
     
end; 






