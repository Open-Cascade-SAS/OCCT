-- Created on: 1996-09-10
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DrawableSUR from TestTopOpeDraw inherits Surface from DrawTrSurf

uses 
    
    Surface     from Geom,
    Color           from Draw,
    Display         from Draw,
    Text3D          from Draw,
    CString         from Standard,
    Pnt             from gp,
    Pnt2d           from gp

is 

    Create (S : Surface from Geom; IsoColor : Color from Draw)
    returns mutable DrawableSUR from TestTopOpeDraw;

    Create (S : Surface from Geom; IsoColor : Color from Draw;
    	    Text : CString from Standard; TextColor : Color from Draw)
    returns mutable DrawableSUR from TestTopOpeDraw;

    Create (S : Surface from Geom; IsoColor : Color from Draw;
            BoundColor,NormalColor : Color from Draw;
    	    Text : CString from Standard; TextColor : Color from Draw;
	    Nu,Nv : Integer;
    	    Discret : Integer; Deflection : Real; DrawMode : Integer;
    	    DispOrigin : Boolean from Standard = Standard_True)
    returns mutable DrawableSUR from TestTopOpeDraw;

    Pnt(me) returns Pnt from gp
    is static;

    Pnt2d(me) returns Pnt2d from gp
    is static;
    
    DrawOn(me; dis : in out Display from Draw)
    is redefined;

    NormalColor(me : mutable; NormalColor : Color from Draw)
    is static;

    DrawNormale(me; dis : in out Display from Draw)
    is static;
    
fields

    myText : Text3D from Draw;
    myNormalColor : Color from Draw;
    
end DrawableSUR;
