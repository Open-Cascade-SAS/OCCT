-- Created on: 2002-01-04
-- Created by: data exchange team
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1

class Subedge from StepShape
inherits Edge from StepShape

    ---Purpose: Representation of STEP entity Subedge

uses
    HAsciiString from TCollection,
    Vertex from StepShape,
    Edge from StepShape

is
    Create returns Subedge from StepShape;
	---Purpose: Empty constructor

    Init (me: mutable; aRepresentationItem_Name: HAsciiString from TCollection;
                       aEdge_EdgeStart: Vertex from StepShape;
                       aEdge_EdgeEnd: Vertex from StepShape;
                       aParentEdge: Edge from StepShape);
	---Purpose: Initialize all fields (own and inherited)

    ParentEdge (me) returns Edge from StepShape;
	---Purpose: Returns field ParentEdge
    SetParentEdge (me: mutable; ParentEdge: Edge from StepShape);
	---Purpose: Set field ParentEdge

fields
    theParentEdge: Edge from StepShape;

end Subedge;
