-- Created on: 1999-11-26
-- Created by: Andrey BETENEV
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0

class CcDesignSecurityClassification from StepAP203
inherits SecurityClassificationAssignment from StepBasic

    ---Purpose: Representation of STEP entity CcDesignSecurityClassification

uses
    SecurityClassification from StepBasic,
    HArray1OfClassifiedItem from StepAP203

is
    Create returns CcDesignSecurityClassification from StepAP203;
	---Purpose: Empty constructor

    Init (me: mutable; aSecurityClassificationAssignment_AssignedSecurityClassification: SecurityClassification from StepBasic;
                       aItems: HArray1OfClassifiedItem from StepAP203);
	---Purpose: Initialize all fields (own and inherited)

    Items (me) returns HArray1OfClassifiedItem from StepAP203;
	---Purpose: Returns field Items
    SetItems (me: mutable; Items: HArray1OfClassifiedItem from StepAP203);
	---Purpose: Set field Items

fields
    theItems: HArray1OfClassifiedItem from StepAP203;

end CcDesignSecurityClassification;
