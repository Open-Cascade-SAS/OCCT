-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class SolidClassifier from BOP

    ---Purpose: 
    --  The  auxiliary class to classify points with 
    --  a solid  
    --	     
uses 

    State from TopAbs,
    Shell from TopoDS,
    Solid from TopoDS,
    Pnt   from gp,
    PSoClassif                      from BOP,
    IndexedDataMapOfSolidClassifier from BOP,
    Builder from BRep
    
is

    Create  
    	returns SolidClassifier from BOP;
    	---Purpose:  
    	--- Empty  Constructor 
    	---
    Clear(me:out)  
    	is static;
    	---Purpose:  
    	--- Clear internal state  
    	---
    LoadSolid(me: out;  
    	    aS : Solid from TopoDS)  
    	is static;
    	---Purpose:  
    	--- Modifier  
    	---
    Classify(me:out;  
    	    aS : Solid from TopoDS;  
    	    aP : Pnt from gp;  
    	    aTol: Real from Standard) 
    returns State from TopAbs
    	is static;
    	---Purpose:  
    	--- Compute the position of point <P> regarding with the
    	--- geometric domain of the solid <S>.  
    	---
    	

    LoadShell(me:out;  
    	    S : Shell from TopoDS) 
    	 is static;
    	---Purpose:  
    	--- Modifier  
    	---
    Classify(me:out;  
    	    aS : Shell from TopoDS;  
    	    aP : Pnt from gp;  
    	    aTol : Real  from  Standard) 
    returns State from TopAbs
    	is static;
    	---Purpose:  
    	--- Compute the position of point <P> regarding with the
    	--- geometric domain of the shell <S>. 
	---
    State(me)  
    	returns State from TopAbs
    	is static;   
    	---Purpose: 
    	--- Returns computed 3D-State   
    	---
    Destroy (me:out); 
    	---C++: alias "Standard_EXPORT virtual ~BOP_SolidClassifier(){Destroy();}"  
    	---Purpose: 
    	--- Destructor   
    	---
    
fields

    myPClassifier   : PSoClassif from BOP;  
    myClassifierMap : IndexedDataMapOfSolidClassifier from BOP;
    myState         : State from TopAbs;    
    myShell         : Shell from TopoDS;
    mySolid         : Solid from TopoDS;
    myBuilder       : Builder from BRep;
    
end SolidClassifier from BOP;
