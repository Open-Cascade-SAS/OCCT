-- Created on: 1993-04-06
-- Created by: Philippe DAUTRY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class AxisPlacement from PGeom2d inherits Geometry from PGeom2d

        ---Purpose :   An  axis  placement  defines a  local cartesian
        --         coordinate  system and   can be used to  locate  an
        --         entity in 3D space.
        --  

uses Ax2d from gp

is


    Create returns mutable AxisPlacement from PGeom2d;
	---Purpose: Initializes the field(s) with default value(s).
	---Level: Internal 


    Create(aAxis: Ax2d from gp) returns mutable AxisPlacement from PGeom2d;
	---Purpose: Initializes the field axis with <aAxis>.
	---Level: Internal 


  Axis (me : mutable; aAxis : Ax2d from gp);
        --- Purpose : Set the field axis with <aAxis>.
	---Level: Internal 


  Axis (me)  returns Ax2d from gp;
        --- Purpose : Returns the value of the field axis.
	---Level: Internal 


fields

  axis : Ax2d from gp;

end;
