-- Created on: 1998-07-29
-- Created by: Christian CAILLET
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package STEPEdit

    ---Purpose : Provides tools to exploit and edit a set of STEP data :
    --           editors, selections ..

uses Standard, TCollection,
     Interface, IFSelect, StepData

is

    class EditContext;
    -- This class is for global context : ApplicationContext,
    --   ProductRelatedProductCategory

    class EditSDR;
    -- This class allows to edit product data for a SDR


    	--  Some useful operators
    	--  They are not classes, they are just based on general tools

    Protocol returns Protocol from Interface;
    ---Purpose : Returns a Protocol fit for STEP (creates the first time)

    NewModel returns StepModel from StepData;
    ---Purpose : Returns a new empty StepModel fit for STEP
    --           i.e. with its header determined from Protocol

    SignType returns Signature from IFSelect;
    ---Purpose : Returns a SignType fit for STEP (creates the first time)

    NewSelectSDR returns SelectSignature from IFSelect;
    ---Purpose : Creates a Selection for ShapeDefinitionRepresentation
    --           By default searches among root entities

    NewSelectPlacedItem returns SelectSignature from IFSelect;
    ---Purpose : Creates a Selection for Placed Items, i.e. MappedItem or
    --           ContextDependentShapeRepresentation, which itself refers to a
    --           RepresentationRelationship with possible subtypes (Shape...
    --           and/or ...WithTransformation)
    --           By default in the whole StepModel

    NewSelectShapeRepr returns SelectSignature from IFSelect;
    ---Purpose : Creates a Selection for ShapeRepresentation and its sub-types,
    --           plus ContextDependentShapeRepresentation (which is not a
    --           sub-type of ShapeRepresentation)
    --           By default in the whole StepModel

end STEPEdit;
