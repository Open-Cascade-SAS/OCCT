-- File:	QAMitutoyoUK.cdl
-- Created:	Tue Mar 19 12:16:49 2002
-- Author:	QA Admin
--		<qa@umnox.nnov.matra-dtv.fr>
---Copyright:	 Matra Datavision 2002

package QAMitutoyoUK
     uses Draw
is
    Commands(DI : in out Interpretor from Draw);
end;
