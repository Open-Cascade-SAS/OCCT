-- File:	Interface_IntVal.cdl
-- Created:	Wed Sep  3 15:25:38 1997
-- Author:	Christian CAILLET
--		<cky@heliox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1997


class IntVal  from Interface    inherits TShared  from MMgt

    ---Purpose : An Integer through a Handle (i.e. managed as TShared)

uses Integer

is

    Create returns mutable IntVal;

    Value (me) returns Integer;

    CValue (me : mutable) returns Integer;
    ---C++ : return &

fields

    theval : Integer;

end IntVal;
