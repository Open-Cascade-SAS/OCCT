-- Created on: 1995-10-23
-- Created by: Mister rmi
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PolygonOnTriangulation from PBRep inherits CurveRepresentation from PBRep


    	---Purpose: A representation by an array of nodes on a 
    	--          triangulation.


uses Location               from PTopLoc,
     PolygonOnTriangulation from PPoly,
     Triangulation          from PPoly

is

    Create(P: PolygonOnTriangulation from PPoly;
    	   T: Triangulation          from PPoly;
	   L: Location               from PTopLoc)
    returns mutable PolygonOnTriangulation from PBRep;
    
    
    IsPolygonOnTriangulation(me) returns Boolean
    	---Purpose: returns True.
    is redefined;

    PolygonOnTriangulation(me) returns any PolygonOnTriangulation from PPoly;

    Triangulation(me) returns any Triangulation from PPoly;
        
fields

    myPolygon       : PolygonOnTriangulation from PPoly;
    myTriangulation : Triangulation          from PPoly;

end PolygonOnTriangulation;
