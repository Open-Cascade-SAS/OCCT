-- Created on: 1993-02-22
-- Created by: Philippe DAUTRY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class Transformation from PGeom inherits Persistent from Standard

        ---Purpose :  The    class Transformation  allows   to  create
        --         Translation, Rotation,   Symmetry,     Scaling  and
        --         complex transformations obtained by  combination of
        --         the  previous elementary   transformations.     The
        --         restriction to  these basic  transformations allows
        --         us to be sure that   an object  will never   change
        --         nature.
        --         
	---See Also : Transformation from Geom.


uses Trsf from gp

is


  Create returns mutable Transformation from PGeom;
        ---Purpose : Creates a transformation with default values.
    	---Level: Internal 


  Create (aTrsf : Trsf from gp) returns mutable Transformation from PGeom;
        ---Purpose :  Creates a transformation with <aTrsf>.
    	---Level: Internal 


  Trsf (me : mutable; aTrsf : Trsf from gp);
        ---Purpose : Set the field trsf with <aTrsf>.
    	---Level: Internal 


  Trsf (me)  returns Trsf from gp;
        ---Purpose : Returns the value of the field trsf.
    	---Level: Internal 


fields

  trsf : Trsf from gp;

end;
