-- Created on: 1997-07-28
-- Created by: Pierre CHALAMET
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class  Texture1Dmanual  from  Graphic3d 

inherits  Texture1D  from  Graphic3d  
 
---Purpose: This class provides the implementation of
-- a manual 1D texture.
-- you MUST provides texture coordinates on
-- your facets if you want to see your
-- texture. 


uses 
    NameOfTexture1D  from  Graphic3d, 
    StructureManager    from  Graphic3d

is 
    Create(SM  :  StructureManager  from  Graphic3d; 
           FileName  :  CString  from  Standard)  returns  mutable  Texture1Dmanual  from  Graphic3d; 
    ---Purpose: Creates a texture from the file FileName.


    Create(SM  :  StructureManager  from  Graphic3d; 
    	   NOT  :  NameOfTexture1D  from  Graphic3d)  returns  mutable  Texture1Dmanual  from  Graphic3d;
    ---Purpose: Create a texture from a predefined texture name set.

end  Texture1Dmanual; 

