-- Created on: 1994-12-21
-- Created by: Christian CAILLET
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class IGESName from IGESSelect    inherits Signature  from IFSelect

    ---Purpose : IGESName is a Signature specific to IGESNorm :
    --           it considers the Name of an IGESEntity as being its ShortLabel
    --           (some sending systems use name, not to identify entities, but
    --           ratjer to classify them)

uses CString, Transient, InterfaceModel

is

    Create returns IGESName;
    ---Purpose : Creates a Signature for IGES Name (reduced to ShortLabel,
    --           without SubscriptLabel or Long Name)

    Value (me; ent : any Transient; model : InterfaceModel) returns CString;
    ---Purpose : Returns the ShortLabel as being the Name of an IGESEntity
    --           If <ent> has no name, it returns empty string ""

end IGESName;
