-- Created on: 2000-02-14
-- Created by: Denis PASCAL
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class CopyShape from TNaming 

	---Purpose: 

uses Shape from TopoDS,
     IndexedDataMapOfTransientTransient from TColStd,
     TranslateTool from TNaming,
     Location from TopLoc

is

    CopyTool (myclass;
              aShape    :  Shape      from TopoDS;
    	      aMap      :  in out  IndexedDataMapOfTransientTransient from TColStd; 
	      aResult   :  in  out Shape  from  TopoDS);
	---Purpose:      Makes  copy  a  set  of  shape(s),  using the  aMap 
	 
	  
    Translate (myclass;
               aShape  : Shape          from TopoDS; 
	       aMap    : in out  IndexedDataMapOfTransientTransient from TColStd; 
	       aResult : in  out Shape  from  TopoDS;
    	       TrTool  : TranslateTool  from TNaming); 
	     
	 ---Purpose: Translates  a  Transient  shape(s)  to  Transient     
	    
    Translate (myclass;
               L : Location from TopLoc; 
     	       aMap :  in out  IndexedDataMapOfTransientTransient from TColStd)   	       
    returns Location from TopLoc; 
     ---Purpose: Translates a Topological  Location  to an  other  Top.
     --          Location 

end CopyShape;
