-- Created on: 1992-02-07
-- Created by: Laurent PAINNOT
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DoubleTab from math
uses Address from Standard
is

    Create(LowerRow, UpperRow, LowerCol, UpperCol: Integer)
    	returns DoubleTab;

    Create(Tab : Address; LowerRow, UpperRow, LowerCol, UpperCol: Integer)
    	returns DoubleTab;

    Init(me : in out; InitValue: Real) is static;

    Create(Other: DoubleTab)
    	returns DoubleTab;

    Allocate(me : in out) is private;
    
    Copy(me; Other: in out DoubleTab)
    	---C++: inline
    is static;

    
    SetLowerRow(me: in out; LowerRow: Integer)
    is static;


    SetLowerCol(me: in out; LowerCol: Integer)
    is static;

        
    Value(me; RowIndex, ColIndex: Integer)
    	---C++: alias operator()
    	---C++: return &
    	---C++: inline
      returns Real
      is static;		
	
	
    Free(me: in out)
        ---C++: alias ~

    is static;
    
    
fields

Addr        : Address;
AddrBuf     : Address[32];
Buf         : Real[512];
isAddrAllocated: Boolean;
isAllocated : Boolean;
LowR        : Integer;
UppR        : Integer;
LowC        : Integer;
UppC        : Integer;

end DoubleTab;	
