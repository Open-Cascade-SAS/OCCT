-- Created on: 1994-06-01
-- Created by: Modelistation
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SetGlobalParameter  from IGESSelect  inherits ModelModifier from IGESSelect

    ---Purpose : Sets a Global (Header) Parameter to a new value, directly given
    --           Controls the form of the parameter (Integer, Real, String
    --           with such or such form), but not the consistence of the new
    --           value regarding the rest of the file.
    --           
    --           The new value is given under the form of a HAsciiString, even
    --           for Integer or Real values. For String values, Hollerith forms
    --           are accepted but not mandatory
    --  Warning : a Null (not set) value is not accepted. For an empty string,
    --           give a Text Parameter which is empty

uses AsciiString from TCollection, HAsciiString from TCollection,
     IGESModel, CopyTool, ContextModif

is

    Create (numpar : Integer) returns mutable SetGlobalParameter;
    ---Purpose : Creates an SetGlobalParameter, to be applied on Global
    --           Parameter <numpar>

    GlobalNumber (me) returns Integer;
    ---Purpose : Returns the global parameter number to which this modifiers
    --           applies

    SetValue (me : mutable; text : mutable HAsciiString);
    ---Purpose : Sets a Text Parameter for the new value

    Value (me) returns mutable HAsciiString;
    ---Purpose : Returns the value to set to the global parameter (Text Param)


    Performing (me; ctx : in out ContextModif;
    	        target  : mutable IGESModel;
                TC      : in out CopyTool);
    ---Purpose : Specific action : only <target> is used : the form of the new
    --           value is checked regarding the parameter number (given at
    --           creation time).

    Label (me) returns AsciiString from TCollection;
    ---Purpose : Returns a text which is
    --           "Sets Global Parameter <numpar> to <new value>"

fields

    thenum : Integer;
    theval : HAsciiString from TCollection;

end SetGlobalParameter;
