-- File:	IntPatch_PolygoTool.cdl
-- Created:	Thu May  6 17:50:02 1993
-- Author:	Jacques GOUSSARD
--		<jag@form4>
---Copyright:	 Matra Datavision 1993


 
class PolygoTool from IntPatch

       	---Purpose: Tool an a polygon to instantiates the Interference
       	--          between 2 polygons.


uses Box2d  from Bnd,
     Pnt2d  from gp,
     Polygo from IntPatch
 

is

    Bounding (myclass; Line : Polygo from IntPatch )

    	returns Box2d from Bnd;
        ---C++: return const &
	---C++: inline


    DeflectionOverEstimation(myclass; Line :Polygo from IntPatch)

    	returns Real from Standard;
	---C++: inline
                         	    	          

    Closed(myclass; Line : Polygo from IntPatch )

    	returns Boolean from Standard;
	---C++: inline


    NbSegments(myclass; Line : Polygo from IntPatch )

    	returns Integer from Standard;
	---C++: inline


    BeginOfSeg(myclass; Line  : Polygo from IntPatch;
                        Index : Integer from Standard)

    	returns Pnt2d from gp;
	---C++: inline


    EndOfSeg(myclass; Line  : Polygo from IntPatch ;
                      Index : Integer from Standard)

    	returns Pnt2d from gp;
	---C++: inline


    Dump(myclass; Line  : Polygo from IntPatch);
    

end PolygoTool;
		 
