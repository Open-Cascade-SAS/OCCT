-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class OrientedPath from StepShape 

inherits Path from StepShape 

uses

	Boolean from Standard, 
	HArray1OfOrientedEdge from StepShape, 
	OrientedEdge from StepShape, 
	HAsciiString from TCollection,
	EdgeLoop from StepShape
is

	Create returns mutable OrientedPath;
	---Purpose: Returns a OrientedPath


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aEdgeList : mutable HArray1OfOrientedEdge from StepShape) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aPathElement : mutable EdgeLoop from StepShape;
	      aOrientation : Boolean from Standard) is virtual;

	-- Specific Methods for Field Data Access --

	SetPathElement(me : mutable; aPathElement : mutable EdgeLoop);
	PathElement (me) returns mutable EdgeLoop;
	SetOrientation(me : mutable; aOrientation : Boolean);
	Orientation (me) returns Boolean;
	SetEdgeList(me : mutable; aEdgeList : mutable HArray1OfOrientedEdge) is redefined;
	EdgeList (me) returns mutable HArray1OfOrientedEdge is redefined;
	EdgeListValue (me; num : Integer) returns mutable OrientedEdge is redefined;
	NbEdgeList (me) returns Integer is redefined;

fields

	pathElement : EdgeLoop from StepShape;
	orientation : Boolean from Standard;

 -- 
 -- NB : field <edge_list> inherited from classe <EdgeLoop> is redeclared.
 --      it shall appears in a physical file as a *.
 --

end OrientedPath;
