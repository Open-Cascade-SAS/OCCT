-- Created on: 1992-09-30
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class QuadricTool from IntSurf

	---Purpose: This class provides a tool on a quadric that can be
	--          used to instantiates the Walking algorithmes (see
	--          package IntWalk) with a Quadric from IntSurf
	--          as implicit surface.

uses Quadric from IntSurf,
     Vec     from gp

is

    Value(myclass; Quad: Quadric from IntSurf;
          X, Y, Z: Real from Standard)
	  
    	---Purpose: Returns the value of the function.
    
    	returns Real from Standard;
	
	---C++: inline
    
    
    Gradient(myclass; Quad: Quadric from IntSurf;
             X, Y, Z: Real from Standard ; V : out Vec from gp);
	     
    	---Purpose: Returns the gradient of the function.

	---C++: inline
    


    ValueAndGradient(myclass; Quad: Quadric from IntSurf;
                     X, Y, Z: Real from Standard;
                     Val: out Real from Standard; Grad: out Vec from gp);
		     
    	---Purpose: Returns the value and the gradient.

	---C++: inline
    

    Tolerance(myclass; Quad: Quadric from IntSurf )
    
	---Purpose: returns the tolerance of the zero of the implicit function

    	returns Real from Standard; 


end QuadricTool;


