-- Created on: 2001-12-28
-- Created by: Andrey BETENEV
-- Copyright (c) 2001-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1

class EdgeBasedWireframeModel from StepShape
inherits GeometricRepresentationItem from StepGeom

    ---Purpose: Representation of STEP entity EdgeBasedWireframeModel

uses
    HAsciiString from TCollection,
    HArray1OfConnectedEdgeSet from StepShape

is
    Create returns EdgeBasedWireframeModel from StepShape;
	---Purpose: Empty constructor

    Init (me: mutable; aRepresentationItem_Name: HAsciiString from TCollection;
                       aEbwmBoundary: HArray1OfConnectedEdgeSet from StepShape);
	---Purpose: Initialize all fields (own and inherited)

    EbwmBoundary (me) returns HArray1OfConnectedEdgeSet from StepShape;
	---Purpose: Returns field EbwmBoundary
    SetEbwmBoundary (me: mutable; EbwmBoundary: HArray1OfConnectedEdgeSet from StepShape);
	---Purpose: Set field EbwmBoundary

fields
    theEbwmBoundary: HArray1OfConnectedEdgeSet from StepShape;

end EdgeBasedWireframeModel;
