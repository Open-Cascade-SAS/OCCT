-- Created on: 1991-05-27
-- Created by: Laurent PAINNOT
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class IntegerRandom from math
   ---Purpose:
   -- This class implements an integer random number generator.

is

   Create(Lower, Upper: Integer)
   ---Purpose:
   -- creates a Integer random generator between the values Lower and Upper.
    
   returns IntegerRandom;
   
    
   Reset(me:in out)
    	---Purpose: reinitializes the random generator

   is static;

   Next(me: in out)
    ---Purpose: returns the next random number.

   returns Integer
   is static;
   
fields

Low:    Integer;
Up:     Integer;
Dummy:  Integer;

end IntegerRandom;
