-- Created on: 1998-11-25
-- Created by: Denis PASCAL
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PlanarDiameter from DrawDim inherits PlanarDimension from DrawDim

	---Purpose: 

uses Vertex  from TopoDS,
     Face    from TopoDS,
     Shape   from TopoDS,
     Color   from Draw,
     Display from Draw

is

    Create (plane  : Face  from TopoDS;
            circle : Shape from TopoDS)
    returns PlanarDiameter from DrawDim;    

    Create (circle : Shape from TopoDS)
    returns PlanarDiameter from DrawDim;
    
    DrawOn(me; dis : in out Display);
    
fields

    myCircle : Shape   from TopoDS;

end PlanarDiameter;
