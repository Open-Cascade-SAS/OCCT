-- Created on: 1992-06-04
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




package Geom2dInt 

	---Purpose: Intersection between two Curves2 from Geom2dAdaptor

        ---Level: Public
        --
        -- All the methods of the classes are public.
        --


uses Standard, gp, TColStd, GeomAbs, Geom2d, Adaptor3d,Adaptor2d, IntCurve

is

   generic class CurveTool;

   class Geom2dCurveTool instantiates CurveTool from Geom2dInt
            (Curve2d      from Adaptor2d);
    	 
   class GInter instantiates IntCurveCurveGen from IntCurve
            (Curve2d         from Adaptor2d,
             Geom2dCurveTool from Geom2dInt);

end Geom2dInt; 
 
