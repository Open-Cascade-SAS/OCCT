-- Created on: 1992-04-03
-- Created by: Laurent BUCHARD
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package IntRes2d


    ---Purpose: This package provides the definition of the results of
    --          the intersection between 2D curves and the definition
    --          of a domain on a 2D curve.
    ---Level: Public 
    -- 
    -- All the methods of all the classes of this package are public.
    --

uses

    Standard, TCollection, gp, StdFail

is


    class IntersectionPoint;
    
    class IntersectionSegment;

    class Transition;

    class Domain;

    deferred class Intersection;

    enumeration Position is Head,Middle,End;

    enumeration TypeTrans is In,Out,Touch,Undecided;

    enumeration Situation is Inside, Outside, Unknown;

    class SequenceOfIntersectionPoint instantiates
    	       Sequence from TCollection (IntersectionPoint);

    class SequenceOfIntersectionSegment instantiates
    	       Sequence from TCollection (IntersectionSegment);


end IntRes2d; 


