-- Created on: 1992-09-28
-- Created by: Remi GILET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MakeHyperbola from GCE2d inherits Root from GCE2d

    ---Purpose :This class implements the following algorithms used to 
    --          create Hyperbola from Geom2d.
    --          * Create an Hyperbola from two apex  and the center.
    --  Defines the main branch of an hyperbola.
    --  The parameterization range is ]-infinite,+infinite[
    --  It is possible to get the other branch and the two conjugate
    --  branches of the main branch.
    --
    --                         ^YAxis                
    --                         |                   
    --                  FirstConjugateBranch     
    --                         |        
    --        Other            |                Main
    --   --------------------- C ------------------------------>XAxis
    --        Branch           |                Branch
    --                         |         
    --                   SecondConjugateBranch
    --                         |         
    --
    --  The major radius is the distance between the Location point
    --  of the hyperbola C and the apex of the main Branch (or the
    --  Other branch). The major axis is the "XAxis".
    --  The minor radius is the distance between the Location point
    --  of the hyperbola C and the apex of the First (or Second)
    --  Conjugate branch. The minor axis is the "YAxis".
    --  The major radius can be lower than the minor radius.

uses Pnt2d     from gp,
     Hypr      from gp,
     Hypr2d    from gp,
     Ax2d      from gp,
     Ax22d     from gp,
     Hyperbola from Geom2d

raises NotDone from StdFail

is

Create (H : Hypr2d from gp) returns MakeHyperbola;
    --- Purpose :
    --  Creates  an Hyperbola from a non persistent one from package gp

Create (MajorAxis   : Ax2d    from gp      ; 
    	MajorRadius : Real    from Standard;
    	MinorRadius : Real    from Standard;
    	Sense       : Boolean from Standard) returns MakeHyperbola;
    --- Purpose :
    --  MajorAxis is the "XAxis" of the hyperbola.
    --  The major radius of the hyperbola is on this "XAxis" and 
    --  the minor radius is on the "YAxis" of the hyperbola.
    --  The status is "NegativeRadius" if MajorRadius < 0.0 or if 
    --  MinorRadius < 0.0

Create (Axis        : Ax22d   from gp      ; 
    	MajorRadius : Real    from Standard;
    	MinorRadius : Real    from Standard) returns MakeHyperbola;
    --- Purpose :
    --  Axis is the local coordinate system of the hyperbola.
    --  The major radius of the hyperbola is on this "XAxis" and 
    --  the minor radius is on the "YAxis" of the hyperbola.
    --  The status is "NegativeRadius" if MajorRadius < 0.0 or if 
    --  MinorRadius < 0.0

Create(S1,S2  : Pnt2d from gp;
       Center : Pnt2d from gp) returns MakeHyperbola;
    ---Purpose: Creates a hyperbol centered on the origin of the coordinate system
    --  Axis, with major and minor radii MajorRadius and
    --   MinorRadius, where the major axis is the "X Axis"
    --   of Axis (Axis is the local coordinate system of the hyperbola).
    --   The implicit orientation of the ellipse is:
    -- -   the sense defined by Axis or H,
    -- -   the sense defined by points Center, S1 and S2,
    -- -   the trigonometric sense if Sense is not given or is true, or
    -- -   the opposite sense if Sense is false.
    -- Warning
    -- If an error occurs (that is, when IsDone returns
    -- false), the Status function returns:
    -- -   gce_NegativeRadius if MajorRadius or
    --   MinorRadius is less than 0.0, or
    -- -   gce_InvertAxis if the major radius defined by
    --   Center and S1 is less than the minor radius
    --   defined by Center, S1 and S2.Make an Hyperbola with its center and two apexes.
	          
		
Value(me) returns Hyperbola from Geom2d
    raises NotDone
    is static;
    ---C++: return const&
    ---Purpose: Returns the constructed hyperbola.
    -- Exceptions: StdFail_NotDone if no hyperbola is constructed.
    
Operator(me) returns Hyperbola from Geom2d
    is static;
    ---C++: return const&
    ---C++: alias "Standard_EXPORT operator Handle_Geom2d_Hyperbola() const;"

fields

    TheHyperbola : Hyperbola from Geom2d;
    --The solution from Geom2d.
    
end MakeHyperbola;
