-- Created on: 2003-09-29
-- Created by: Alexander SOLOVYOV and Sergey LITONIN
-- Copyright (c) 2003-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DummySensitiveEntity from MeshVS inherits SensitiveEntity from SelectBasics

	---Purpose: This class allows to create owners to all elements or nodes,
        -- both hidden and shown, but these owners user cannot select "by hands"
        -- in viewer. They means for internal application tasks, for example, receiving
        -- all owners, both for hidden and shown entities.
uses
  EntityOwner   from SelectBasics,
  ListOfBox2d   from SelectBasics,
  PickArgs      from SelectBasics,
  Array1OfPnt2d from TColgp,

  Box2d         from Bnd

is
   Create   ( OwnerId : EntityOwner from SelectBasics ) returns mutable DummySensitiveEntity from MeshVS;

   Areas    ( me: mutable;
              aresult: in out ListOfBox2d from SelectBasics ) is redefined;

   Matches (me : mutable;
            thePickArgs : PickArgs from SelectBasics;
            theMatchDMin, theMatchDepth : out Real from Standard)
    returns Boolean is redefined;

   Matches  ( me: mutable;
              XMin, YMin, XMax, YMax, aTol: Real ) returns Boolean is redefined;

   Matches  ( me: mutable;
              Polyline : Array1OfPnt2d from TColgp;
              aBox     : Box2d from Bnd;
              aTol     : Real    ) returns Boolean is redefined;

   Is3D     ( me ) returns Boolean is redefined;

   NeedsConversion ( me ) returns Boolean is redefined;

   MaxBoxes ( me ) returns Integer is redefined;

end DummySensitiveEntity;
