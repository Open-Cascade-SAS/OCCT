-- Created on: 2002-01-04
-- Created by: data exchange team
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1

class OrientedSurface from StepGeom
inherits Surface from StepGeom

    ---Purpose: Representation of STEP entity OrientedSurface

uses
    HAsciiString from TCollection

is
    Create returns OrientedSurface from StepGeom;
	---Purpose: Empty constructor

    Init (me: mutable; aRepresentationItem_Name: HAsciiString from TCollection;
                       aOrientation: Boolean);
	---Purpose: Initialize all fields (own and inherited)

    Orientation (me) returns Boolean;
	---Purpose: Returns field Orientation
    SetOrientation (me: mutable; Orientation: Boolean);
	---Purpose: Set field Orientation

fields
    theOrientation: Boolean;

end OrientedSurface;
