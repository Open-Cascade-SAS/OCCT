-- Created on: 2002-10-30
-- Created by: Michael SAZONOV
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package BinMDataStd 

        ---Purpose: Storage and Retrieval drivers for modelling attributes.

uses BinMDF,
     BinObjMgt,
     TDF,
     CDM

is
        ---Category: Storage/Retrieval drivers for TDataStd attributes
        --           =======================================

    class NameDriver;

    class IntegerDriver;

    class RealDriver;

    class IntegerArrayDriver;

    class RealArrayDriver;

    class UAttributeDriver;

    class DirectoryDriver;

    class CommentDriver;

    class VariableDriver;

    class ExpressionDriver;

    class RelationDriver;

    class NoteBookDriver;

    class TreeNodeDriver;

    class ExtStringArrayDriver; 

      
    -- Extension 
    
    class TickDriver;  
    
    class AsciiStringDriver;  
    
    class IntPackedMapDriver;
    
    -- Lists: 
    
    class IntegerListDriver; 
    
    class RealListDriver; 
    
    class ExtStringListDriver; 
    
    class BooleanListDriver; 
    
    class ReferenceListDriver;
    
    -- Arrays: 
    
    class BooleanArrayDriver; 
    
    class ReferenceArrayDriver; 
    
    class ByteArrayDriver;  
              
    class NamedDataDriver;  
    
    
    AddDrivers (theDriverTable : ADriverTable  from BinMDF;
                aMsgDrv        : MessageDriver from CDM);
        ---Purpose: Adds the attribute drivers to <theDriverTable>. 
	 
    SetDocumentVersion (DocVersion  : Integer from Standard); 
    
    DocumentVersion returns Integer from Standard; 
    
end BinMDataStd;
