-- Created on: 1997-02-11
-- Created by: Alexander BRIVIN
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Texture2 from Vrml 

	---Purpose: defines a Texture2 node of VRML specifying properties of geometry
	--          and its appearance.
    	--  This  property  node  defines  a  texture  map  and  parameters  for  that  map   
	--  The  texture  can  be  read  from  the  URL  specified  by  the  filename  field. 
	--  To  turn  off  texturing,  set  the  filename  field  to  an  empty  string  ("").
    	--  Textures  can  alsobe  specified  inline  by  setting  the  image  field   
	--  to  contain  the  texture  data.  
    	--  By  default  : 
	--    myFilename ("")
	--    myImage (0 0 0)
	--    myWrapS (Vrml_REPEAT)
	--    myWrapT (Vrml_REPEAT) 

uses
 
    SFImage      from  Vrml, 
    Texture2Wrap from  Vrml, 
    AsciiString  from  TCollection

is
 
    Create  returns  Texture2 from Vrml;
 
    Create  (  aFilename : AsciiString from TCollection; 
    	       aImage    : SFImage      from  Vrml; 
    	       aWrapS    : Texture2Wrap from  Vrml; 
    	       aWrapT    : Texture2Wrap from  Vrml) 
    	returns  Texture2 from Vrml;

    SetFilename   ( me : in out; aFilename : AsciiString from TCollection );
    Filename   ( me )  returns  AsciiString from TCollection;
 
    SetImage   ( me : in out; aImage : SFImage  from  Vrml );
    Image   ( me )  returns SFImage  from  Vrml;

    SetWrapS   ( me : in out; aWrapS : Texture2Wrap from  Vrml );
    WrapS   ( me )  returns  Texture2Wrap from  Vrml;

    SetWrapT   ( me : in out; aWrapT : Texture2Wrap from  Vrml );
    WrapT   ( me )  returns  Texture2Wrap from  Vrml;

    Print  ( me;  anOStream: in out OStream from Standard) returns OStream from Standard;
    ---C++:  return  & 

fields
 
    myFilename  :  AsciiString  from  TCollection;	-- file to read texture from
    myImage     :  SFImage      from  Vrml;      	-- The texture
    myWrapS     :  Texture2Wrap from  Vrml;
    myWrapT     :  Texture2Wrap from  Vrml;

end Texture2;
