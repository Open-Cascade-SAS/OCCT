-- Created on: 2002-12-10
-- Created by: data exchange team
-- Copyright (c) 2002-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V2.0

class SymmetricTensor23d from StepFEA
inherits SelectType from StepData

    ---Purpose: Representation of STEP SELECT type SymmetricTensor23d

uses
    SelectMember from StepData,
    HArray1OfReal from TColStd,
    HArray1OfReal from TColStd

is
    Create returns SymmetricTensor23d from StepFEA;
	---Purpose: Empty constructor

    CaseNum (me; ent: Transient) returns Integer;
	---Purpose: Recognizes a kind of SymmetricTensor23d select type
	--          return 0 

    CaseMem (me; ent: SelectMember from StepData) returns Integer is redefined;
	---Purpose: Recognizes a items of select member SymmetricTensor23dMember
	--          1 -> IsotropicSymmetricTensor23d
	--          2 -> OrthotropicSymmetricTensor23d
	--          3 -> AnisotropicSymmetricTensor23d
	--          0 else


     NewMember(me) returns SelectMember from StepData is redefined;
	---Purpose: Returns a new select member the type SymmetricTensor23dMember

    SetIsotropicSymmetricTensor23d(me: in out; aVal :Real);
	---Purpose: Set Value for IsotropicSymmetricTensor23d

    IsotropicSymmetricTensor23d (me) returns Real;
	---Purpose: Returns Value as IsotropicSymmetricTensor23d (or Null if another type)

    SetOrthotropicSymmetricTensor23d(me: in out; aVal :HArray1OfReal from TColStd);
	---Purpose: Set Value for OrthotropicSymmetricTensor23d

    OrthotropicSymmetricTensor23d (me) returns HArray1OfReal from TColStd;
	---Purpose: Returns Value as OrthotropicSymmetricTensor23d (or Null if another type)

    SetAnisotropicSymmetricTensor23d(me: in out; aVal :HArray1OfReal from TColStd);
	---Purpose: Set Value for AnisotropicSymmetricTensor23d

    AnisotropicSymmetricTensor23d (me) returns HArray1OfReal from TColStd;
	---Purpose: Returns Value as AnisotropicSymmetricTensor23d (or Null if another type)

end SymmetricTensor23d;
