-- Created on: 1993-01-09
-- Created by: CKY / Contract Toubro-Larsen ( SIVA )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class ConeFrustum from IGESSolid  inherits IGESEntity

        ---Purpose: defines ConeFrustum, Type <156> Form Number <0>
        --          in package IGESSolid
        --          The Cone Frustum is defined by the center of the
        --          larger circular face of the frustum, its radius, a unit
        --          vector in the axis direction, a height in this direction
        --          and a second circular face with radius which is lesser
        --          than the first face.

uses

        Pnt             from gp,
        Dir             from gp,
        XYZ             from gp

is

        Create returns mutable ConeFrustum;

        -- Specific Methods pertaining to the class

        Init (me     : mutable;
              Ht     : Real;
              R1     : Real;
              R2     : Real;
              Center : XYZ;
              anAxis : XYZ);
        ---Purpose : This method is used to set the fields of the class
        --           ConeFrustum
        --       - Ht     : the Height of cone
        --       - R1     : Radius of the larger face
        --       - R2     : Radius of the smaller face (default 0)
        --       - Center : Center of the larger face (default (0,0,0))
        --       - anAxis : Unit vector in axis direction (default (0,0,1))

        Height (me) returns Real;
        ---Purpose : returns the height of the cone frustum

        LargerRadius (me) returns Real;
        ---Purpose : returns the radius of the larger face of the cone frustum

        SmallerRadius (me) returns Real;
        ---Purpose : returns the radius of the second face of the cone frustum

        FaceCenter (me) returns Pnt;
        ---Purpose : returns the center of the larger face of the cone frustum

        TransformedFaceCenter (me) returns Pnt;
        ---Purpose : returns the center of the larger face of the cone frustum
        -- after applying TransformationMatrix

        Axis (me) returns Dir;
        ---Purpose : returns the direction of the axis of the cone frustum

        TransformedAxis (me) returns Dir;
        ---Purpose : returns the direction of the axis of the cone frustum
        -- after applying TransformationMatrix

fields

--
-- Class    : IGESSolid_ConeFrustum
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class ConeFrustum.
--
-- Reminder : A ConeFrustum instance is defined by :
--            The Cone Frustum is defined by the center of the
--            larger circular face of the frustum(X1,Y1,Z1), its radius(R1),
--            a unit vector in the axis direction(I1,J1,K1),a height in this
--            direction(Height) and a second circular face with radius(R2)
--            R1 > R2
--

        theHeight     : Real;

        theR1         : Real;
            -- the radius of the larger face of the cone frustum

        theR2         : Real;
            -- the radius of the smaller face of the cone frustum
    
        theFaceCenter : XYZ;
            --  the larger face center coordinates

        theAxis       : XYZ;
            --  the Unit vector in axis direction

end ConeFrustum;
