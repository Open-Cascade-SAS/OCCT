-- Created on: 1992-04-29
-- Created by: Remi LEQUETTE
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Text3D from Draw inherits Drawable3D from Draw

	---Purpose: 

uses Pnt from gp,
    Color from Draw,
    Display from Draw,
    AsciiString from TCollection

is

    Create(p : Pnt; T : CString; col : Color)
    returns mutable Text3D from Draw;
    
    Create(p : Pnt; T : CString; col : Color;
    	   moveX : Real; moveY : Real)
    returns mutable Text3D from Draw;

    SetPnt(me : mutable; p : Pnt);
   
    DrawOn(me; dis : in out Display);

fields

    myPoint : Pnt          from gp;
    myColor : Color        from Draw;
    myText  : AsciiString  from TCollection;
    mymoveX : Real      from Standard;
    mymoveY : Real      from Standard;
    
end Text3D;
