-- Created on: 1992-04-07
-- Created by: Christian CAILLET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class NameEntity  from IGESData  inherits IGESEntity

    ---Purpose : a NameEntity is a kind of IGESEntity which can provide a Name
    --           under alphanumeric (String) form, from Properties list
    --           an effective Name entity must inherit it

uses  HAsciiString from TCollection

is

    Value (me) returns HAsciiString from TCollection  is deferred;
    ---Purpose : Retyrns the alphanumeric value of the Name, to be defined

end NameEntity;
