-- Created on: 1999-01-25
-- Created by: Xuan PHAM PHU
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class TOOL from TopOpeBRepDS
uses
    Edge from TopoDS,
    Shape from TopoDS,
    ListOfShape from TopTools,
    Config from TopOpeBRepDS,
    HDataStructure from TopOpeBRepDS,
    DataMapOfShapeListOfShapeOn1State from TopOpeBRepDS
is

    EShareG(myclass; HDS : HDataStructure; E: Edge from TopoDS; 
     	    lEsd : out ListOfShape from TopTools)
    returns Integer;
    -- Fills up <lEsd> with edges sharing geometric domain with <E>, 
    -- using interferences attached to <E>.
    -- Returns <lEsd>'s length.

    ShareG(myclass; HDS : HDataStructure; is1,is2 : Integer)
    returns Boolean;
    -- Returns true if shapes <is1> and <is2> share geometric domain.

    GetEsd(myclass; HDS : HDataStructure; S : Shape; ie : Integer; iesd : out Integer)
    returns Boolean;
    -- Gets edge<iesd> in shape <S>, edge<ie> shares geometric domain with edge<iesd>
    -- Returns true if <iesd> is found

    ShareSplitON(myclass; HDS : HDataStructure; MspON : DataMapOfShapeListOfShapeOn1State;
    	      	 i1, i2 : Integer; spON : out Shape)
    returns Boolean;
    -- Gets <spON> splitON shared  by  shapes  <i1>  an <i2> (shapes same domain) 
    -- Returns true if <spON> is found.

    GetConfig(myclass; HDS : HDataStructure; MEspON : DataMapOfShapeListOfShapeOn1State;
    	      ie, iesd : Integer; conf : out Integer)
    returns Boolean;
    -- Gives relative orientation conf = 1 : SAMEORIENTED
    --                                   2 : DIFFORIENTED.
    -- edges <ie>, <iesd> are same domain.
    -- Returns true if <conf> is found.

end TOOL;
