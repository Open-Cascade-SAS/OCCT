-- Created on: 1996-01-09
-- Created by: Denis PASCAL
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class PlanarDimension from DrawDim inherits Dimension from DrawDim

	---Purpose: Dimensions between point, line and circle ON a plane

uses Face from TopoDS

is

    SetPlane (me : mutable; plane : Face from TopoDS);
    
    GetPlane (me)
    returns Face from TopoDS;


--    Point (myclass; s : Shape from TopoDS; p : in out Pnt from gp)

--    returns Boolean from Standard;    


--    Line (myclass; s : Shape from TopoDS; l : in out Lin from gp)

--    returns Boolean from Standard;    


--    Circle (myclass; s : Shape from TopoDS; c : in out Circ from gp)

--    returns Boolean from Standard;    


--    Ellipse (myclass; s : Shape from TopoDS; c : in out Elips from gp)

--    returns Boolean from Standard;


fields

    myPlane : Face from TopoDS  is protected;
    
end PlanarDimension;
