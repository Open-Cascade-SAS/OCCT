-- Created on: 1995-04-25
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Builder from LocOpe

	---Purpose: Provides    a  basic  tool    to  implement  local
	--          topological operations.

uses
    Shape          from TopoDS,
    ListOfShape    from TopTools,
--    HBuilder       from TopOpeBRepBuild,
--    DSAccess       from BRepAlgo,
    HistoryCollector from BOP,
    TopOpe         from BRepAlgo, 
    MapOfShape     from TopTools  
  
     
raises
    NotDone           from StdFail,
    ConstructionError from Standard


is

    Create
	---Purpose: Empty constructor.
    	returns Builder from LocOpe;
	
	
    Create(S: Shape from TopoDS)
	---Purpose: Creates a builder for local operations on <S>.
    	returns Builder from LocOpe
	raises ConstructionError from Standard;
	--- The exception is raised if <S> is a null shape.


    Create(S: Shape from TopoDS; Tool: Shape from TopoDS)
	---Purpose: Creates a builder for local operations between <S>
	--          and  <Tool>.
    	returns Builder from LocOpe
	raises ConstructionError from Standard;
	--- The exception is raised if <S> or <Tool> is a null shape .


    Init(me: in out; S: Shape from TopoDS)
	---Purpose: Initializes a builder for local operations on <S>.
	raises ConstructionError from Standard
	--- The exception is raised if <S> is a null shape.
    	is static;


    Init(me: in out; S: Shape from TopoDS; Tool: Shape from TopoDS)
	---Purpose: Initializes a builder for local operations between
	--          <S>  and <Tool>.
	raises ConstructionError from Standard
	--- The exception is raised if <S> or <Tool>is a null shape.
    	is static;


    Perform(me: in out; Tool : Shape       from TopoDS;
                        L    : ListOfShape from TopTools;
                        Fuse : Boolean     from Standard)

	---Purpose: Performs the local operation on the formerly given
	--          shape.  <L> defines   a   set  of faces  of    the
	--          shape. The whole tool is used. The list may not be
	--          empty.   The  boolean  <Fuse>   gives the type  of
	--          operation. If set  to Standard_True, the operation
	--          is  a fusion.    If  set  to   Standard_False, the
	--          operation is a cutting one.
	--          
	--          The Perform process stops just before constructing
	--          any result in order to authorize  the selection of
	--          parts of the tool.  After a call to Perform, it is
	--          possible   to call     BuilPartsOfTool,       then
	--          RemovePart/ActivatePart to select valid parts, and
	--          it  is necessary to  call PerformResult to get any
	--          result. 

    	raises ConstructionError from Standard
	-- The exception is raised if <Tool> is null or same as the shape.

    	is static;


    Perform(me: in out; LShape : ListOfShape from TopTools;
                        LTool  : ListOfShape from TopTools;
                        Fuse   : Boolean from Standard)

	---Purpose: Performs the local operation on the formerly given
	--          shape and tool.  <LShape>  defines a set  of faces
	--          of  the shape.  <LTool> defines  a set of faces of
	--          the  tool.  The boolean  <Fuse>  gives the type of
	--          operation.  If set to Standard_True, the operation
	--          is  a  fusion.    If set   to  Standard_False, the
	--          operation   is  a cutting  one. If <LShape> (resp.
	--          <LTool>) is empty, the whole shape (resp. tool) is
	--          used. 
	--          
	--          The Perform process stops just before constructing
	--          any result in order to authorize  the selection of
	--          parts of the tool.  After a call to Perform, it is
	--          possible   to call     BuilPartsOfTool,       then
	--          RemovePart/ActivatePart to select valid parts, and
	--          it  is necessary to  call PerformResult to get any
	--          result. 

    	is static;



    BuildPartsOfTool(me: in out)
	---Purpose: Builds every valid parts of the tool.
    	raises NotDone from StdFail
	-- The exception is raised if no call to Perform has been done.
    	is static;
    

    PartsOfTool(me)
	---Purpose: Returns  the list of  the  parts of tool.  Each of
	--          this part is a TopoDS_Shell.
    	returns ListOfShape from TopTools
	---C++: return const&
    	raises NotDone from StdFail
	-- The exception is raised if no  call to BuildPartsOfTool has
	-- been done. 
	is static;


    RemovePart(me: in out; S: Shape from TopoDS)
	---Purpose: Removes <S> from the list of valid parts of tool.
    	raises NotDone from StdFail
	-- The exception is raised if no  call to BuildPartsOfTool has
	-- been done. 
    	is static;


    ActivatePart(me: in out; S: Shape from TopoDS)
	---Purpose: Removes <S>  from  the list  of  invalid parts  of
	--          tool. By default, all parts  of tool are valid for
	--          the local operation.
    	raises NotDone from StdFail
	-- The exception is raised if no  call to BuildPartsOfTool has
	-- been done. 
    	is static;
	
	

    PerformResult(me: in out)
	---Purpose: Invalidates the given parts of  tools if any,  and
	--          performs the result of the local operation.
    	raises NotDone from StdFail
	-- The exception is raised if no call to Perform has been done.
    	is static;


    IsDone(me)
	---Purpose: Returns  Standard_True  if the operation  has been
	--          successfuly done.
    	returns Boolean from Standard
	---C++: inline
	is static;

    IsInvDone(me)
	---Purpose: Returns  Standard_True  if the Invalidate Parts 
	--          operation  has been successfuly done.
    	returns Boolean from Standard
	---C++: inline
	is static;

    ResultingShape(me)
	---Purpose: Returns the result of the operation.

    	returns Shape from  TopoDS
	---C++: return const&
	---C++: inline
	raises NotDone from StdFail
	-- The exception is raised if IsDone returns Standard_False.
	is static;
    
    
    OriginalShape(me)
	---Purpose: Returns the shape on which the operation is defined.
    	returns Shape from TopoDS
	---C++: return const&
	---C++: inline
	is static;


    Tool(me)
	---Purpose: Returns the "tool" used to perform the local operation.
    	returns Shape from TopoDS
	---C++: return const&
	---C++: inline
	is static;


--    Builder(me)  
--    	returns HBuilder from TopOpeBRepBuild

    History(me)	    
    	returns HistoryCollector from BOP
	---C++: inline
	---C++: return const&
	is static;


--- Private implementation methods
--  

    InvalidateParts(me: in out)
    
    	is static;

    Edges(me)

    	returns ListOfShape from TopTools
	---C++: return const&
	is static;
	
    TgtEdges(me)

    	returns ListOfShape from TopTools
	---C++: return const&
	is static;


fields

    myDone    : Boolean        from Standard;
    myShape   : Shape          from TopoDS;
    myTool    : Shape          from TopoDS;
    myResult  : Shape          from TopoDS;
    myParts   : ListOfShape    from TopTools;
    myRemoved : ListOfShape    from TopTools;
    myPdone   : Boolean        from Standard;
    myPerfdone: Boolean        from Standard;
    myInvDone : Boolean        from Standard;
    myFuse    : Boolean        from Standard;
    myEdges   : ListOfShape    from TopTools;
    myTgtEdges: ListOfShape    from TopTools;
--    myAlgo    : DSAccess       from BRepAlgo;
    myAlgo    : TopOpe         from BRepAlgo;
    myShapeMap: MapOfShape     from TopTools;
    myToolMap : MapOfShape     from TopTools;

end Builder;



