-- File:        BoundaryCurve.cdl
-- Created:     Fri Dec  1 11:11:15 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class BoundaryCurve from StepGeom 

inherits CompositeCurveOnSurface from StepGeom 

uses

	HAsciiString from TCollection, 
	HArray1OfCompositeCurveSegment from StepGeom, 
	Logical from StepData
is

	Create returns mutable BoundaryCurve;
	---Purpose: Returns a BoundaryCurve


end BoundaryCurve;
