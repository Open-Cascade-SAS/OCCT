-- File:	BRepExtrema_ExtPC.cdl
-- Created:	Fri Dec  3 16:01:30 1993
-- Author:	Christophe MARION
--		<cma@sdsun1>
---Copyright:	 Matra Datavision 1993

class ExtPC from BRepExtrema

uses
    Integer from Standard,
    Real    from Standard,
    Boolean from Standard,
    Vertex  from TopoDS,
    Edge    from TopoDS,
    ExtPC   from Extrema,
    Pnt     from gp,
    HCurve  from BRepAdaptor
     
raises 
    NotDone      from StdFail,
    OutOfRange   from Standard,
    TypeMismatch from Standard

is
    Create returns ExtPC from BRepExtrema;

    Create(V : Vertex from TopoDS;
           E : Edge   from TopoDS)
    	---Purpose: It calculates all the distances.
    returns ExtPC from BRepExtrema;

    Initialize(me: in out; E : Edge from TopoDS)
    	---Purpose: 
    is static;
    
    Perform(me: in out; V : Vertex from TopoDS)
    	---Purpose: An exception is raised if the fields have not been
    	--          initialized.
    raises TypeMismatch from Standard
    is static;
    
    IsDone(me) returns Boolean from Standard
    	---Purpose: True if the distances are found.
    is static;
    
    NbExt(me) returns Integer from Standard
    	---Purpose: Returns the number of extremum distances.
    raises NotDone from StdFail
    is static;

    IsMin(me; N : Integer from Standard) returns Boolean from Standard
    	---Purpose: Returns True if the <N>th extremum distance is a
    	--          minimum.
    raises NotDone    from StdFail,
    	   OutOfRange from Standard
    is static;
    
    SquareDistance(me; N : Integer from Standard) returns Real from Standard
    	---Purpose: Returns the value of the <N>th extremum square distance.
    raises NotDone    from StdFail,
    	   OutOfRange from Standard
    is static;
    
    Parameter(me; N : Integer from Standard) returns Real from Standard
    	---Purpose: Returns the parameter  on the  edge  of the  <N>th
    	--          extremum distance.
    raises NotDone    from StdFail,
    	   OutOfRange from Standard
    is static;
    
    Point(me; N : Integer from Standard) returns Pnt from gp
    	---Purpose: Returns the Point of the <N>th extremum distance.
    raises NotDone    from StdFail, 
    	   OutOfRange from Standard
    is static;
    
    TrimmedSquareDistances(me; dist1 : out Real from Standard;
                         dist2 : out Real from Standard;
                         pnt1  : out Pnt  from gp;
                         pnt2  : out Pnt  from gp)
    	---Purpose: if the curve is a trimmed curve,
    	--          dist1 is a square distance between <P> and the point
    	--          of parameter FirstParameter <pnt1> and
    	--          dist2 is a square distance between <P> and the point
    	--          of parameter LastParameter <pnt2>.
    is static;
    
fields
    myExtrem  : ExtPC  from Extrema;
    myHC      : HCurve  from BRepAdaptor;
end ExtPC;
