-- Created on: 1992-05-07
-- Created by: Modelistation
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package StdFail 

uses Standard

is

    exception NotDone inherits Failure from Standard;
    exception Undefined inherits Failure from Standard;
    exception UndefinedDerivative inherits DomainError from Standard;
    exception UndefinedValue inherits DomainError from Standard;
    exception InfiniteSolutions inherits Failure from Standard;

end StdFail;

    


