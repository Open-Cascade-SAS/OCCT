-- Created on: 1993-10-14
-- Created by: Christian CAILLET
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class ToolReferenceDesignator  from IGESAppli

    ---Purpose : Tool to work on a ReferenceDesignator. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses ReferenceDesignator from IGESAppli,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolReferenceDesignator;
    ---Purpose : Returns a ToolReferenceDesignator, ready to work


    ReadOwnParams (me; ent : mutable ReferenceDesignator;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : ReferenceDesignator;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : ReferenceDesignator;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a ReferenceDesignator <ent>, from
    --           its specific (own) parameters

    OwnCorrect (me; ent : mutable ReferenceDesignator) returns Boolean  is static;
    ---Purpose : Sets automatic unambiguous Correction on a ReferenceDesignator
    --           (NbPropertyValues forced to 1, Level cleared if Subordinate != 0)

    DirChecker (me; ent : ReferenceDesignator) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : ReferenceDesignator;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : ReferenceDesignator; entto : mutable ReferenceDesignator;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : ReferenceDesignator;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolReferenceDesignator;
