-- Created on: 1996-08-30
-- Created by: Xavier BENVENISTE
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Interpolate from GeomLib

	---Purpose: this class is used to construct a BSpline curve by
	--          interpolation  of points  at given parameters  The
	--          continuity   of the curve   is degree -  1 and the
	--          method used when boundary  condition are not given
	--          is to use odd degrees  and null the derivatives on
	--          both sides from degree -1 down to (degree+1) / 2
	--          When even degree is given the returned curve is of
	--          degree - 1 so that the degree of the curve is odd 
    	

uses
    Array1OfPnt         from TColgp,
    Array1OfReal        from TColStd,
    InterpolationErrors from GeomLib,
    BSplineCurve        from Geom

raises

    NotDone    from StdFail,
    OutOfRange from Standard
    
is

    Create( Degree     : Integer from Standard ;
    	    NumPoints  : Integer from Standard ;
	    Points     : Array1OfPnt from TColgp ;
	    Parameters : Array1OfReal from TColStd) 
	     
    returns Interpolate from GeomLib ;
    
    IsDone(me) returns Boolean from Standard
    	---Purpose: 
    	-- returns if everything went OK
	---C++: inline
    is static;


    Error(me) returns InterpolationErrors from GeomLib 
    ---Purpose: returns the error type if any 
    ---C++: inline	      
    --          
    is static ;

    Curve(me) 
    ---Purpose:  returns the interpolated curve of the requested degree 

    returns BSplineCurve from Geom
    raises
    	OutOfRange from Standard,
	NotDone    from StdFail
    is static;
 
    
    
fields

    myCurve : BSplineCurve from Geom ;
    myIsDone : Boolean from Standard ;
    myError  : InterpolationErrors  from GeomLib  ;
    
end Interpolate ;

