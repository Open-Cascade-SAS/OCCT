-- Created on: 2004-02-04
-- Created by: Sergey KUUL
-- Copyright (c) 2004-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SplitCommonVertex from ShapeFix inherits Root from ShapeFix

	---Purpose: Two wires have common vertex - this case is valid in BRep model
        --          and isn't valid in STEP => before writing into STEP it is necessary
        --          to split this vertex (each wire must has one vertex)

uses
    Shape from TopoDS
    
is
    Create returns SplitCommonVertex;
    ---Purpose :

    Init(me: mutable; S : Shape from TopoDS); 
    ---Purpose :
    
    Perform(me:mutable);	
    ---Purpose :
    
    Shape(me : mutable) returns Shape from TopoDS;
    ---Purpose :

fields

    myShape    : Shape from TopoDS;
    myResult   : Shape from TopoDS;
    myStatus   : Integer; -- error status

end SplitCommonVertex;
