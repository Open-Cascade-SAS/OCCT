-- Created on: 1997-10-29
-- Created by: Roman BORISOV
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred  class SparseMatrix from FEmTool  inherits  TShared  from  MMgt

	---Purpose: Sparse Matrix definition

uses 
    Vector  from  math

raises   
    NotDone  from  StdFail	
   
is    
    Init(me:  mutable;  Value  :  Real) 
    is  deferred; 
     
    ChangeValue(me:  mutable;  I,  J  :  Integer) 
     ---C++: return &
    returns  Real is  deferred; 
     
    Decompose(me  :  mutable)   
    ---Purpose: To make a Factorization of <me>
    returns  Boolean
    is  deferred;
        
    Solve(me;  B  :  Vector;  X  :  in  out  Vector) 
    ---Purpose: Direct Solve of AX = B   
    raises  NotDone from  StdFail --  if  <me> is not decomposed
    is  deferred;  
     
    Prepare(me  :  mutable) 
     ---Purpose: Make Preparation to iterative solve  
    returns  Boolean
    is  deferred;
     
    Solve(me;  B          :  Vector;   
               Init       :  Vector;  
	       X          :  out  Vector;
               Residual   :  out  Vector; 
               Tolerance  :  Real  =  1.0e-8;
	       NbIterations: Integer = 50)
    ---Purpose: Iterative solve  of AX = B
    raises  NotDone from  StdFail  --  if  <me> is not prepared;
    is  deferred;  
     
    
    Multiplied(me; X: Vector; MX  :  in  out  Vector) 
    ---Purpose: returns the product of a SparseMatrix by a vector.
    --          An exception is raised if the dimensions are different
    is  deferred;    
    
    RowNumber(me)
    	---Purpose: returns the row range of a matrix.
    returns Integer
    is deferred;

    
    ColNumber(me)
    	---Purpose: returns the column range of the matrix.
    returns Integer
    is deferred;  
  
end SparseMatrix;
