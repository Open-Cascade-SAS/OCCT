-- File:        OpenShell.cdl
-- Created:     Mon Dec  4 12:02:28 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWOpenShell from RWStepShape

	---Purpose : Read & Write Module for OpenShell

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     OpenShell from StepShape,
     EntityIterator from Interface

is

	Create returns RWOpenShell;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable OpenShell from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : OpenShell from StepShape);

	Share(me; ent : OpenShell from StepShape; iter : in out EntityIterator);

end RWOpenShell;
