-- Created on: 1996-09-18
-- Created by: Jacques MINOT
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class OffsetPresentation from DsgPrs

        ---Purpose: A framework to define display of offsets.
uses
    Presentation from Prs3d,
    Pnt from gp,
    Dir from gp,
    Drawer from Prs3d,
    ExtendedString from TCollection,
    ArrowSide from DsgPrs
is  
    Add( myclass; aPresentation: Presentation from Prs3d;
    	    	  aDrawer: Drawer from Prs3d;
		  aText: ExtendedString from TCollection;
                  AttachmentPoint1: Pnt from gp;
		  AttachmentPoint2: Pnt from gp;
		  aDirection: Dir from gp;
		  aDirection2: Dir from gp;
		  OffsetPoint: Pnt from gp);
	---Purpose: Defines the display of elements showing offset shapes.
    	-- These include the two points of attachment
    	-- AttachmentPoint1 and AttachmentPoint1, the two
    	-- directions aDirection and aDirection2, and the offset point OffsetPoint.
    	-- These arguments are added to the presentation
    	-- object aPresentation. Their display attributes are
    	-- defined by the attribute manager aDrawer.

    AddAxes( myclass; aPresentation: Presentation from Prs3d;
    	    	  aDrawer: Drawer from Prs3d;
		  aText: ExtendedString from TCollection;
                  AttachmentPoint1: Pnt from gp;
		  AttachmentPoint2: Pnt from gp;
		  aDirection: Dir from gp;
		  aDirection2: Dir from gp;
		  OffsetPoint: Pnt from gp);
	---Purpose: draws the representation of axes alignement Constraint
	--          between the point AttachmentPoint1 and the
	--          point AttachmentPoint2, along direction 
	--          aDirection, using the offset point OffsetPoint.

end OffsetPresentation;
