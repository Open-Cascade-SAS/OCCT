-- Created on: 1992-03-04
-- Created by: Laurent BUCHARD
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package IntCurve

    ---Purpose: This package provides algorithmes to intersect 2D curves,
    --          with domains.
    --          
    --          class IntConicConic : Algorithm used to intersect 2 conics 
    --                                from gp with domains.
    --                                
    --          class IntConicCurveGen : Generic algorithm used to intersect 
    --                                   a conic from gp, and a parametrised
    --                                   curve.
    --                                   The parametrised Curve can 
    --                                   not be a Composite curve and 
    --                                   can not be a conic.
    --                                   
    --          class IntCurveCurveGen : Generic algorithm used to intersect 2
    --                                   curves. The resources on a curve are
    --                                   discribed in the class CurveTool.
    --
    --          class UserIntConicCurveGen: Generic algorithm used to  
    --                                      intersect a Conic from gp 
    --                                      and a parametrised curve. 
    --                                      This curve can be either a  
    --                                      composite curve or a conic. 
    --


    ---Level: Advanced 
    -- 
    -- The Classes <PConicTool,
    --              IConicTool,
    --              PConic,
    --              ProjectOnPConicTool,
    --              IntConicCurveGen, 
    --              ProjPCurGen,
    --              UserIntConicCurveGen,
    --              IntPolyPolyGen,
    --              Polygon2dGen,
    --              DistBetweenPCurvesGen>    are  Internal 
    --
    -- The Classe   <IntCurveCurveGen>        is   Advanced 
    --
    --



uses Standard , math, gp, TColgp, GeomAbs,
     IntImpParGen, IntRes2d, Extrema,
     StdFail, Bnd, Intf, TColStd
     

is 

    class IntConicConic;
    ---Purpose: Intersection between 2 conics from gp.

    generic class DistBetweenPCurvesGen;
    
    generic class Polygon2dGen;

    generic class IntPolyPolyGen,ThePolygon2d,
                                 TheDistBetweenPCurves, 
    	    	    	    	 ExactIntersectionPoint;

    generic class UserIntConicCurveGen;

    generic class ProjPCurGen,TheCurveLocator,TheLocateExtPC;
    
    generic class IntConicCurveGen,TheIntersector;
    ---Purpose: Intersection between a conic from gp and a bounded parametric curve.

    generic class IntCurveCurveGen,TheProjPCur,
                                   TheIntConicCurve,
                                   IntConicCurve,
                                   TheIntPCurvePCurve;
				   
    ---Purpose: Intersection between 2 2d curves.
    
    private class ProjectOnPConicTool;
    
    class PConic;

    class IConicTool;

    private class PConicTool;
	      
    private class IntImpConicParConic
         instantiates Intersector from IntImpParGen
             (IConicTool           from IntCurve,
	      PConic               from IntCurve,
	      PConicTool           from IntCurve,
    	      ProjectOnPConicTool  from IntCurve);
	

 	
end IntCurve;    

