-- Created on: 1991-06-24
-- Created by: Christophe MARION
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- modified by jct (15/04/97)  add of  ModificationCommands




package GeomliteTest 

	---Purpose: this  package  provides  elementary commands for  curves  and
	--          surface.
uses
    Draw,
    Standard

is

    AllCommands(I : in out Interpretor from Draw);
	---Purpose: defines all geometric commands.
    
    CurveCommands(I : in out Interpretor from Draw);
	---Purpose: defines curve commands.
    
    SurfaceCommands(I : in out Interpretor from Draw);
	---Purpose: defines surface commands.
    
    API2dCommands(I : in out Interpretor from Draw);
	---Purpose: defines commands to test the Geom2dAPI
	--          - Intersection
	--          - Extrema
	--          - Projection
	--          - Approximation, interpolation 
    ApproxCommands(I : in out Interpretor from Draw);
	---Purpose: defines constrained curves commands.

    ModificationCommands(I : in out Interpretor from Draw);
	---Purpose: defines curves and surfaces modification commands.
	--          - Curve extension to point
	--          - Surface extension by length
    
    
end GeomliteTest;
