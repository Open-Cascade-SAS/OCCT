-- Created on: 1992-11-17
-- Created by: Remi LEQUETTE
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




generic class FaceClassifier from TopClass 
    (TheFaceExplorer as any;
     TheEdge as any;
     TheIntersection2d as any)

	---Purpose: Provides an algorithm to classify a  point in a 2D
	--          face (or in the UV space of a face on a surface).

uses
    Pnt2d from gp,
    Position from IntRes2d,
    State from TopAbs
    
raises
    DomainError

    class FClass2d instantiates Classifier2d from TopClass
    	(TheEdge, TheIntersection2d);

is
    Create returns FaceClassifier from TopClass;
	---Purpose: Empty constructor, undefined algorithm.
	
    Create(F : in out TheFaceExplorer; P : Pnt2d from gp; Tol : Real)
    returns FaceClassifier from TopClass;
	---Purpose: Creates an algorithm to classify the Point  P with
	--          Tolerance <T> on the face described by <F>.
	
    Perform(me : in out;
    	    F : in out TheFaceExplorer; P : Pnt2d from gp; Tol : Real)
	---Purpose: Classify  the Point  P  with  Tolerance <T> on the
	--          face described by <F>.
    is static;
    
    State(me) returns State from TopAbs
	---Purpose: Returns the result of the classification.
    is static;
    
    Rejected(me) returns Boolean
	---Purpose: Returns  True when  the   state was computed by  a
	--          rejection. The state is OUT.
	---C++: inline
    is static;
    
    NoWires(me) returns Boolean
	---Purpose: Returns True if  the face  contains  no wire.  The
	--          state is IN.
	---C++: inline
    is static;
    
    Edge(me) returns TheEdge
	---Purpose: Returns   the    Edge  used   to    determine  the
	--          classification. When the State is ON  this  is the
	--          Edge containing the point.
	---C++: return const &
    raises
    	DomainError -- when no edge was used (rejected or nowires)
    is static;
    
    EdgeParameter(me) returns Real from Standard
	---Purpose: Returns the parameter on Edge() used to determine  the
	--          classification.
    raises
    	DomainError -- when no edge was used (rejected or nowires)
    is static;
    
    Position(me) returns Position from IntRes2d
	---Purpose: Returns the  position of  the   point on the  edge
	--          returned by Edge.
	---C++: inline
    is static;
	
fields

    myClassifier    : FClass2d  is protected;
    myEdge          : TheEdge  is protected;
    myEdgeParameter : Real from Standard  is protected;
    myPosition      : Position from IntRes2d  is protected;
    rejected        : Boolean from Standard  is protected;
    nowires         : Boolean from Standard  is protected;

end FaceClassifier;

