-- Created on: 1995-09-01
-- Created by: Bruno DUMORTIER
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class OffsetAncestors from BRepFill 

	---Purpose: this class is used to find the generating shapes
	--          of an OffsetWire.

uses
    OffsetWire          from BRepFill,
    Shape               from TopoDS,
    Edge                from TopoDS,	
    DataMapOfShapeShape from TopTools
    
raises
    NotDone from StdFail
    
is
    Create returns OffsetAncestors from BRepFill;
    
    Create ( Paral : in out OffsetWire from BRepFill)
    returns OffsetAncestors from BRepFill;
    
    Perform ( me : in out; Paral : in out OffsetWire from BRepFill)
    is static;
    
    IsDone( me)
    returns Boolean from Standard
    is static;

    HasAncestor (me; S1 : Edge from TopoDS)	    
    returns Boolean from Standard
    is static;

    Ancestor    (me ; S1 : Edge from TopoDS)
	---Purpose: may return a Null Shape if S1 is not a subShape
	--          of <Paral>;
	---C++: return const &
    returns Shape from TopoDS
    raises
    	NotDone from StdFail
	---Purpose: if Perform is not done.
    is static;
    
fields

    myIsPerform : Boolean             from Standard;
    myMap       : DataMapOfShapeShape from TopTools;
    
end OffsetAncestors;
