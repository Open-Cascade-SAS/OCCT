-- Created on: 1994-11-30
-- Created by: Frederic MAUPAS
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MakeStepFace from TopoDSToStep 
    inherits Root from TopoDSToStep

    ---Purpose: This class implements the mapping between classes 
    --          Face from TopoDS and TopologicalRepresentationItem from
    --          StepShape. 
  
uses Face                          from TopoDS,
     TopologicalRepresentationItem from StepShape,
     Tool                          from TopoDSToStep,
     MakeFaceError                 from TopoDSToStep,
     FinderProcess                 from Transfer
          
raises NotDone from StdFail
     
is 

    Create returns MakeStepFace;
    
    Create (F           : Face from TopoDS;
            T           : in out Tool from TopoDSToStep;
            FP          : FinderProcess from Transfer)
         returns MakeStepFace;
    
    Init(me          : in out;
         F           : Face from TopoDS;
         T           : in out Tool from TopoDSToStep;
         FP          : FinderProcess from Transfer);
	    	    
    Value (me) returns TopologicalRepresentationItem from StepShape
    	raises NotDone
    	is static;
    	---C++: return const&
    
    Error(me) returns MakeFaceError from TopoDSToStep;

fields

    myResult : TopologicalRepresentationItem from StepShape;

    myError  : MakeFaceError from TopoDSToStep;
    
end MakeStepFace;


