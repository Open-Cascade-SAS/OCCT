-- Created on: 2000-05-30
-- Created by: Sergey MOZOKHIN
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package XSDRAWSTLVRML

	---Purpose:

uses Draw, MeshVS, StlMesh, TColStd, TCollection, Standard, TopoDS

is

    class DataSource;

    class DrawableMesh;

    class ElemNodesMap instantiates DataMap from TCollection
            ( Integer from Standard, DataMapOfIntegerInteger from TColStd, MapIntegerHasher from TColStd );

    class CoordsMap instantiates DataMap from TCollection
            ( Integer from Standard, DataMapOfIntegerReal from TColStd, MapIntegerHasher from TColStd );

    class ToVRML;
    ---Purpose: A utility which writes a Shape to VRML format

    InitCommands (theCommands : in out Interpretor from Draw);
    ---Purpose : Inits commands for writing to STL and VRML formats

    Factory (theDI : out Interpretor from Draw);
    ---Purpose: Loads all Draw commands of TKXSDRAW. Used for plugin.

end XSDRAWSTLVRML;
