-- Created on: 1994-09-19
-- Created by: Gilles DEBARBOUILLE
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



generic class Node from Dynamic (Item as Transient)

	---Purpose: This generic class    is a light  way  to  store a
	--          persistent   homogeneous  collection  of   objects
	--          inside another persistent object.

inherits

    TShared from MMgt
    

is

    Create returns mutable Node from Dynamic;
    
    ---Level: Advanced 
    
    ---Purpose: Returns an empty instance of this class.

    Create(anitem : any Item) returns mutable Node from Dynamic;
    
    ---Level: Advanced 
    
    ---Purpose: Returns an instance  of  this class  initialized  with
    --          <anitem> as object.

    Object(me : mutable ; anitem : any Item)
    
    ---Level: Advanced 
    
    ---Purpose: Sets to <me> the object <anitem>.
    
    is static;
    
    Object(me) returns any Item
    
    ---Level: Advanced 
    
    ---Purpose: Returns the object into <me>.
    
    is static;
    
    Next(me : mutable ; anode : Node from Dynamic)
    
    ---Level: Advanced 
    
    ---Purpose: Links to <me> the node <anode>.
    
    is static;
    
    Next(me) returns any Node from Dynamic
    
    ---Level: Advanced 
    
    ---Purpose: Returns the node linked to <me>.
    
    is static;
    
fields

    thenextnode : Node from Dynamic;
    theitem     : Item;

end Node;



