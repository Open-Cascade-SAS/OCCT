-- Created on: 1997-02-12
-- Created by: Alexander BRIVIN
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class PointLight from Vrml 

	---Purpose:defines a point  light node of VRML specifying
	--         properties of lights. 
    	--  This  node  defines  a  point  light  source   at  a  fixed  3D  location
    	--  A  point  source  illuminates equally  in  all  directions;   
    	--  that  is  omni-directional.
    	--  Color is  written  as  an  RGB  triple.
    	--  Light intensity must be in the range 0.0 to 1.0, inclusive.  

uses
 
    Color   from Quantity, 
    Vec     from gp

is
                                                    --  defaults  :
    Create returns PointLight from Vrml; 
    	    	    	    	    	    	    --  myOnOff(Standard_TRUE)
 						    --  myIntensity(1)
						    --  myColor(1 1 1)
						    --  myLocation(0 0 1)

    Create  (  aOnOff     :   Boolean from  Standard; 
    	       aIntensity :   Real    from  Standard; 
    	       aColor     :   Color   from  Quantity; 
    	       aLocation  :   Vec     from  gp ) 
    	returns PointLight from Vrml; 
     
    SetOnOff ( me : in out;  aOnOff : Boolean from  Standard );
    OnOff ( me )  returns Boolean  from  Standard;

    SetIntensity ( me : in out;  aIntensity : Real from  Standard );
    Intensity ( me )  returns Real  from  Standard;

    SetColor ( me : in out;  aColor :  Color   from  Quantity );
    Color ( me )  returns  Color   from  Quantity;

    SetLocation ( me : in out;  aLocation : Vec  from  gp );
    Location ( me )  returns Vec  from  gp;

    Print  ( me;  anOStream: in out OStream from Standard) returns OStream from Standard;
    ---C++:  return  & 

fields
 
    myOnOff     :   Boolean from  Standard; -- Whether light is on
    myIntensity :   Real    from  Standard; -- Source intensity (0 to 1)
    myColor     :   Color   from  Quantity; -- RGB source color
    myLocation  :   Vec     from  gp;       -- Illumination Location vector

end PointLight;

