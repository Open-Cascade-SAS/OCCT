-- Created on: 1993-05-26
-- Created by: Laurent BOURESCHE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



deferred generic class Tool from Sweep (TheShape as any)

    ---Purpose: This  is a signature  class  describing the indexation
    --          and type analysis  services required by  the Directing
    --          and Generating Shapes of Swept Primitives.
    --          

uses

    ShapeEnum from TopAbs,
    Orientation from TopAbs

raises 

    OutOfRange from Standard

is

    Initialize(aShape: TheShape);
	---Purpose: Initialize the tool  with <aShape>.  The IndexTool
	--          must prepare an indexation for  all  the subshapes
	--          of this shape.

    NbShapes(me) returns Integer
	---Purpose: Returns the number of subshapes in the shape.
    is deferred;

    Index(me; aShape : TheShape) returns Integer
	---Purpose: Returns the index of <aShape>.
    is deferred;
    
    Shape(me; anIndex : Integer from Standard) returns TheShape
	---Purpose: Returns the Shape of index anIndex
    is deferred;
    
    Type(me; aShape : TheShape) returns ShapeEnum from TopAbs
	---Purpose: Returns the type of <aShape>.
    is deferred;
    
    Orientation(me; aShape : TheShape) returns Orientation from TopAbs
	---Purpose: Returns the Orientation of <aShape>.
    is deferred;
    
    SetOrientation(me; aShape : in out TheShape; Or : Orientation from TopAbs) 
	---Purpose: Set the Orientation of <aShape> with Or.
    is deferred;

------------------------------------------
--- Methods used for Directing Shapes only
------------------------------------------

    HasFirstVertex(me) returns Boolean from Standard
	---Purpose: Returns true if there is a First Vertex in the Shape.
    is deferred;

    HasLastVertex(me) returns Boolean from Standard
	---Purpose: Returns true if there is a Last Vertex in the Shape.
    is deferred;

    FirstVertex(me) returns TheShape
	---Purpose: Returns the first vertex.
    is deferred;

    LastVertex(me) returns TheShape
	---Purpose: Returns the last vertex.
    is deferred;

end Tool from Sweep;
