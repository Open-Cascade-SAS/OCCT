-- File:	RWStepFEA_RWNodeDefinition.cdl
-- Created:	Sun Dec 15 10:59:25 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWNodeDefinition from RWStepFEA

    ---Purpose: Read & Write tool for NodeDefinition

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    NodeDefinition from StepFEA

is
    Create returns RWNodeDefinition from RWStepFEA;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : NodeDefinition from StepFEA);
	---Purpose: Reads NodeDefinition

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: NodeDefinition from StepFEA);
	---Purpose: Writes NodeDefinition

    Share (me; ent : NodeDefinition from StepFEA;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWNodeDefinition;
