-- Created on: 1992-10-08
-- Created by: Isabelle GRIGNON
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package GeomAdaptor 

	---Purpose: this package contains the  geometric definition of
	--          curve and surface necessary to use algorithmes.

uses 
    Geom,
    GeomAbs,
    Adaptor3d,
    gp,
    Standard,
    TColStd,
    Geom2dAdaptor,
    TColgp,
    Precision

is
      class Curve; 

      class Surface;

      private class GHSurface instantiates GenHSurface from Adaptor3d
      	    (Surface from GeomAdaptor);
	    
      class HSurface;

      private class GHCurve instantiates GenHCurve from Adaptor3d
            (Curve from GeomAdaptor);
      
      class HCurve;
	---Purpose: Inherited  from    GHCurve.   Provides a  curve
	--          handled by reference.

    
      MakeCurve( C : Curve from Adaptor3d)
	---Purpose: Build a Geom_Curve using the informations from the 
	--          Curve from Adaptor3d
      returns Curve from Geom;
      
      MakeSurface( S : Surface from Adaptor3d)
	---Purpose: Build a Geom_Surface using the informations from the 
	--          Surface from Adaptor3d
      returns Surface from Geom;
      
end GeomAdaptor;
