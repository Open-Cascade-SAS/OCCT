-- File:	StepBasic_DocumentRepresentationType.cdl
-- Created:	Wed May 10 15:09:06 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class DocumentRepresentationType from StepBasic
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity DocumentRepresentationType

uses
    HAsciiString from TCollection,
    Document from StepBasic

is
    Create returns DocumentRepresentationType from StepBasic;
	---Purpose: Empty constructor

    Init (me: mutable; aName: HAsciiString from TCollection;
                       aRepresentedDocument: Document from StepBasic);
	---Purpose: Initialize all fields (own and inherited)

    Name (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Name
    SetName (me: mutable; Name: HAsciiString from TCollection);
	---Purpose: Set field Name

    RepresentedDocument (me) returns Document from StepBasic;
	---Purpose: Returns field RepresentedDocument
    SetRepresentedDocument (me: mutable; RepresentedDocument: Document from StepBasic);
	---Purpose: Set field RepresentedDocument

fields
    theName: HAsciiString from TCollection;
    theRepresentedDocument: Document from StepBasic;

end DocumentRepresentationType;
