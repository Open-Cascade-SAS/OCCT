-- Created on: 1993-10-26
-- Created by: Christian CAILLET
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class FileProtocol  from IGESData    inherits  Protocol  from IGESData

    ---Purpose : This class allows to define complex protocols, in order to
    --           treat various sub-sets (or the complete set) of the IGES Norm,
    --           such as Solid + Draw (which are normally independant), etc...
    --           While it inherits Protocol from IGESData, it admits
    --           UndefinedEntity too

uses Protocol from Interface

is

    Create returns mutable FileProtocol;
    ---Purpose : Returns an empty FileProtocol

    Add (me : mutable; protocol : Protocol from IGESData);
    ---Purpose : Adds a resource

    NbResources (me) returns Integer  is redefined;
    ---Purpose : Gives the count of Resources : the count of Added Protocols

    Resource (me; num : Integer) returns Protocol from Interface  is redefined;
    ---Purpose : Returns a Resource, given a rank (rank of call to Add)

fields

    theresource : Protocol from IGESData;
    thenext     : FileProtocol from IGESData;

end FileProtocol;
