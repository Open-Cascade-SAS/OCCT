-- Created by: NW,JPB,CAL
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package Aspect

        ---Version:

        ---Purpose: This package contains the group of graphic elements common
        --          to different types of visualisers. It allows the description
        --          of a screen background, a window, an edge, and groups of
        --          graphic attributes that can be used in describing 2D
        --          and 3D objects.

        ---Keywords: Window, Aspect, FillArea, Line, Marker, Edge
        --           Highlight, Hatch, Background, GradientBackground, Color map,
        --           Type map, Width map, Font map
        ---Warning:
        ---References:

uses
        TCollection,
        TColStd,
        TShort,
        Quantity,
        TColQuantity,
        Resource,
        MMgt

is
        ---------------------------
        -- Category: Imported types
        ---------------------------
        imported FStream;
        -- waiting for RBA creating this class in Standard ...  

        imported IFStream;
        -- G002A study 

        imported CLayer2d;

        ---Category: Imported types

        primitive Handle;
        primitive Drawable;

        primitive Display;

        primitive RenderingContext;

        imported GraphicCallbackProc;

        -- 22-03-04 OCC4895 SAN High-level interface for controlling polygon offsets
        imported PolygonOffsetMode;

        -----------------------
        -- Category: Exceptions
        -----------------------

        exception AspectLineDefinitionError inherits OutOfRange;
        ---Category: Exceptions

        exception AspectFillAreaDefinitionError inherits OutOfRange;
        ---Category: Exceptions

        exception AspectMarkerDefinitionError inherits OutOfRange;
        ---Category: Exceptions

        exception BadAccess inherits DomainError;
        ---Category: Exceptions

        exception IdentDefinitionError inherits OutOfRange;
        ---Category: Exceptions

        exception WindowDefinitionError inherits OutOfRange;
        ---Category: The exceptions

        exception WindowError inherits OutOfRange;
        ---Category: The exceptions

        exception DriverDefinitionError inherits OutOfRange;
        ---Category: The exceptions

        exception GraphicDeviceDefinitionError inherits OutOfRange;
        ---Category: The exceptions

        exception DisplayConnectionDefinitionError inherits OutOfRange;
        ---Category: The exceptions

        ---------------------------
        -- Category: Classes Aspect
        ---------------------------

        deferred class AspectLine;
        ---Category: Classes Aspect

        deferred class AspectMarker;
        ---Category: Classes Aspect

        deferred class AspectFillArea;
        ---Category: Classes Aspect

        --------------------
        -- Category: Classes
        --------------------

        class Background;
        ---Category: Classes

        class GradientBackground;
        ---Category: Classes

        class GenId;
        ---Category: Classes

        deferred class Window;
        ---Category: Classes

        deferred class Grid;
        class RectangularGrid;
        class CircularGrid;

        deferred class ColorScale;

        imported DisplayConnection;

        imported DisplayConnection_Handle;

        -------------------------
        -- Category: Enumerations
        -------------------------

        enumeration HatchStyle is       HS_HORIZONTAL,
                                        HS_HORIZONTAL_WIDE,
                                        HS_VERTICAL,
                                        HS_VERTICAL_WIDE,
                                        HS_DIAGONAL_45,
                                        HS_DIAGONAL_45_WIDE,
                                        HS_DIAGONAL_135,
                                        HS_DIAGONAL_135_WIDE,
                                        HS_GRID,
                                        HS_GRID_WIDE,
                                        HS_GRID_DIAGONAL,
                                        HS_GRID_DIAGONAL_WIDE
        end HatchStyle;
        ---Purpose: Definition of all available hatch styles.
        --
        --          HS_HORIZONTAL
        --          HS_HORIZONTAL_WIDE
        --          HS_VERTICAL
        --          HS_VERTICAL_WIDE
        --          HS_DIAGONAL_45
        --          HS_DIAGONAL_45_WIDE
        --          HS_DIAGONAL_135
        --          HS_DIAGONAL_135_WIDE
        --          HS_GRID
        --          HS_GRID_WIDE
        --          HS_GRID_DIAGONAL
        --          HS_GRID_DIAGONAL_WIDE
        --
        ---Category: Enumerations

        enumeration InteriorStyle is    IS_EMPTY,
                                        IS_HOLLOW,
                                        IS_HATCH,
                                        IS_SOLID,
                                        IS_HIDDENLINE,
                                        IS_POINT
        end InteriorStyle;
        ---Purpose: Definition of interior types for primitive
        --          faces.
        --
        --          IS_EMPTY    no interior.
        --          IS_HOLLOW   display the boundaries of the surface.
        --          IS_HATCH    display hatched with a hatch style.
        --          IS_SOLID    display the interior entirely filled.
        --          IS_HIDDENLINE       display in hidden lines removed.
        --          IS_POINT            display only vertices.
        --
        ---Category: Enumerations

        enumeration TypeOfConstraint is TOC_BOTTOM_LEFT,
                                        TOC_BOTTOM_RIGHT,
                                        TOC_TOP_LEFT, 
                                        TOC_TOP_RIGHT
        end TypeOfConstraint;
        ---Purpose: Definition of the attachment for the layers
        --
        ---Category: Enumerations

        enumeration TypeOfDrawMode is   TODM_REPLACE,
                                        TODM_ERASE,
                                        TODM_XOR,
                                        TODM_XORLIGHT
        end TypeOfDrawMode;
        ---Purpose: Definition of the draw modes
        --
        ---Category: Enumerations

        enumeration TypeOfEdge is       TOE_VISIBLE,
                                        TOE_INVISIBLE
        end TypeOfEdge;
        ---Purpose: Definition of edge visibility
        --
        --          TOE_VISIBLE         Edge is displayed
        --          TOE_INVISIBLE       Edge is not displayed
        --
        ---Category: Enumerations

        enumeration TypeOfHighlightMethod is    TOHM_COLOR,
                                                TOHM_BOUNDBOX
        end TypeOfHighlightMethod;
        ---Purpose: Definition of a highlight method
        --
        --          TOHM_COLOR          drawn in the highlight color
        --                              (default white)
        --          TOHM_BOUNDBOX       enclosed by the boundary box
        --                              (default white)
        --
        ---Category: Enumerations

        enumeration TypeOfLine is       TOL_SOLID,
                                        TOL_DASH,
                                        TOL_DOT,
                                        TOL_DOTDASH,
                                        TOL_USERDEFINED
        end TypeOfLine;
        ---Purpose: Definition of line types
        --
        --          TOL_SOLID           continuous
        --          TOL_DASH            dashed 2.0,1.0 (MM)
        --          TOL_DOT             dotted 0.2,0.5 (MM)
        --          TOL_DOTDASH         mixed  10.0,1.0,2.0,1.0 (MM)
        --          TOL_USERDEFINED     defined by Users
        ---Category: Enumerations

        enumeration WidthOfLine is      WOL_THIN,
                                        WOL_MEDIUM,
                                        WOL_THICK,
                                        WOL_VERYTHICK,
                                        WOL_USERDEFINED
        end WidthOfLine;
        ---Purpose: Definition of line types
        --
        --          WOL_THIN            thin line (1 pixel width)
        --          WOL_MEDIUM          medium width of 0.5 MM
        --          WOL_THICK           thick width of 0.7 MM
        --          WOL_VERYTHICK       very thick width of 1.5 MM
        --          WOL_USERDEFINED     defined by Users
        ---Category: Enumerations

        enumeration TypeOfStyleText is  TOST_NORMAL,
                                        TOST_ANNOTATION
        end TypeOfStyleText;
        ---Purpose: Define the style of the text.       
        --
        --          TOST_NORMAL         Default text. The text is displayed like any other graphic object.
        --                              This text can be hidden by another object that is nearest from the 
        --                              point of view. 
        --          TOST_ANNOTATION     The text is always visible. The texte is displayed 
        --                              over the other object according to the priority.
        ---Category: Enumerations

        enumeration TypeOfDisplayText is        TODT_NORMAL,
                                                TODT_SUBTITLE,
                                                TODT_DEKALE,
                                                TODT_BLEND,
                                                TODT_DIMENSION
        end TypeOfDisplayText;
        ---Purpose: Define the display type of the text.        
        --
        --          TODT_NORMAL         Default display. Text only.     
        --          TODT_SUBTITLE       There is a subtitle under the text.
        --          TODT_DEKALE         The text is displayed with a 3D style.
        --          TODT_BLEND          The text is displayed in XOR.
        --          TODT_DIMENSION      Dimension line under text will be invisible. 
        ---Category: Enumerations

        enumeration TypeOfMarker is     TOM_POINT,
                                        TOM_PLUS,
                                        TOM_STAR,
                                        TOM_X,
                                        TOM_O,
                                        TOM_O_POINT,
                                        TOM_O_PLUS,
                                        TOM_O_STAR,
                                        TOM_O_X,
                                        TOM_RING1,
                                        TOM_RING2,
                                        TOM_RING3,
                                        TOM_BALL,
                                        TOM_USERDEFINED 
        end TypeOfMarker;
        ---Purpose: Definition of types of markers
        --
        --          TOM_POINT   point   .
        --          TOM_PLUS    plus    +
        --          TOM_STAR    star    *
        --          TOM_X       cross   x
        --          TOM_O       circle  O
        --          TOM_O_POINT a point in a circle
        --          TOM_O_PLUS  a plus in a circle
        --          TOM_O_STAR  a star in a circle
        --          TOM_O_X     a cross in a circle
        --          TOM_RING1   a large ring
        --          TOM_RING2   a medium ring
        --          TOM_RING3   a small ring
        --          TOM_BALL    a ball with 1 color and different saturations
        --          TOM_USERDEFINED     defined by Users
        --
        ---Category: Enumerations

        enumeration TypeOfUpdate is     TOU_ASAP,
                                        TOU_WAIT
        end TypeOfUpdate;
        ---Purpose: Definition of screen refresh mode
        --
        --          TOU_ASAP    as soon as possible
        --          TOU_WAIT    on demand (Update)
        --
        ---Category: Enumerations

        enumeration TypeOfDeflection is TOD_RELATIVE,
                                        TOD_ABSOLUTE
        end TypeOfDeflection;
        ---Purpose: Defines if the maximal chordial deflection used when
        --          drawing an object is absolute  or relative to the size 
        --          of the object.

        enumeration TypeOfResize is     TOR_UNKNOWN,
                                        TOR_NO_BORDER,
                                        TOR_TOP_BORDER,
                                        TOR_RIGHT_BORDER,
                                        TOR_BOTTOM_BORDER,
                                        TOR_LEFT_BORDER,
                                        TOR_TOP_AND_RIGHT_BORDER,
                                        TOR_RIGHT_AND_BOTTOM_BORDER,
                                        TOR_BOTTOM_AND_LEFT_BORDER,
                                        TOR_LEFT_AND_TOP_BORDER
        end TypeOfResize;
        ---Purpose: Defines the type of Resize Window method applied
        --          by the user.

        enumeration TypeOfPrimitive is
                                        TOP_UNKNOWN,
                                        TOP_POLYLINE,
                                        TOP_POLYGON,
                                        TOP_SEGMENTS,
                                        TOP_ARCS,
                                        TOP_POLYARCS,
                                        TOP_POINTS,
                                        TOP_MARKERS
        end TypeOfPrimitive;
        ---Purpose:

        enumeration GridDrawMode is GDM_Lines,
                                    GDM_Points,
                                    GDM_None
        end GridDrawMode;
        ---Purpose: Defines the grid draw mode. The grid may be drawn
        --          by using lines or points.

        enumeration GridType is GT_Rectangular,
                                GT_Circular
        end GridType;
        ---Purpose: Defines the grid type : Rectangular or Circular.

        enumeration TypeOfTriedronEcho is       TOTE_NONE,
                                                TOTE_ORIGIN,
                                                TOTE_AXIS_X,
                                                TOTE_AXIS_Y,
                                                TOTE_AXIS_Z,
                                                TOTE_TEXT_X,
                                                TOTE_TEXT_Y,
                                                TOTE_TEXT_Z, 
                                                TOTE_01,
                                                TOTE_02,
                                                TOTE_03,
                                                TOTE_04,
                                                TOTE_05,
                                                TOTE_06,
                                                TOTE_07,
                                                TOTE_08,
                                                TOTE_09,
                                                TOTE_10
        end TypeOfTriedronEcho;
        ---Purpose: Definition of the Triedron echo zone to highlight
        --
        --          TOTE_NONE           no echo zone
        --          TOTE_ORIGIN         a box on origin of the Triedron
        --          TOTE_AXIS_X         highlights the X axis
        --          TOTE_AXIS_Y         highlights the Y axis
        --          TOTE_AXIS_Z         highlights the Z axis
        --          TOTE_TEXT_X         highlights the X character
        --          TOTE_TEXT_Y         highlights the Y character
        --          TOTE_TEXT_Z         highlights the Z character
        --          TOTE_01 to TOTE_10  not yet implemented.
        ---Category: The enumerations


        enumeration TypeOfTriedronPosition is   TOTP_CENTER,
                                                TOTP_LEFT_LOWER,
                                                TOTP_LEFT_UPPER,
                                                TOTP_RIGHT_LOWER,
                                                TOTP_RIGHT_UPPER,
                                                TOTP_01,
                                                TOTP_02,
                                                TOTP_03,
                                                TOTP_04,
                                                TOTP_05,
                                                TOTP_06,
                                                TOTP_07,
                                                TOTP_08,
                                                TOTP_09,
                                                TOTP_10
        end TypeOfTriedronPosition;
        ---Purpose: Definition of the Triedron position in the views
        --
        --          TOTP_CENTER         at the center of the view
        --          TOTP_LEFT_LOWER     at the left lower corner
        --          TOTP_LEFT_UPPER     at the left upper corner
        --          TOTP_RIGHT_LOWER    at the right lower corner
        --          TOTP_RIGHT_UPPER    at the right upper corner
        --          TOTP_01 to TOTP_10  not yet implemented.
        ---Category: The enumerations

        enumeration TypeOfLayer is      TOL_OVERLAY, 
                                        TOL_UNDERLAY
        end TypeOfLayer;
        ---Purpose: Modes of drawing for the objects in a layer
        --
        --          TOL_OVERLAY, the graphic of the layer is draw
        --                       after the 3d graphic.
        --          TOL_UNDERLAY, the graphic of the layer is draw
        --                       before the 3d graphic.
        ---Category: The enumerations

        enumeration TypeOfFacingModel is TOFM_BOTH_SIDE,
                                         TOFM_BACK_SIDE,
                                         TOFM_FRONT_SIDE
        end TypeOfFacingModel;

        enumeration FillMethod is
          FM_NONE,
          FM_CENTERED,
          FM_TILED,
          FM_STRETCH
        end FillMethod;
        ---Purpose: Defines the fill methods to
        --      write bitmaps in a window.

        enumeration GradientFillMethod is
          GFM_NONE,
          GFM_HOR,
          GFM_VER,
          GFM_DIAG1,
          GFM_DIAG2,
          GFM_CORNER1,
          GFM_CORNER2,
          GFM_CORNER3,
          GFM_CORNER4
        end GradientFillMethod;
        ---Purpose: Defines the fill methods to
        --      write gradient background in a window.

        enumeration TypeOfColorScaleData is
          TOCSD_AUTO,
          TOCSD_USER
        end TypeOfColorScaleData;
        ---Purpose: Defines the using type of colors and labels

        enumeration TypeOfColorScalePosition is
          TOCSP_NONE,
          TOCSP_LEFT,
          TOCSP_RIGHT,
          TOCSP_CENTER
        end TypeOfColorScalePosition;
        ---Purpose: Defines the type of position for color scale labels

        enumeration TypeOfColorScaleOrientation is
          TOCSO_NONE,
          TOCSO_LEFT,
          TOCSO_RIGHT,
          TOCSO_CENTER
        end TypeOfColorScaleOrientation;
        ---Purpose: Defines the type of color scale orientation

        enumeration PrintAlgo is
          PA_STRETCH,
          PA_TILE
        end PrintAlgo;
        ---Purpose: Defines print algorithm
        --          Aspect_PrintAlgo:
        --          1) PA_STRETCH - Stretch offscreen printing frame
        --                          if its dimensions are smaller than
        --                          the printer's printing area dimensions;
        --                          This algorithm is more reliable as it
        --                          works on any hardware and is recommended
        --                          to be used with average printing resolutions,
        --                          as it more RAM memory dependent than PA_TILE;
        --                          Stretching is performend using bicubic interpolation
        --                          algorithm from FreeImage library if OCCT is built
        --                          with FreeImage support, otherwise Windows API 
        --                          StretchBlt() function in STRETCH_HALFTONE mode
        --                          is used;
        --          2) PA_TILE    - If the offscreen printing frame dimensions
        --                          are smaller than the printer's printing
        --                          area dimensions - use multiple printing
        --                          frames to cover the whole printing area
        enumeration XAtom is
          XA_DELETE_WINDOW
        end XAtom;
        ---Purpose: Defines custom identifiers(atoms) for X window custom named properties
        ---------------------------------
        -- Category: Instantiated classes
        ---------------------------------

        class SequenceOfColor instantiates
                Sequence from TCollection(Color from Quantity);

end Aspect;
