-- Created on: 1996-01-09
-- Created by: Laurent PAINNOT
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


private class FuncExtSS from Extrema

 inherits FunctionSetWithDerivatives from math
    ---Purpose: Function to find extrema of the 
    --          distance between two surfaces.

uses    POnSurf           from Extrema,
	SequenceOfPOnSurf from Extrema,
	SequenceOfReal    from TColStd,
	Pnt               from gp,
	Vector            from math,
	Matrix            from math,
	Surface           from Adaptor3d,
    	SurfacePtr        from Adaptor3d

raises  OutOfRange from Standard

is
    Create returns FuncExtSS;

    Create (S1, S2: Surface from Adaptor3d) returns FuncExtSS;
    	---Purpose:

    Initialize(me: in out; S1, S2: Surface from Adaptor3d)
    	---Purpose: sets the field mysurf of the function.
    is static;
    
    ------------------------------------------------------------
    -- In all next methods, an exception is raised if the fields 
    -- were not initialized.

    NbVariables (me) returns Integer;

    NbEquations (me) returns Integer;

    Value (me: in out; UV: Vector; F: out Vector) returns Boolean;
    	---Purpose: Calculate Fi(U,V).

    Derivatives (me: in out; UV: Vector; DF: out Matrix)
    	returns Boolean;
    	---Purpose: Calculate Fi'(U,V).

    Values (me: in out; UV: Vector; F: out Vector; DF: out Matrix)
    	returns Boolean;
    	---Purpose: Calculate Fi(U,V) and Fi'(U,V).

    GetStateNumber (me: in out) returns Integer
    	---Purpose: Save the found extremum.
    	is redefined;

    NbExt (me) returns Integer;
    	---Purpose: Return the number of found extrema.

    SquareDistance (me; N: Integer) returns Real
    	---Purpose: Return the value of the Nth distance.
    	raises  OutOfRange;
	    	-- if N < 1 or N > NbExt(me).

    PointOnS1 (me; N: Integer) returns POnSurf
    	---Purpose: Return the Nth extremum on S1.
    	raises  OutOfRange;
	    	-- if N < 1 or N > NbExt(me).

    PointOnS2 (me; N: Integer) returns POnSurf
    	---Purpose: Renvoie le Nieme extremum sur S2.
    	raises  OutOfRange;
	    	-- si N < 1 ou N > NbExt(me).

    Bidon(me) returns SurfacePtr from Adaptor3d
    is static private;


fields
    myS1   : SurfacePtr from Adaptor3d;
    myS2   : SurfacePtr from Adaptor3d;
    
    myP1   : Pnt from gp;
    myP2   : Pnt from gp;

    myU1    : Real;          -- current value of U on S1
    myV1    : Real;          -- current value of V on S1
    myU2    : Real;          -- current value of U on S2
    myV2    : Real;          -- current value of V on S2

    mySqDist:  SequenceOfReal    from TColStd;
    myPoint1: SequenceOfPOnSurf from Extrema;
    myPoint2: SequenceOfPOnSurf from Extrema;
    
    myS1init: Boolean;
    myS2init: Boolean;

end FuncExtSS;
