-- Created on: 1997-02-12
-- Created by: Alexander BRIVIN
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class WWWInline from Vrml 

	---Purpose: defines a WWWInline node of VRML specifying group properties.
    	--  The  WWWInline  group  node  reads  its  children  from  anywhere  in  the   
    	--  World  Wide  Web.
	--  Exactly  when  its  children  are  read  is  not  defined; 
	--  reading  the  children  may  be  delayed  until  the  WWWInline  is  actually 
    	--  displayed. 
	--  WWWInline  with  an  empty  ("")  name  does  nothing. 
	--  WWWInline  behaves  like  a  Separator,  pushing  the  traversal  state 
	--  before  traversing  its  children  and  popping  it  afterwards.
    	--  By  defaults: 
	--    myName  ("")
	--    myBboxSize (0,0,0)
	--    myBboxCenter  (0,0,0)

uses
 
    AsciiString   from   TCollection,
    Vec           from   gp 

is
 
    Create returns  WWWInline from Vrml; 

    Create  ( aName        :   AsciiString from  TCollection; 
    	      aBboxSize    :   Vec         from  gp;
    	      aBboxCenter  :   Vec         from  gp )
    	returns  WWWInline from Vrml; 

    SetName ( me : in out; aName : AsciiString from TCollection );
    Name ( me )  returns  AsciiString from TCollection;

    SetBboxSize ( me : in out; aBboxSize  : Vec  from  gp);
    BboxSize ( me )  returns   Vec  from  gp;

    SetBboxCenter ( me : in out; aBboxCenter  : Vec  from  gp);
    BboxCenter ( me )  returns  Vec  from  gp;

    Print  ( me;  anOStream: in out OStream from Standard) returns OStream from Standard;
    ---C++:  return  & 

fields
 
    myName        :   AsciiString from TCollection;   -- URL name
    myBboxSize    :   Vec         from gp;            -- Size of 3D bounding box
    myBboxCenter  :   Vec         from gp;            -- Center of 3D bounding box
    
end WWWInline;

