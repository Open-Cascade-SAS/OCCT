-- Created by: Peter KURNEV
-- Copyright (c) 2010-2014 OPEN CASCADE SAS
-- Copyright (c) 2007-2010 CEA/DEN, EDF R&D, OPEN CASCADE
-- Copyright (c) 2003-2007 OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN, CEDRAT,
--                         EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PassKey from BOPDS 

	---Purpose: 
	--  The class BOPDS_PassKey is to provide 
        --  possibility to map objects that  
    	--  have a set of integer IDs as a base        

uses
    Shape from TopoDS, 
    ListOfInteger from BOPCol,
    PInteger from BOPCol, 
    BaseAllocator from BOPCol

--raises

is 
    Create  
    	returns PassKey from BOPDS; 
    ---C++: inline 
    ---C++: alias "virtual ~BOPDS_PassKey();" 
    	---Purpose:  
    	--- Empty contructor  
    	---   
	 
    Create (theAllocator: BaseAllocator from BOPCol)  
    	returns PassKey from BOPDS;  
    ---C++: inline 
	---Purpose:  
    	---  Contructor    
    	---  theAllocator - the allocator to manage the memory     
    	---  
	      
    Create(Other:PassKey from BOPDS) 
    	returns PassKey from BOPDS; 
    ---C++: inline    
    ---C++: alias "BOPDS_PassKey& operator =(const BOPDS_PassKey& Other);" 
    	---Purpose:  
    	---  Copy Contructor 
	 
    Clear(me:out); 
    ---C++: inline  
    	---Purpose:  
    	---  Clear the contents 
	 
    SetIds(me:out; 
    	    theI1  :Integer from Standard); 
    ---C++: inline      
     	---Purpose: 
	--- Modifier 
	--- Sets one Id <theI1>   
	
    SetIds(me:out; 
    	    theI1 :Integer from Standard; 
    	    theI2 :Integer from Standard);  
    ---C++: inline      
     	---Purpose: 
	--- Modifier 
	--- Sets two Id <theI1>,<theI2>    
	
    SetIds(me:out; 
    	    theI1 :Integer from Standard;    
    	    theI2 :Integer from Standard;    
    	    theI3 :Integer from Standard);  
    ---C++: inline  
    	---Purpose: 
	--- Modifier 
	--- Sets three Id <theI1>,<theI2>,<theI3>    
    SetIds(me:out; 
    	    theI1 :Integer from Standard;    
    	    theI2 :Integer from Standard;    
    	    theI3 :Integer from Standard;    
    	    theI4 :Integer from Standard); 
    ---C++: inline  
    	---Purpose: 
	--- Modifier 
	--- Sets four Id <theI1>,<theI2>,<theI3>,<theI4>    
    SetIds(me:out; 
    	    theLI:ListOfInteger from BOPCol); 
	---Purpose: 
	--- Modifier 
	--- Sets the list of Id <theLI> 

    NbIds(me) 
	returns Integer  from Standard; 
    ---C++: inline  
    	---Purpose: 
	--- Selector
	--- Returns the number of Ids> 
     
    IsEqual(me; 
    	    theOther:PassKey from BOPDS) 
	returns Boolean from Standard;   		     
    ---C++: inline 
     	---Purpose: 
	--- Query
	--- Returns true if the PassKey is equal to <the theOther> 

    HashCode(me; 
	    theUpper : Integer  from Standard)  
    	returns Integer from Standard;   	 
    ---C++: inline	 
    	---Purpose: 
	--- Query
	--- Returns hash  code 
 
    Id(me; 
    	    theIndex: Integer  from Standard)  
    	returns  Integer from Standard;
    ---C++: inline  
    	---Purpose: 
	--- Selector
	--- Returns Id of index <theIndex>  
     
    Ids(me; 
    	    theI1 :out Integer from Standard;    
    	    theI2 :out Integer from Standard);
    ---C++: inline 
    	---Purpose:  
    	--- Selector
	--- Returns the first two Ids <theI1>,<theI2> 
	
    Dump(me; 
    	aHex:Integer from Standard=0);
     
    Allocate(me:out; 
    	    theSize:Integer from Standard) 
    	returns PInteger from BOPCol 
    	is protected; 
    ---C++: inline
	
fields  
    myAllocator : BaseAllocator from BOPCol is protected;
    myNbIds: Integer from Standard is protected;  
    mySum  : Integer from Standard is protected;  
    myPtr  : PInteger from BOPCol is protected;  
     
end PassKey;
