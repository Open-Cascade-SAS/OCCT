-- File:	StepToGeom_MakeTransformation3d.cdl
-- Created:	Tue Feb 16 11:14:36 1999
-- Author:	Andrey BETENEV
---Copyright:	 Matra Datavision 1999

class MakeTransformation3d from StepToGeom

    ---Purpose: Convert cartesian_transformation_operator_3d to gp_Trsf

uses
    CartesianTransformationOperator3d from StepGeom,
    Trsf from gp

is

    Convert ( myclass; SCTO : CartesianTransformationOperator3d from StepGeom;
                       CT : out Trsf from gp )
    returns Boolean from Standard;

end MakeTransformation3d;
