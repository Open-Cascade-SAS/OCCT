-- Created on: 1993-07-06
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MakeEdge from BRepBuilderAPI  inherits MakeShape from BRepBuilderAPI

	---Purpose: Provides methods to build edges.
	--          
	--          The   methods have  the  following   syntax, where
	--          TheCurve is one of Lin, Circ, ...
	--          
	--          Create(C : TheCurve)
	--            
	--            Makes an edge on  the whole curve.  Add vertices
	--            on finite curves.
	--            
	--          Create(C : TheCurve; p1,p2 : Real)
	--          
	--            Make an edge  on the curve between parameters p1
	--            and p2. if p2 < p1 the edge will be REVERSED. If
	--            p1  or p2 is infinite the  curve will be open in
	--            that  direction. Vertices are created for finite
	--            values of p1 and p2.
	--            
	--          Create(C : TheCurve; P1, P2 : Pnt from gp)
	--          
	--            Make an edge on the curve  between the points P1
	--            and P2. The  points are projected on   the curve
	--            and the   previous method is  used. An  error is
	--            raised if the points are not on the curve.
	--            
	--          Create(C : TheCurve; V1, V2 : Vertex from TopoDS)
	--          
	--            Make an edge  on the curve  between the vertices
	--            V1 and V2. Same as the  previous but no vertices
	--            are created. If a vertex is  Null the curve will
	--            be open in this direction.

uses
    EdgeError from BRepBuilderAPI,
    Edge      from TopoDS,
    Vertex    from TopoDS,
    Pnt       from gp,
    Lin       from gp,
    Circ      from gp,
    Elips     from gp,
    Hypr      from gp,
    Parab     from gp,
    Curve     from Geom2d,
    Curve     from Geom,
    Surface   from Geom,
    MakeEdge  from BRepLib
    
raises
    NotDone from StdFail
    
is

    Create returns MakeEdge from BRepBuilderAPI;

    ----------------------------------------
    -- Points
    ----------------------------------------

    Create(V1, V2 : Vertex from TopoDS)                    
	---Level: Public
    returns MakeEdge from BRepBuilderAPI;

    Create(P1, P2 : Pnt from gp)                           
	---Level: Public
    returns MakeEdge from BRepBuilderAPI;


    ----------------------------------------
    -- Lin
    ----------------------------------------
	
    Create(L : Lin from gp)                                
	---Level: Public
    returns MakeEdge from BRepBuilderAPI;

    Create(L : Lin from gp; p1,p2 : Real)                  
	---Level: Public
    returns MakeEdge from BRepBuilderAPI;

    Create(L : Lin from gp; P1,P2 : Pnt from gp)           
	---Level: Public
    returns MakeEdge from BRepBuilderAPI;

    Create(L : Lin from gp; V1, V2 : Vertex from TopoDS)   
	---Level: Public
    returns MakeEdge from BRepBuilderAPI;

    ----------------------------------------
    -- Circ
    ----------------------------------------
	
    Create(L : Circ from gp)                               
	---Level: Public
    returns MakeEdge from BRepBuilderAPI;

    Create(L : Circ from gp; p1,p2 : Real)                 
	---Level: Public
    returns MakeEdge from BRepBuilderAPI;

    Create(L : Circ from gp; P1,P2 : Pnt from gp)          
	---Level: Public
    returns MakeEdge from BRepBuilderAPI;

    Create(L : Circ from gp; V1, V2 : Vertex from TopoDS)  
	---Level: Public
    returns MakeEdge from BRepBuilderAPI;

	
    ----------------------------------------
    -- Elips
    ----------------------------------------

    Create(L : Elips from gp)                               
	---Level: Public
    returns MakeEdge from BRepBuilderAPI;

    Create(L : Elips from gp; p1,p2 : Real)                 
	---Level: Public
    returns MakeEdge from BRepBuilderAPI;

    Create(L : Elips from gp; P1,P2 : Pnt from gp)          
	---Level: Public
    returns MakeEdge from BRepBuilderAPI;

    Create(L : Elips from gp; V1, V2 : Vertex from TopoDS)  
	---Level: Public
    returns MakeEdge from BRepBuilderAPI;

    ----------------------------------------
    -- Hypr
    ----------------------------------------

    Create(L : Hypr from gp)                               
	---Level: Public
    returns MakeEdge from BRepBuilderAPI;

    Create(L : Hypr from gp; p1,p2 : Real)                 
	---Level: Public
    returns MakeEdge from BRepBuilderAPI;

    Create(L : Hypr from gp; P1,P2 : Pnt from gp)          
	---Level: Public
    returns MakeEdge from BRepBuilderAPI;

    Create(L : Hypr from gp; V1, V2 : Vertex from TopoDS)  
	---Level: Public
    returns MakeEdge from BRepBuilderAPI;

    ----------------------------------------
    -- Parab
    ----------------------------------------

    Create(L : Parab from gp)                               
	---Level: Public
    returns MakeEdge from BRepBuilderAPI;

    Create(L : Parab from gp; p1,p2 : Real)                 
	---Level: Public
    returns MakeEdge from BRepBuilderAPI;

    Create(L : Parab from gp; P1,P2 : Pnt from gp)          
	---Level: Public
    returns MakeEdge from BRepBuilderAPI;

    Create(L : Parab from gp; V1, V2 : Vertex from TopoDS)  
	---Level: Public
    returns MakeEdge from BRepBuilderAPI;

    ----------------------------------------
    -- Curve
    ----------------------------------------

    Create(L : Curve from Geom)                               
	---Level: Public
    returns MakeEdge from BRepBuilderAPI;

    Create(L : Curve from Geom; p1,p2 : Real)                 
	---Level: Public
    returns MakeEdge from BRepBuilderAPI;

    Create(L : Curve from Geom; 
    P1,P2 : Pnt from gp)
	---Level: Public                        
    returns MakeEdge from BRepBuilderAPI;

    Create(L : Curve from Geom; 
    V1, V2 : Vertex from TopoDS)
	---Level: Public
    returns MakeEdge from BRepBuilderAPI;

    Create(L : Curve from Geom; 
    P1,P2 : Pnt from gp; p1,p2 : Real)                        
	---Level: Public
    returns MakeEdge from BRepBuilderAPI;

    Create(L : Curve from Geom; 
    V1, V2 : Vertex from TopoDS;
    p1, p2 :Real)       
	---Level: Public                                      
    returns MakeEdge from BRepBuilderAPI;

    ----------------------------------------
    -- Curve and surface
    ----------------------------------------

    Create(L : Curve from Geom2d; S : Surface from Geom)
    	---Level: Public
    returns MakeEdge from BRepBuilderAPI;

    Create(L : Curve from Geom2d; S : Surface from Geom; p1,p2 : Real)
    	---Level: Public
    returns MakeEdge from BRepBuilderAPI;

    Create(L : Curve from Geom2d; S : Surface from Geom; 
    P1,P2 : Pnt from gp)
	---Level: Public                        
    returns MakeEdge from BRepBuilderAPI;

    Create(L : Curve from Geom2d; S : Surface from Geom; 
    V1, V2 : Vertex from TopoDS)
	---Level: Public
    returns MakeEdge from BRepBuilderAPI;

    Create(L : Curve from Geom2d; S : Surface from Geom; 
    P1,P2 : Pnt from gp; p1,p2 : Real)                        
	---Level: Public
    returns MakeEdge from BRepBuilderAPI;

    Create(L : Curve from Geom2d; S : Surface from Geom; 
    V1, V2 : Vertex from TopoDS;
    p1, p2 :Real)       
	---Level: Public                                      
    returns MakeEdge from BRepBuilderAPI;

 
    	---Purpose: The general method to directly create an edge is to give
    	-- -      a 3D curve C as the support (geometric domain) of the edge,
    	-- -      two vertices V1 and V2 to limit the curve (definition of the restriction of
    	--    the edge), and
    	-- -      two real values p1 and p2 which are the parameters for the vertices V1 and V2
    	--    on the curve.
    	-- The curve may be defined as a 2d curve in the parametric space of a surface: a
    	-- pcurve. The surface on which the edge is built is then kept at the level of the edge.
    	-- The default tolerance will be associated with this edge.
    	-- Rules applied to the arguments:
    	-- For the curve:
    	-- -      The curve must not be a 'null handle'.
    	-- -      If the curve is a trimmed curve the basis curve is used.
    	-- For the vertices:
    	-- -      Vertices may be null shapes. When V1 or V2 is null the edge is open in the
    	--    corresponding direction and the parameter value p1 or p2 must be infinite
    	--    (remember that Precision::Infinite() defines an infinite value).
    	-- -      The two vertices must be identical if they have the same 3D location.
    	--    Identical vertices are used in particular when the curve is closed.
    	-- For the parameters:
    	-- -      The parameters must be in the parametric range of the curve (or the basis
    	--    curve if the curve is trimmed). If this condition is not satisfied the edge is not
    	--    built, and the Error function will return BRepAPI_ParameterOutOfRange.
    	-- -      Parameter values must not be equal. If this condition is not satisfied (i.e.
    	--    if | p1 - p2 | ) the edge is not built, and the Error function will return
    	--    BRepAPI_LineThroughIdenticPoints.
    	-- Parameter values are expected to be given in increasing order:
    	--      C->FirstParameter() 
    	-- - If the parameter values are given in decreasing order the vertices are switched,
    	-- i.e. the "first vertex" is on the point of parameter p2 and the "second vertex" is
    	-- on the point of parameter p1. In such a case, to keep the original intent of the
    	-- construction, the edge will be oriented "reversed".
    	-- - On a periodic curve the parameter values p1 and p2 are adjusted by adding or
    	-- subtracting the period to obtain p1 in the parametric range of the curve, and p2]
    	-- such that [ p1 , where Period is the period of the curve.
    	-- - A parameter value may be infinite. The edge is open in the corresponding
    	-- direction. However the corresponding vertex must be a null shape. If this condition
    	-- is not satisfied the edge is not built, and the Error function will return
    	-- BRepAPI_PointWithInfiniteParameter.
    	-- - The distance between the vertex and the point evaluated on the curve with the
    	-- parameter, must be lower than the precision of the vertex. If this condition is not
    	-- satisfied the edge is not built, and the Error function will return
    	-- BRepAPI_DifferentsPointAndParameter.
    	--  Other edge constructions
    	-- - The parameter values can be omitted, they will be computed by projecting the
    	-- vertices on the curve. Note that projection is the only way to evaluate the
    	-- parameter values of the vertices on the curve: vertices must be given on the curve,
    	-- i.e. the distance from a vertex to the curve must be less than or equal to the
    	-- precision of the vertex. If this condition is not satisfied the edge is not built,
    	-- and the Error function will return BRepAPI_PointProjectionFailed.
    	-- -      3D points can be given in place of vertices. Vertices will be created from the
    	--    points (with the default topological precision Precision::Confusion()). 
    	-- Note:
    	-- -      Giving vertices is useful when creating a connected edge.
    	-- -      If the parameter values correspond to the extremities of a closed curve,
    	--    points must be identical, or at least coincident. If this condition is not
    	--    satisfied the edge is not built, and the Error function will return
    	--   BRepAPI_DifferentPointsOnClosedCurve.
    	-- -      The vertices or points can be omitted if the parameter values are given. The
    	--    points will be computed from the parameters on the curve.
    	-- The vertices or points and the parameter values can be omitted. The first and last
    	--   parameters of the curve will then be used.   
        ----------------------------------------
    --  Auxiliary methods
    ----------------------------------------

    Init(me : in out; C      : Curve from Geom)
	---Level: Public
    is static;
    
    Init(me : in out; C      : Curve from Geom;
		      p1, p2 : Real)
	---Level: Public
    is static;		      
	
    Init(me : in out; C      : Curve from Geom;
    	    	      P1, P2 : Pnt   from gp)
	---Level: Public
    is static;		      
	
    Init(me : in out; C      : Curve  from Geom;
    	              V1, V2 : Vertex from TopoDS)
	---Level: Public
    is static;
	
    Init(me : in out; C      : Curve from Geom;
    	    	      P1, P2 : Pnt   from gp;
		      p1, p2 : Real)
	---Level: Public
    is static;		      
	
    Init(me : in out; C      : Curve  from Geom;
    	              V1, V2 : Vertex from TopoDS;
		      p1, p2 : Real)
	---Level: Public
    is static;
	
    Init(me : in out; C      : Curve from Geom2d; S : Surface from Geom)
	---Level: Public
    is static;
    
    Init(me : in out; C      : Curve from Geom2d; S : Surface from Geom;
		      p1, p2 : Real)
	---Level: Public
    is static;		      
	
    Init(me : in out; C      : Curve from Geom2d; S : Surface from Geom;
    	    	      P1, P2 : Pnt   from gp)
	---Level: Public
    is static;		      
	
    Init(me : in out; C      : Curve  from Geom2d; S : Surface from Geom;
    	              V1, V2 : Vertex from TopoDS)
	---Level: Public
    is static;
	
    Init(me : in out; C      : Curve from Geom2d; S : Surface from Geom;
    	    	      P1, P2 : Pnt   from gp;
		      p1, p2 : Real)
	---Level: Public
    is static;		      
	
    Init(me : in out; C      : Curve  from Geom2d; S : Surface from Geom;
    	              V1, V2 : Vertex from TopoDS;
		      p1, p2 : Real)
	---Level: Public
    is static;
    	---Purpose: Defines or redefines the arguments for the construction of an edge.
    	-- This function is currently used after the empty constructor BRepAPI_MakeEdge().	

    ----------------------------------------
    --  Results
    ----------------------------------------

    IsDone(me) returns Boolean
	---Purpose: Returns true if the edge is built.
    is redefined;

    Error(me) returns EdgeError from BRepBuilderAPI
	---Purpose: Returns the construction status
        -- -   BRepBuilderAPI_EdgeDone if the edge is built, or
    	-- -   another value of the BRepBuilderAPI_EdgeError
    	--   enumeration indicating the reason of construction failure.
    is static;

    Edge(me) returns Edge from TopoDS
	---C++: return const &
	---C++: alias "Standard_EXPORT operator TopoDS_Edge() const;"
    	--- Purpose:
    	-- Returns the constructed edge.
    	-- Exceptions StdFail_NotDone if the edge is not built.
    raises
    	NotDone from StdFail
    is static;
    
    Vertex1(me) returns Vertex from TopoDS
	---Purpose: Returns the first vertex of the edge. May be Null.
	--          
	---C++: return const &
	---Level: Public
    is static;
    
    Vertex2(me) returns Vertex from TopoDS
		---C++: return const &
    	---Purpose: Returns the second vertex of the edge. May be Null.
	--          
	-- Warning
    	-- The returned vertex in each function corresponds respectively to
    	-- -   the lowest, or
    	-- -   the highest parameter on the curve along which the edge is built.
    	--  It does not correspond to the first or second vertex
    	-- given at the time of the construction, if the edge is oriented reversed.
    	-- Exceptions
    	-- StdFail_NotDone if the edge is not built.
    is static; 
    
fields

    myMakeEdge : MakeEdge  from BRepLib;

end MakeEdge;
