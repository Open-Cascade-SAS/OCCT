-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class CameraModelD3 from StepVisual 

inherits CameraModel from StepVisual 

uses

	Axis2Placement3d from StepGeom, 
	ViewVolume from StepVisual, 
	HAsciiString from TCollection
is

	Create returns mutable CameraModelD3;
	---Purpose: Returns a CameraModelD3


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aViewReferenceSystem : mutable Axis2Placement3d from StepGeom;
	      aPerspectiveOfVolume : mutable ViewVolume from StepVisual) is virtual;

	-- Specific Methods for Field Data Access --

	SetViewReferenceSystem(me : mutable; aViewReferenceSystem : mutable Axis2Placement3d);
	ViewReferenceSystem (me) returns mutable Axis2Placement3d;
	SetPerspectiveOfVolume(me : mutable; aPerspectiveOfVolume : mutable ViewVolume);
	PerspectiveOfVolume (me) returns mutable ViewVolume;

fields

	viewReferenceSystem : Axis2Placement3d from StepGeom;
	perspectiveOfVolume : ViewVolume from StepVisual;

end CameraModelD3;
