-- Created on: 1993-09-22
-- Created by: Didier PIFFAULT
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Vertex from BRepMesh 

  ---Purpose: 


uses    Boolean from Standard,
        Integer from Standard,
        Real from Standard,
        XY from gp,
        DegreeOfFreedom from BRepMesh


is        Create     returns Vertex from BRepMesh;

          Create         (UV      : in XY from gp;
                          Locat3d : in Integer from Standard;
                          Move    : in DegreeOfFreedom from BRepMesh)
            returns Vertex from BRepMesh;


          Create         (U, V    : Real from Standard;
                          Move    : in DegreeOfFreedom from BRepMesh)
            returns Vertex from BRepMesh;


          Initialize     (me      : in out;
                          UV      : in XY from gp; 
                          Locat3d : in Integer from Standard;
                          Move    : in DegreeOfFreedom from BRepMesh)
            is static;


          Coord          (me) 
            returns XY from gp
            ---C++: return const &
            ---C++: inline
            is static;


          Location3d    (me) 
            returns Integer from Standard
            ---C++: inline
            is static;


          Movability     (me)
            returns DegreeOfFreedom from BRepMesh
            ---C++: inline
            is static;

          SetMovability  (me   : in out;
                          Move : DegreeOfFreedom from BRepMesh)
            is static;


          HashCode       (me;
                          Upper : Integer from Standard)
            returns Integer from Standard
            ---C++: function call
            is static;


          IsEqual        (me; Other : Vertex from BRepMesh)
            returns Boolean from Standard
            ---C++: alias operator ==
            is static;


        fields  myUV         : XY from gp;
                myLocation   : Integer from Standard;
                myMovability : DegreeOfFreedom from BRepMesh;

end Vertex;
