-- File:        AutoDesignOrganizationAssignment.cdl
-- Created:     Fri Dec  1 11:11:14 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class AutoDesignOrganizationAssignment from StepAP214 

inherits OrganizationAssignment from StepBasic 

uses

	HArray1OfAutoDesignGeneralOrgItem from StepAP214, 
	AutoDesignGeneralOrgItem from StepAP214, 
	Organization from StepBasic, 
	OrganizationRole from StepBasic
is

	Create returns mutable AutoDesignOrganizationAssignment;
	---Purpose: Returns a AutoDesignOrganizationAssignment


	Init (me : mutable;
	      aAssignedOrganization : mutable Organization from StepBasic;
	      aRole : mutable OrganizationRole from StepBasic) is redefined;

	Init (me : mutable;
	      aAssignedOrganization : mutable Organization from StepBasic;
	      aRole : mutable OrganizationRole from StepBasic;
	      aItems : mutable HArray1OfAutoDesignGeneralOrgItem from StepAP214) is virtual;

	-- Specific Methods for Field Data Access --

	SetItems(me : mutable; aItems : mutable HArray1OfAutoDesignGeneralOrgItem);
	Items (me) returns mutable HArray1OfAutoDesignGeneralOrgItem;
	ItemsValue (me; num : Integer) returns AutoDesignGeneralOrgItem;
	NbItems (me) returns Integer;

fields

	items : HArray1OfAutoDesignGeneralOrgItem from StepAP214; -- a SelectType

end AutoDesignOrganizationAssignment;
