-- Created on: 1993-03-24
-- Created by: JCV
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class BezierCurve from Geom2d inherits BoundedCurve from Geom2d

        --- Purpose : Describes a rational or non-rational Bezier curve
    	-- - a non-rational Bezier curve is defined by a table
    	--   of poles (also called control points),
    	-- - a rational Bezier curve is defined by a table of
    	--   poles with varying weights.
    	-- These data are manipulated by two parallel arrays:
    	-- - the poles table, which is an array of gp_Pnt2d points, and
    	-- - the weights table, which is an array of reals.
    	-- The bounds of these arrays are 1 and "the number of poles" of the curve.
    	-- The poles of the curve are "control points" used to deform the curve.
    	-- The first pole is the start point of the curve, and the
    	-- last pole is the end point of the curve. The segment
    	-- which joins the first pole to the second pole is the
    	-- tangent to the curve at its start point, and the
    	-- segment which joins the last pole to the
    	-- second-from-last pole is the tangent to the curve
    	-- at its end point.
    	-- It is more difficult to give a geometric signification
    	-- to the weights but they are useful for providing
    	-- exact representations of the arcs of a circle or
    	-- ellipse. Moreover, if the weights of all the poles are
    	-- equal, the curve is polynomial; it is therefore a
    	-- non-rational curve. The non-rational curve is a
    	-- special and frequently used case. The weights are
    	-- defined and used only in case of a rational curve.
    	-- The degree of a Bezier curve is equal to the
    	-- number of poles, minus 1. It must be greater than or
    	-- equal to 1. However, the degree of a
    	-- Geom2d_BezierCurve curve is limited to a value
    	-- (25) which is defined and controlled by the system.
    	-- This value is returned by the function MaxDegree.
    	-- The parameter range for a Bezier curve is [ 0, 1 ].
    	-- If the first and last control points of the Bezier
    	-- curve are the same point then the curve is closed.
    	-- For example, to create a closed Bezier curve with
    	-- four control points, you have to give a set of control
    	-- points P1, P2, P3 and P1.
    	-- The continuity of a Bezier curve is infinite.
    	-- It is not possible to build a Bezier curve with
    	-- negative weights. We consider that a weight value
    	-- is zero if it is less than or equal to
    	-- gp::Resolution(). We also consider that
    	-- two weight values W1 and W2 are equal if:
    	-- |W2 - W1| <= gp::Resolution().
    	--  Warning
    	-- - When considering the continuity of a closed
    	--   Bezier curve at the junction point, remember that
    	--   a curve of this type is never periodic. This means
    	--   that the derivatives for the parameter u = 0
    	--   have no reason to be the same as the
    	--   derivatives for the parameter u = 1 even if the curve is closed.
    	-- - The length of a Bezier curve can be null.


uses  Array1OfReal        from TColStd,
      HArray1OfReal       from TColStd,
      Array1OfPnt2d       from TColgp,
      Ax2d                from gp,
      Pnt2d               from gp, 
      HArray1OfPnt2d      from TColgp, 
      Vec2d               from gp, 
      Trsf2d              from gp,
      Geometry            from Geom2d,
      Shape               from GeomAbs


raises ConstructionError from Standard,
       DimensionError    from Standard,
       RangeError        from Standard,
       OutOfRange        from Standard


is 




  Create (CurvePoles : Array1OfPnt2d from TColgp) returns mutable BezierCurve
        --- Purpose :
        --  Creates a non rational Bezier curve with a set of poles :
        --  CurvePoles.  The weights are defaulted to all being 1. 
    	--    Raises ConstructionError if the number of poles is greater than MaxDegree + 1
        --  or lower than 2.
     raises ConstructionError;
   

  Create (CurvePoles  : Array1OfPnt2d from TColgp;
    	  PoleWeights : Array1OfReal from TColStd) 
     returns mutable BezierCurve
        --- Purpose :
        --  Creates a rational Bezier curve with the set of poles
        --  CurvePoles and the set of weights  PoleWeights .
        --  If all the weights are identical the curve is considered 
        --  as non rational.  Raises ConstructionError if 
        --  the number of poles is greater than  MaxDegree + 1 or lower
        --  than 2 or CurvePoles and CurveWeights have not the same length
        --  or one weight value is lower or equal to Resolution from
        --  package gp.
     raises ConstructionError;
     

  Increase (me : mutable; Degree : Integer)
        --- Purpose :
        --  Increases the degree of a bezier curve. Degree is the new 
        --  degree of <me>.
    	--    raises ConstructionError if Degree is greater than MaxDegree or lower than 2 
        --  or lower than the initial degree of <me>.

     raises ConstructionError;
      


  InsertPoleAfter (me : mutable; Index : Integer; P : Pnt2d;
     	    	   Weight : Real = 1.0)
        --- Purpose :
        --  Inserts a pole with its weight in the set of poles after the
        --  pole of range Index. If the curve was non rational it can
        --  become rational if all the weights are not identical.
     raises OutOfRange,
        --- Purpose : Raised if Index is not in the range [0, NbPoles]
            ConstructionError;
        --- Purpose : 
        --  Raised if the resulting number of poles is greater than 
        --  MaxDegree + 1.


  InsertPoleBefore (me : mutable; Index : Integer; P : Pnt2d;
    	    	    Weight : Real = 1.0)
        --- Purpose :
        --  Inserts a pole with its weight in the set of poles after 
        --  the pole of range Index. If the curve was non rational it
        --  can become rational if all the weights are not identical.
     raises OutOfRange,
        --- Purpose : Raised if Index is not in the range [1, NbPoles+1]
            ConstructionError;
        --- Purpose : 
        --  Raised if the resulting number of poles is greater than 
        --  MaxDegree + 1.


  RemovePole (me : mutable; Index : Integer)
        --- Purpose : Removes the pole of range Index.
        --  If the curve was rational it can become non rational.
     raises OutOfRange,
        --- Purpose : Raised if Index is not in the range [1, NbPoles]
            ConstructionError;
         -- Purpose : Raised if Degree is lower than 2.


  Reverse (me : mutable);
        --- Purpose :
        --  Reverses the direction of parametrization of <me>
        --  Value (NewU) =  Value (1 - OldU)


  ReversedParameter(me; U : Real) returns Real;
	---Purpose: Returns the  parameter on the  reversed  curve for
	--          the point of parameter U on <me>.
	--          
	--          returns 1-U


  Segment (me : mutable; U1, U2 : Real);
        --- Purpose :
        --  Segments the curve between U1 and U2 which can be out
        --  of the bounds of the curve. The curve is oriented from U1
        --  to U2.
        --  The control points are modified, the first and the last point
        --  are not the same but the parametrization range is [0, 1] 
        --  else it could not be a Bezier curve.
        -- Warnings :
        --  Even if <me> is not closed it can become closed after the 
        --  segmentation for example if U1 or U2 are out of the bounds 
        --  of the curve <me> or if the curve makes loop.
        --  After the segmentation the length of a curve can be null.


  SetPole (me : mutable; Index : Integer; P : Pnt2d)
        --- Purpose :
        --  Substitutes the pole of range index with P.
        --  If the curve <me> is rational the weight of range Index 
        --  is not modified.
     raises OutOfRange;
        --- Purpose : raiseD if Index is not in the range [1, NbPoles]


  SetPole (me : mutable; Index : Integer; P : Pnt2d; Weight : Real)
        --- Purpose :
        --  Substitutes the pole and the weights of range Index.
        --  If the curve <me> is not rational it can become rational 
        --  if all the weights are not identical.
        --  If the curve was rational it can become non rational if
        --  all the weights are identical.
     raises OutOfRange,
        --- Purpose : Raised if Index is not in the range [1, NbPoles]
            ConstructionError;
        --- Purpose : Raised if Weight <= Resolution from package gp


  SetWeight (me : mutable; Index : Integer; Weight : Real)
        --- Purpose :
        --  Changes the weight of the pole of range Index.
        --  If the curve <me> is not rational it can become rational 
        --  if all the weights are not identical.
        --  If the curve was rational it can become non rational if
        --  all the weights are identical.
     raises OutOfRange,
        --- Purpose : Raised if Index is not in the range [1, NbPoles]
            ConstructionError;
        --- Purpose : Raised if Weight <= Resolution from package gp



  IsClosed (me)   returns Boolean;
        --- Purpose :
        --  Returns True if the distance between the first point 
        --  and the last point of the curve is lower or equal to
        --  the Resolution from package gp.


  IsCN (me; N : Integer)   returns Boolean;
        --- Purpose : Continuity of the curve, returns True. 


  IsPeriodic (me)   returns Boolean;
        --- Purpose : 
        --  Returns False. A BezierCurve cannot be periodic in this
        --  package


  IsRational (me)   returns Boolean;
        --- Purpose :
        --  Returns false if all the weights are identical. The tolerance
        --  criterion is Resolution from package gp.


  Continuity (me)   returns Shape from GeomAbs;
        --- Purpose :  Returns GeomAbs_CN, which is the continuity of any Bezier curve.


  Degree (me)   returns Integer;
        --- Purpose : 
        --  Returns the polynomial degree of the curve. It is the number 
        --  of poles less one.  In this package the Degree of a Bezier
        --  curve cannot be greater than "MaxDegree".






  D0 (me; U : Real; P : out Pnt2d);

  D1 (me; U : Real; P : out Pnt2d; V1 : out Vec2d);

  D2 (me; U : Real; P : out Pnt2d; V1, V2 : out Vec2d);

  D3 (me; U : Real; P : out Pnt2d; V1, V2, V3 : out Vec2d);

  DN (me; U : Real; N : Integer)  returns Vec2d
        --- Purpose :  For this Bezier curve, computes
    	-- - the point P of parameter U, or
    	-- - the point P and one or more of the following values:
    	--   - V1, the first derivative vector,
    	--   - V2, the second derivative vector,
    	--   - V3, the third derivative vector.
    	-- Note: the parameter U can be outside the bounds of the curve.
    	--     Raises RangeError if N < 1.
     raises RangeError;

  EndPoint (me) returns Pnt2d;
        --- Purpose :    Returns the end point or start point of this Bezier curve.
      

  FirstParameter (me) returns Real;
        --- Purpose : Returns the value of the first  parameter of this
    	-- Bezier curve. This is  0.0, which gives the start point of this Bezier curve.


  LastParameter (me) returns Real;
        --- Purpose : Returns the value of the last  parameter of this
    	-- Bezier curve. This is  1.0, which gives the end point of this Bezier curve.


  NbPoles (me)  returns Integer;

    	---Purpose: Returns the number of poles for this Bezier curve.
    
  Pole (me; Index : Integer) returns Pnt2d
        --- Purpose : Returns the pole of range Index.
     raises OutOfRange;
        --- Purpose : Raised if Index is not in the range [1, NbPoles]


  Poles (me; P : out Array1OfPnt2d from TColgp)
        --- Purpose : Returns all the poles of the curve.
     raises DimensionError;
        --- Purpose : 
        --  Raised if the length of P is not equal to the number of poles.


  StartPoint (me)  returns Pnt2d;
        --- Purpose :
        --  Returns Value (U=1), it is the first control point
        --  of the curve.


  Weight (me; Index : Integer)   returns Real  
        --- Purpose : Returns the weight of range Index.
     raises OutOfRange;
        --- Purpose : Raised if Index is not in the range [1, NbPoles]


  Weights (me; W : out Array1OfReal from TColStd)
        --- Purpose : Returns all the weights of the curve.
     raises DimensionError;
        --- Purpose : 
        --  Raised if the length of W is not equal to the number of poles.
        



  Transform (me : mutable; T : Trsf2d);

    	---Purpose: Applies the transformation T to this Bezier curve.
	     

  MaxDegree (myclass)   returns Integer;
        --- Purpose:
        --  Returns the value of the maximum polynomial degree of a 
        --  BezierCurve. This value is 25.



  Resolution(me          : mutable; 
    	     ToleranceUV : Real;
             UTolerance  : out Real);
	---Purpose:  Computes for this Bezier curve the parametric
    	-- tolerance UTolerance for a given tolerance
    	-- Tolerance3D (relative to dimensions in the plane).
    	-- If f(t) is the equation of this Bezier curve,
    	-- UTolerance ensures that
	--           | t1 - t0| < Utolerance ===> 
	--           |f(t1) - f(t0)| < ToleranceUV

  Copy (me)  returns mutable like me;
    	---Purpose: Creates a new object which is a copy of this Bezier curve.     

  Init (me : mutable; Poles   :  HArray1OfPnt2d  from TColgp;
    	              Weights : HArray1OfReal    from TColStd) 
  
        ---Purpose : Set  poles  to  Poles,  weights to  Weights  (not
        --         copied). If Weights is   null  the  curve is    non
        --         rational. Create the arrays of coefficients.  Poles
        --         and    Weights  are   assumed   to  have the  first
        --         coefficient 1.
        --         
        --         Update rational and closed.
        --         
  raises ConstructionError -- if nbpoles < 2 or nbboles > MaDegree + 1

  is static private;
  
  CoefficientsOK(me; U : Real) returns Boolean
  
        ---Purpose : returns true if the coefficients have been
        --           computed with the right value of cacheparameter
        --           for the given U value.
        -- 
        is static private;
  
  UpdateCoefficients(me : mutable; U : Real from Standard = 0.0)
    	---Purpose: Recompute the coeficients.
  is static private;



fields

   rational : Boolean;
   closed   : Boolean;
   poles    : HArray1OfPnt2d from TColgp;
   weights  : HArray1OfReal from TColStd;

   coeffs   : HArray1OfPnt2d from TColgp;
   wcoeffs  : HArray1OfReal from TColStd;

   validcache      : Integer;
   -- = 1 the cache is valid 
   -- = 0 the cache is invalid
   parametercache    : Real;
   -- Parameter at which the Taylor expension is stored in 
   -- the cache, often 0., sometimes 1..
   spanlenghtcache   : Real;
   -- always 1. for the moment.

   -- usefull to evaluate the parametric resolution
   maxderivinv   : Real from Standard;
   maxderivinvok : Boolean from Standard;

end;
