-- File:	IGESGeom_ToolOffsetSurface.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolOffsetSurface  from IGESGeom

    ---Purpose : Tool to work on a OffsetSurface. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses OffsetSurface from IGESGeom,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolOffsetSurface;
    ---Purpose : Returns a ToolOffsetSurface, ready to work


    ReadOwnParams (me; ent : mutable OffsetSurface;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : OffsetSurface;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : OffsetSurface;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a OffsetSurface <ent>, from
    --           its specific (own) parameters

    DirChecker (me; ent : OffsetSurface) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : OffsetSurface;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : OffsetSurface; entto : mutable OffsetSurface;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : OffsetSurface;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolOffsetSurface;
