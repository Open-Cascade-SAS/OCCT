-- Created on: 1994-03-25
-- Created by: Jean Marc LACHAUME
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class IsoBuilder from DBRep

	---Purpose: Creation of isoparametric curves.

inherits Hatcher from Geom2dHatch

uses

    Face from TopoDS ,
    Face from DBRep ,
    Array1OfReal    from TColStd ,
    Array1OfInteger from TColStd
    

is

    Create (TopologicalFace : Face    from TopoDS ;
    	    Infinite        : Real    from Standard ;
    	    NbIsos          : Integer from Standard)

    	---Purpose: Creates the builder.

    	returns IsoBuilder from DBRep ;


    NbDomains (me)

    	---Purpose: Returns the total number of domains.

    	---C++: inline

    	returns Integer from Standard
    	is static ;


    LoadIsos (me; Face : mutable Face from DBRep)

    	---Purpose: Loading of the isoparametric curves in the
    	--          Data Structure of a drawable face.

    	is static ;


fields

    myInfinite : Real            from Standard ;
    myUMin     : Real            from Standard ;
    myUMax     : Real            from Standard ;
    myVMin     : Real            from Standard ;
    myVMax     : Real            from Standard ;
    myUPrm     : Array1OfReal    from TColStd ;
    myUInd     : Array1OfInteger from TColStd ;    
    myVPrm     : Array1OfReal    from TColStd ;
    myVInd     : Array1OfInteger from TColStd ;    
    myNbDom    : Integer         from Standard ;
    
end IsoBuilder;
