-- Created on: 1994-12-16
-- Created by: Frederic MAUPAS
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class TranslatePolyLoop from StepToTopoDS
    inherits Root from StepToTopoDS
    
    ---Purpose:
    --         

uses

    PolyLoop               from StepShape,
    TranslatePolyLoopError from StepToTopoDS,
    Tool                   from StepToTopoDS,
    Surface                from Geom,
    Face                   from TopoDS,
    Shape                  from TopoDS
    
raises NotDone from StdFail

is

    Create returns TranslatePolyLoop;
    
    Create (PL : PolyLoop    from StepShape;
    	    T  : in out Tool from StepToTopoDS;
    	    S  : Surface     from Geom;
    	    F  : Face        from TopoDS)
    	returns TranslatePolyLoop;
	    
    Init (me : in out;
    	  PL : PolyLoop from StepShape;
    	  T  : in out Tool from StepToTopoDS;
    	  S  : Surface     from Geom;
    	  F  : Face        from TopoDS);

    Value (me) returns Shape from TopoDS
    	raises NotDone
	is static;
	---C++: return const &

    Error (me) returns TranslatePolyLoopError from StepToTopoDS;
    
fields

    myError  : TranslatePolyLoopError from StepToTopoDS;
    
    myResult : Shape                  from TopoDS;
    
end TranslatePolyLoop;
