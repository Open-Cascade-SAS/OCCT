-- Created by: Peter KURNEV
-- Copyright (c) 2010-2014 OPEN CASCADE SAS
-- Copyright (c) 2007-2010 CEA/DEN, EDF R&D, OPEN CASCADE
-- Copyright (c) 2003-2007 OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN, CEDRAT,
--                         EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class BuilderSolid from BOPAlgo 
    inherits BuilderArea from BOPAlgo 
 
---Purpose: The algorithm to build solids from set of faces  

uses 
    BaseAllocator from BOPCol,
    Solid from TopoDS 
    
--raises

is 
    Create  
    returns BuilderSolid from BOPAlgo; 
    ---C++: alias "Standard_EXPORT virtual ~BOPAlgo_BuilderSolid();" 
     
      
    Create (theAllocator: BaseAllocator from BOPCol) 
    returns BuilderSolid from BOPAlgo; 
      
    SetSolid(me:out; 
            theSolid:Solid from TopoDS); 
    ---Purpose: Sets the source solid <theSolid>   
     
    Solid(me) 
    	 returns Solid from TopoDS; 
    ---C++:  return const &	 
    ---Purpose: Returns the source solid 
     
    Perform(me:out)  
    ---Purpose:  Performs the algorithm 
    is redefined;  
 
    PerformShapesToAvoid(me:out) 
    ---Purpose:  Collect the faces that 
    --           a) are internal        	 
    --           b) are the same and have different orientation         
    is redefined protected; 
	 
    PerformLoops(me:out) 
    ---Purpose: Build draft shells 
    --          a)myLoops - draft shells that consist of  
    --                       boundary faces 
    --          b)myLoopsInternal - draft shells that contains 
    --                               inner faces 
    is redefined protected;  
	 
    PerformAreas(me:out)   
    ---Purpose: Build draft solids that contains boundary faces   
    is redefined protected;  

    PerformInternalShapes(me:out)   
    ---Purpose: Build finalized solids with internal shells   
    is redefined protected;   

fields 
    mySolid:Solid from TopoDS is protected;       
  
end BuilderSolid; 
