-- Created on: 1993-02-02
-- Created by: Christian CAILLET
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class GeneralModule  from StepData
         inherits GeneralModule from Interface

    ---Purpose : Specific features for General Services adapted to STEP

uses Transient ,
     EntityIterator , CopyTool, Check, ShareTool

is

    	--  Reconduction because limitation cdl  --

    FillSharedCase (me; casenum : Integer; ent : Transient;
    	iter : in out EntityIterator)  is deferred;
    ---Purpose : Specific filling of the list of Entities shared by an Entity
    --           <ent>. Can use the internal utility method Share, below

    CheckCase (me; casenum : Integer; ent : Transient; shares : ShareTool;
    	       ach : in out Check)  is deferred;
    ---Purpose : Specific Checking of an Entity <ent>

    CopyCase (me; casenum : Integer;
    	      entfrom : Transient; entto : Transient;
    	      TC : in out CopyTool)  is deferred;
    ---Purpose : Specific Copy ("Deep") from <entfrom> to <entto> (same type)
    --           by using a TransferControl which provides its working Map.
    --           Use method Transferred from TransferControl to work

--    ImpliedCase (me; casenum : Integer;
--    	         entfrom : Transient; entto : Transient;
--    	         TC : CopyTool);
    ---Purpose : Specific Copying of Implied References
    --           A Default is provided which does nothing (must current case !)
    --           Already copied references (by CopyFrom) must remain unchanged
    --           Use method Search from TransferControl to work

end GeneralModule;
