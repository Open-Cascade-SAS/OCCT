-- File:	RWStepRepr_RWAssemblyComponentUsage.cdl
-- Created:	Mon Jul  3 19:47:50 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class RWAssemblyComponentUsage from RWStepRepr

    ---Purpose: Read & Write tool for AssemblyComponentUsage

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    AssemblyComponentUsage from StepRepr

is
    Create returns RWAssemblyComponentUsage from RWStepRepr;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : AssemblyComponentUsage from StepRepr);
	---Purpose: Reads AssemblyComponentUsage

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: AssemblyComponentUsage from StepRepr);
	---Purpose: Writes AssemblyComponentUsage

    Share (me; ent : AssemblyComponentUsage from StepRepr;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWAssemblyComponentUsage;
