-- Created on: 1993-11-09
-- Created by: Modelistation
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class CompBezierCurves2dToBSplineCurve2d from Convert 

	---Purpose: Converts a list  of connecting Bezier Curves 2d to  a
	--          BSplineCurve 2d.
	--          if possible, the continuity of the BSpline will be 
	--          increased to more than C0.


uses
    SequenceOfReal            from TColStd,
    SequenceOfInteger         from TColStd,
    Array1OfReal              from TColStd,
    Array1OfInteger           from TColStd,
    Array1OfPnt2d             from TColgp,
    SequenceOfPnt2d           from TColgp,
    SequenceOfArray1OfPoles2d from Convert


raises
    ConstructionError from Standard

    -------------------------------------------------------------------------
    --- Don't forget to use the method Perform before accessing the Result.
    -------------------------------------------------------------------------

is
    Create( AngularTolerance : Real = 1.0e-4 )
    returns CompBezierCurves2dToBSplineCurve2d from Convert;
    	---Purpose: Constructs a framework for converting a sequence of
    	-- adjacent non-rational Bezier curves into a BSpline curve.
    	-- Knots will be created on the computed BSpline curve at
    	-- each junction point of two consecutive Bezier curves. The
    	-- degree of continuity of the BSpline curve will be increased at
    	-- the junction point of two consecutive Bezier curves if their
    	-- tangent vectors at this point are parallel. AngularTolerance
    	-- (given in radians, and defaulted to 1.0 e-4) will be used
    	-- to check the parallelism of the two tangent vectors.
    	-- Use the following functions:
    	-- -   AddCurve to define in sequence the adjacent Bezier
    	--  curves to be converted,
    	-- -   Perform to compute the data needed to build the BSpline curve,
    	-- -   and the available consultation functions to access the
    	--  computed data. This data may be used to construct the BSpline curve.
  
    AddCurve( me    : in out;
              Poles : Array1OfPnt2d from TColgp)
    is static;
    	--- Purpose: Adds the Bezier curve defined by the table of poles Poles, to
    	--  the sequence (still contained in this framework) of adjacent
    	-- Bezier curves to be converted into a BSpline curve.
    	-- Only polynomial (i.e. non-rational) Bezier curves are
    	-- converted using this framework.
    	-- If this is not the first call to the function (i.e. if this framework
    	-- still contains data in its sequence of Bezier curves), the
    	-- degree of continuity of the BSpline curve will be increased at
    	-- the time of computation at the first point of the added Bezier
    	-- curve (i.e. the first point of the Poles table). This will be the
    	-- case if the tangent vector of the curve at this point is
    	-- parallel to the tangent vector at the end point of the
    	-- preceding Bezier curve in the sequence of Bezier curves still
    	-- contained in this framework. An angular tolerance given at
    	-- the time of construction of this framework, will be used to
    	-- check the parallelism of the two tangent vectors. This
    	-- checking procedure, and all the relative computations will be
    	-- performed by the function Perform.
    	-- When the sequence of adjacent Bezier curves is complete,
    	-- use the following functions:
    	-- -   Perform to compute the data needed to build the BSpline curve,
    	-- -   and the available consultation functions to access the
    	--  computed data. This data may be used to construct the BSpline curve.
    	--  Warning
    	-- The sequence of Bezier curves treated by this framework is
    	-- automatically initialized with the first Bezier curve when the
    	-- function is first called. During subsequent use of this function,
    	-- ensure that the first point of the added Bezier curve (i.e. the
    	-- first point of the Poles table) is coincident with the last point
    	-- of the sequence (i.e. the last point of the preceding Bezier
    	-- curve in the sequence) of Bezier curves still contained in
    	-- this framework. An error may occur at the time of
    	-- computation if this condition is not satisfied. Particular care
    	-- must be taken with respect to the above, as this condition is
    	-- not checked either when defining the sequence of Bezier
    	-- curves or at the time of computation.


    Perform(me: in out)
    	---Purpose: Computes all the data needed to build a BSpline curve
    	-- equivalent to the sequence of adjacent Bezier curves still
    	-- contained in this framework.
    	-- A knot is inserted on the computed BSpline curve at the
    	-- junction point of two consecutive Bezier curves. The
    	-- degree of continuity of the BSpline curve will be increased
    	-- at the junction point of two consecutive Bezier curves if
    	-- their tangent vectors at this point are parallel. An angular
    	-- tolerance given at the time of construction of this
    	-- framework is used to check the parallelism of the two
    	-- tangent vectors.
    	-- Use the available consultation functions to access the
    	-- computed data. This data may then be used to construct
    	-- the BSpline curve.
    	-- Warning
    	-- Ensure that the curves in the sequence of Bezier curves
    	-- contained in this framework are adjacent. An error may
    	-- occur at the time of computation if this condition is not
    	-- satisfied. Particular care must be taken with respect to the
    	-- above as this condition is not checked, either when
    	-- defining the Bezier curve sequence or at the time of computation.
    is static;

    
    Degree(me) returns Integer from Standard
    is static;
    	---Purpose: Returns the degree of the BSpline curve whose data is
    	-- computed in this framework.
    	-- Warning
    	-- Take particular care not to use this function before the
    	-- computation is performed (Perform function), as this
    	-- condition is not checked and an error may therefore occur.
    
    NbPoles(me) returns Integer from Standard
    is static;
   	---Purpose: Returns the number of poles of the BSpline curve whose
    	-- data is computed in this framework.
    	-- Warning
    	-- Take particular care not to use this function before the
    	-- computation is performed (Perform function), as this
    	-- condition is not checked and an error may therefore occur.
 
    Poles(me; Poles : in out Array1OfPnt2d from TColgp)
    is static;
 	--- Purpose: Loads the Poles table with the poles of the BSpline curve
    	-- whose data is computed in this framework.
    	-- Warning
    	-- -   Do not use this function before the computation is
    	--  performed (Perform function).
    	-- -   The length of the Poles array must be equal to the
    	--  number of poles of the BSpline curve whose data is
    	--  computed in this framework.
    	-- Particular care must be taken with respect to the above, as
    	-- these conditions are not checked, and an error may occur.
 
    NbKnots(me) returns Integer from Standard
    is static;
 	--- Purpose: Returns the number of knots of the BSpline curve whose
    	-- data is computed in this framework.
    	-- Warning
    	-- Take particular care not to use this function before the
    	-- computation is performed (Perform function), as this
    	-- condition is not checked and an error may therefore occur.
 
    KnotsAndMults(me;
                  Knots : in out Array1OfReal    from TColStd;
		  Mults : in out Array1OfInteger from TColStd)
    is static; 
    	--- Purpose: Loads the Knots table with the knots
    	-- and the Mults table with the corresponding multiplicities
    	-- of the BSpline curve whose data is computed in this framework.
    	-- Warning
    	-- -   Do not use this function before the computation is
    	--  performed (Perform function).
    	-- -   The length of the Knots and Mults arrays must be equal
    	--  to the number of knots in the BSpline curve whose data is
    	--  computed in this framework.
    	-- Particular care must be taken with respect to the above as
    	-- these conditions are not checked, and an error may occur.
 
    
fields
    mySequence          : SequenceOfArray1OfPoles2d from Convert;
    CurvePoles          : SequenceOfPnt2d           from TColgp;
    CurveKnots          : SequenceOfReal            from TColStd;
    KnotsMultiplicities : SequenceOfInteger         from TColStd;
    myDegree            : Integer                   from Standard;
    myAngular           : Real                      from Standard;
    myDone              : Boolean                   from Standard;

end CompBezierCurves2dToBSplineCurve2d;
