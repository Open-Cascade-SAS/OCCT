-- Created on: 1995-12-08
-- Created by: Laurent BOURESCHE
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class CornerState from GeomFill 

	---Purpose: Class  (should    be  a  structure)   storing  the
	--          informations         about     continuity, normals
	--          parallelism,  coons conditions and bounds tangents
	--          angle on the corner of contour to be filled.

is

    Create returns CornerState from GeomFill;
    Gap(me) returns Real from Standard;
    Gap(me : in out; G : Real from Standard);
    TgtAng(me) returns Real from Standard;
    TgtAng(me : in out; Ang : Real from Standard);
    HasConstraint(me) returns Boolean from Standard;
    Constraint(me : in out);
    NorAng(me) returns Real from Standard;
    NorAng(me : in out; Ang : Real from Standard);
    IsToKill(me; Scal : out Real from Standard) 
    returns Boolean from Standard;
    DoKill(me : in out; Scal : Real from Standard);
    
fields

    gap           : Real from Standard;
    tgtang        : Real from Standard;
    isconstrained : Boolean from Standard;
    norang        : Real from Standard;
    scal          : Real from Standard;
    coonscnd      : Boolean from Standard;

end CornerState;
