-- Created on: 1997-05-06
-- Created by: Yves FRICAUD
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



private class IteratorOnShapesSet from TNaming 

	---Purpose: 

uses
    ShapesSet               from TNaming,
    Shape                   from TopoDS,
    MapIteratorOfMapOfShape from TopTools
    
raises
    NoMoreObject from Standard,
    NoSuchObject from Standard

is
    Create returns IteratorOnShapesSet;
         ---C++: inline

    Create (S : ShapesSet from TNaming) returns IteratorOnShapesSet;    	
    	 ---C++: inline
    
    Init (me : in out; S : ShapesSet from TNaming);
	---Purpose: Initialize the iteration
    	---C++: inline
    
    More (me) returns Boolean;
	---Purpose: Returns True if there is a current Item in
	--          the iteration.
    	---C++: inline
    
    Next (me : in out)
    	---Purpose: Move to the next Item 
    	---C++: inline
    raises
	NoMoreObject from Standard;
    
    Value(me) returns Shape from TopoDS
    	---C++: return const&
    raises
	NoSuchObject from Standard;


fields
    myIt    : MapIteratorOfMapOfShape from TopTools;

end IteratorOnShapesSet;
