-- File:        Block.cdl
-- Created:     Mon Dec  4 12:02:23 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWBlock from RWStepShape

	---Purpose : Read & Write Module for Block

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     Block from StepShape,
     EntityIterator from Interface

is

	Create returns RWBlock;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable Block from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : Block from StepShape);

	Share(me; ent : Block from StepShape; iter : in out EntityIterator);

end RWBlock;
