-- Created on: 1993-05-14
-- Created by: Laurent PAINNOT
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

generic class ComputeCLine from Approx 
    	    	    (MultiLine as any;
    	    	     LineTool  as any) --as TheLineTool from AppCont(MultiLine)


uses ParametrizationType       from Approx,
     SequenceOfReal            from TColStd,
     HArray1OfReal             from TColStd,
     SequenceOfMultiCurve      from AppParCurves,
     MultiCurve                from AppParCurves,
     Constraint                from AppParCurves,
     Vector                    from math
     
     

private class MyLeastSquare instantiates LeastSquare from AppCont
    	    	    	    	       (MultiLine,
			    	    	LineTool);
							  
is


    Create(Line:            MultiLine; 
    	   degreemin:       Integer    = 3;
           degreemax:       Integer    = 8;
    	   Tolerance3d:     Real       = 1.0e-5; 
    	   Tolerance2d:     Real       = 1.0e-5;
	   cutting:         Boolean    = Standard_False;
    	   FirstC:          Constraint = AppParCurves_TangencyPoint;
    	   LastC:           Constraint = AppParCurves_TangencyPoint)
	   
	---Purpose: The MultiLine <Line> will be approximated until tolerances
	--          will be reached.
	--          The approximation will be done from degreemin to degreemax
	--          with a cutting if the corresponding boolean is True.

    returns ComputeCLine;




    Create(degreemin:    Integer    = 3;
    	   degreemax:    Integer    = 8;
    	   Tolerance3d:  Real       = 1.0e-05; 
    	   Tolerance2d:  Real       = 1.0e-05; 
	   cutting:      Boolean    = Standard_False;
    	   FirstC:       Constraint = AppParCurves_TangencyPoint;
    	   LastC:        Constraint = AppParCurves_TangencyPoint)
	   
	---Purpose: Initializes the fields of the algorithm.

    returns ComputeCLine;


    Perform(me: in out; Line: MultiLine)
	---Purpose: runs the algorithm after having initialized the fields.
    
    is static;


    Compute(me: in out; Line: MultiLine; Ufirst, Ulast: Real;
    	    TheTol3d, TheTol2d: in out Real)
	---Purpose: is internally used by the algorithms.

    returns Boolean
    is static private;
    
    
    SetDegrees(me: in out; degreemin, degreemax: Integer)
    	---Purpose: changes the degrees of the approximation.
    
    is static;
    
    
    SetTolerances(me: in out; Tolerance3d, Tolerance2d: Real)
    	---Purpose: Changes the tolerances of the approximation.
    
    is static;
    

    SetConstraints(me: in out; FirstC, LastC: Constraint)
    	---Purpose: Changes the constraints of the approximation.
    
    is static;
    
    
    IsAllApproximated(me) 
    	---Purpose: returns False if at a moment of the approximation,
    	--          the status NoApproximation has been sent by the user
    	--          when more points were needed.
    
    returns Boolean
    is static;
    
    IsToleranceReached(me)
    	---Purpose: returns False if the status NoPointsAdded has been sent.
    
    returns Boolean
    is static;
    

    Error(me; Index: Integer; tol3d: in out Real; tol2d: in out Real)
    	---Purpose: returns the tolerances 2d and 3d of the <Index> MultiCurve.

    is static;
    

    NbMultiCurves(me)
    	---Purpose: Returns the number of MultiCurve doing the approximation
    	--          of the MultiLine.
    returns Integer
    is static;


    Value(me; Index: Integer = 1)
    	---Purpose: returns the approximation MultiCurve of range <Index>.

    returns MultiCurve from AppParCurves;

	    
    Parameters(me; Index: Integer; firstp, lastp: in out Real)
    	---purpose: returns the first and last parameters of the 
    	--          <Index> MultiCurve.
    is static;
	    

fields


myMultiCurves: SequenceOfMultiCurve from AppParCurves;    
myfirstparam:  SequenceOfReal       from TColStd;
mylastparam:   SequenceOfReal       from TColStd;
TheMultiCurve: MultiCurve from AppParCurves;
alldone:       Boolean;
tolreached:    Boolean;
Tolers3d:      SequenceOfReal from TColStd;
Tolers2d:      SequenceOfReal from TColStd;
mydegremin:    Integer;
mydegremax:    Integer;
mytol3d:       Real;
mytol2d:       Real;
currenttol3d:  Real;
currenttol2d:  Real;
mycut:         Boolean;
myfirstC:      Constraint;
mylastC:      Constraint;


end ComputeCLine;
