-- Created on: 1994-11-16
-- Created by: Marie Jose MARTZ
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class GeomPoint from GeomToIGES inherits GeomEntity from GeomToIGES

    ---Purpose: This class implements the transfer of the Point Entity from Geom
    --          to IGES . These are :
    --          . Point
    --              * CartesianPoint 

  
uses

    Point          from Geom,
    CartesianPoint from Geom,
    Point          from IGESGeom,
    GeomEntity     from GeomToIGES
     
is 
    
    Create returns GeomPoint from GeomToIGES;


    Create(GE : GeomEntity from GeomToIGES)  
    	 returns GeomPoint from GeomToIGES;
    ---Purpose : Creates a tool GeomPoint ready to run and sets its
    --         fields as GE's.

    TransferPoint            (me    : in out;
                              start : Point from Geom)
    	 returns mutable Point from IGESGeom;
    ---Purpose :  Transfert  a  Point from Geom to IGES. If this
    --            Entity could not be converted, this member returns a NullEntity.

    TransferPoint            (me    : in out;
                              start : CartesianPoint from Geom)
    	 returns mutable Point from IGESGeom;
    ---Purpose :  Transfert  a  CartesianPoint from Geom to IGES. If this
    --            Entity could not be converted, this member returns a NullEntity.


end GeomPoint;


