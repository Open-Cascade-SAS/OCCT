-- Created on: 1993-07-06
-- Created by: Jean Louis FRENKEL
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Modified:    stt: 25-02-98: S3558 ajout ViewStdAdapter
--              stt: 08-04-98: suppr ViewStdAdapter


package V2d
---Purpose: this package furnishes the services needed to build a
--          2d mono-view visualizer on a windowing system.
uses

    Quantity,
    Graphic2d,
    Aspect,
    PlotMgt,
    MMgt,
    TCollection,
    TColStd,
    Viewer

is

    class Viewer;
    private pointer ViewerPointer to Viewer from V2d;
    
    class View;
    ---Purpose: allows the creation of a view in a window driver.
    ---         describes all the commands available for a view.
    --          
    
    class DefaultMap;
    ---Purpose: furnishes default color, font, and width map.
    
    enumeration TypeOfWindowResizingEffect is TOWRE_ENLARGE_SPACE,
                                              TOWRE_ENLARGE_OBJECTS
    ---Purpose: determines the desired type of effect after the resizing
    --          of a window.
    end TypeOfWindowResizingEffect;

    ---Purpose: drawing of the grid.

    private class BackgroundGraphicObject;

    private class RectangularGrid;
    private class CircularGrid;

    private class CircularGraphicGrid;
    private class RectangularGraphicGrid;

    Draw(aViewer: Viewer from V2d);
    ---Purpose: Test

end V2d;
