-- File:	MakeScale.cdl
-- Created:	Mon Sep 28 11:53:08 1992
-- Author:	Remi GILET
--		<reg@sdsun2>
---Copyright:	 Matra Datavision 1992

class MakeScale

from GC

    ---Purpose: This class implements an elementary construction algorithm for
    -- a scaling transformation in 3D space. The result is a
    -- Geom_Transformation transformation.
    -- A MakeScale object provides a framework for:
    -- -   defining the construction of the transformation,
    -- -   implementing the construction algorithm, and
    -- -   consulting the result.
        
uses Pnt            from gp,
     Transformation from Geom,
     Real           from Standard
     
is

Create(Point : Pnt from gp      ;
       Scale : Real  from Standard) returns MakeScale;
    ---Purpose: Constructs a scaling transformation with
    -- -   Point as the center of the transformation, and
    -- -   Scale as the scale factor.       
    
Value(me) returns Transformation from Geom
    is static;
    ---Purpose: Returns the constructed transformation.
    ---C++: return const&

Operator(me) returns Transformation from Geom
    is static;
    ---C++: return const&
    ---C++: alias "Standard_EXPORT operator Handle_Geom_Transformation() const;"

fields

    TheScale : Transformation from Geom;

end MakeScale;

