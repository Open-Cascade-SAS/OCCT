-- Created on: 1993-03-10
-- Created by: JCV
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Direction from Geom inherits Vector from Geom

        ---Purpose :
        --  The class Direction specifies a vector that is never null.
        --  It is a unit vector.


uses  Dir      from gp,
      Pnt      from gp, 
      Trsf     from gp,
      Vec      from gp,
      Geometry from Geom

raises ConstructionError from Standard

is


  Create (X, Y, Z :Real)  returns Direction
        ---Purpose : Creates a unit vector with it 3 cartesian coordinates.
     raises ConstructionError;
        ---Purpose : 
        --  Raised if Sqrt( X*X + Y*Y + Z*Z) <= Resolution from gp.

  Create (V : Dir) returns Direction;
        ---Purpose : Creates a transient copy of <me>.


  SetCoord (me : mutable; X, Y, Z : Real)
        ---Purpose : Sets <me> to X,Y,Z coordinates.
     raises ConstructionError;
        ---Purpose : 
        --  Raised if Sqrt( X*X + Y*Y + Z*Z) <= Resolution from gp.


  SetDir (me : mutable; V : Dir);
        ---Purpose : Converts the gp_Dir unit vector V into this unit vector.


  SetX (me : mutable; X : Real)
        ---Purpose : Changes the X coordinate of <me>.
     raises ConstructionError;
        ---Purpose : 
        --  Raised if Sqrt( X*X + Y*Y + Z*Z) <= Resolution from gp.


  SetY (me : mutable; Y : Real)
        ---Purpose : Changes the Y coordinate of <me>.
     raises ConstructionError;
        ---Purpose : 
        --  Raised if Sqrt( X*X + Y*Y + Z*Z) <= Resolution from gp.


  SetZ (me : mutable; Z : Real)
        ---Purpose : Changes the Z coordinate of <me>.
     raises ConstructionError;
        ---Purpose : 
        --  Raised if Sqrt( X*X + Y*Y + Z*Z) <= Resolution from gp.


  Dir (me) returns Dir;
        ---Purpose :
        --  Returns the non transient direction with the same 
        --  coordinates as <me>.


  Magnitude (me)   returns Real;
        ---Purpose : returns 1.0 which is the magnitude of any unit vector.


  SquareMagnitude (me)   returns Real;
        ---Purpose : returns 1.0 which is the square magnitude of any unit vector.    
    
  Cross (me : mutable; Other : Vector)
        ---Purpose :
        --  Computes the cross product between <me> and <Other>.
     raises ConstructionError;
        ---Purpose :
        --  Raised if the two vectors are parallel because it is
        --  not possible to have a direction with null length.


  CrossCross (me : mutable; V1, V2 : Vector)
        ---Purpose :
        --  Computes the triple vector product  <me> ^(V1 ^ V2).
     raises ConstructionError;
        ---Purpose :
        --  Raised if V1 and V2 are parallel or <me> and (V1 ^ V2) are
        --  parallel


  Crossed (me; Other : Vector)  returns like me
        ---Purpose :
        --  Computes the cross product between <me> and <Other>.
        --  A new direction is returned.

     raises ConstructionError
        ---Purpose :
        --  Raised if the two vectors are parallel because it is 
        --  not possible to have a direction with null length.
     is static;
     

  CrossCrossed (me; V1, V2 : Vector)   returns like me
        ---Purpose :
        --  Computes the triple vector product <me> ^(V1 ^ V2).
     raises ConstructionError
        ---Purpose :
        --  Raised if V1 and V2 are parallel or <me> and (V1 ^ V2) are
        --  parallel
     is static;
 

  Transform (me : mutable; T : Trsf);
    	---Purpose: Applies the transformation T to this unit vector, then normalizes it.
  
  Copy (me) returns like me;
    	---Purpose: Creates a new object which is a copy of this unit vector.
end;

