-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ColourRgb from StepVisual 

inherits ColourSpecification from StepVisual 

uses

	Real from Standard, 
	HAsciiString from TCollection
is

	Create returns ColourRgb;
	---Purpose: Returns a ColourRgb


	Init (me : mutable;
	      aName : HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      aName : HAsciiString from TCollection;
	      aRed : Real from Standard;
	      aGreen : Real from Standard;
	      aBlue : Real from Standard) is virtual;

	-- Specific Methods for Field Data Access --

	SetRed(me : mutable; aRed : Real);
	Red (me) returns Real;
	SetGreen(me : mutable; aGreen : Real);
	Green (me) returns Real;
	SetBlue(me : mutable; aBlue : Real);
	Blue (me) returns Real;

fields

	red : Real from Standard;
	green : Real from Standard;
	blue : Real from Standard;

end ColourRgb;
