-- File:	Draw_Box.cdl
-- Created:	Fri Mar 10 14:18:31 1995
-- Author:	Remi LEQUETTE
--		<rle@phobox>
---Copyright:	 Matra Datavision 1995



class Box from Draw inherits Drawable3D from Draw

	---Purpose: 

uses Pnt from gp,
    Color from Draw,
    Display from Draw

is

    Create(p1,p2 : Pnt; col : Color)
    returns mutable Box;
    
    DrawOn(me; dis : in out Display);
    
    First(me) returns Pnt from gp
	---C++: return const&
    is static;

    First(me : mutable; P : Pnt from gp)
    is static;

    Last(me) returns Pnt from gp
	---C++: return const&
    is static;

    Last(me : mutable; P : Pnt from gp)
    is static;

fields

    myFirst : Pnt;
    myLast  : Pnt;
    myColor : Color;
    
end Box;
