-- Created by: DAUTRY Philippe
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

--      	--------------------

---Version:	0.0
--Version	Date		Purpose
--		0.0	Nov 27 1997	Creation

class TreeBrowser from DDataStd inherits Drawable3D from Draw

	---Purpose: Browses a TreeNode from TDataStd.
	--          =================================

uses

    Label               from TDF,
    TreeNode            from TDataStd,
    Interpretor         from Draw,
    Display             from Draw,
    AsciiString         from TCollection

is

    Create  (root : Label from TDF)
    returns TreeBrowser from DDataStd;
    
    DrawOn (me; dis : in out Display);
    
    Copy (me) 
    returns Drawable3D from Draw
    is redefined;

    Dump (me; S : in out OStream) 
    is redefined;

    Whatis (me; I : in out Interpretor from Draw)
    is redefined;

    ---Purpose: Specific methods
    --          ================

    Label (me : mutable; root : Label from TDF);
    
    Label (me) 
    returns Label from TDF;

    OpenRoot (me)
    ---Purpose: Returns   a   string composed with  the   TreeNode  of
    --          <myLabel>.
     returns AsciiString from TCollection;

    OpenNode (me; L : Label from TDF)
    ---Purpose:  Returns a string composed   with the sub-TreeNodes of
    --          <L>
    returns AsciiString from TCollection;

    OpenNode (me; aTreeNode :        TreeNode    from TDataStd;
    	    	  aList     : in out AsciiString from TCollection)  
    ---Purpose: Returns a string composed with the sub-TreeNodes
    --          of <aTreeNode>. Used to implement other methods.
    is private;

fields

    myRoot : Label from TDF;

end TreeBrowser;
