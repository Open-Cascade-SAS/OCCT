-- Created on: 1993-01-09
-- Created by: CKY / Contract Toubro-Larsen ( Kiran )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Direction from IGESGeom  inherits IGESEntity

        ---Purpose: defines IGESDirection, Type <123> Form <0>
        --          in package IGESGeom
        --          A direction entity is a non-zero vector in Euclidean 3-space
        --          that is defined by its three components (direction ratios)
        --          with respect to the coordinate axes. If x, y, z are the
        --          direction ratios then (x^2 + y^2 + z^2) > 0

uses

        Vec         from gp,
        XYZ         from gp

is

        Create returns mutable Direction;

        -- Specific Methods pertaining to the class

        Init (me : mutable; aDirection : XYZ);
        ---Purpose : This method is used to set the fields of the class
        --           Direction
        --       - aDirection : Direction ratios, Z is 0 by default

        Value (me) returns Vec;

        TransformedValue (me) returns Vec;
        ---Purpose : returns the Direction value after applying Transformation matrix

fields

--
-- Class    : IGESGeom_Direction
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class Direction.
--
-- Reminder : A Direction instance is defined by :
--            The three direction ratios along the three coordinate axes

        theDirection : XYZ;

end Direction;
