-- File:	IGESAppli_ToolPartNumber.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolPartNumber  from IGESAppli

    ---Purpose : Tool to work on a PartNumber. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses PartNumber from IGESAppli,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolPartNumber;
    ---Purpose : Returns a ToolPartNumber, ready to work


    ReadOwnParams (me; ent : mutable PartNumber;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : PartNumber;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : PartNumber;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a PartNumber <ent>, from
    --           its specific (own) parameters

    OwnCorrect (me; ent : mutable PartNumber) returns Boolean  is static;
    ---Purpose : Sets automatic unambiguous Correction on a PartNumber
    --           (NbPropertyValues forced to 4)

    DirChecker (me; ent : PartNumber) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : PartNumber;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : PartNumber; entto : mutable PartNumber;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : PartNumber;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolPartNumber;
