-- Created by: Peter KURNEV
-- Copyright (c) 2010-2012 OPEN CASCADE SAS
-- Copyright (c) 2007-2010 CEA/DEN, EDF R&D, OPEN CASCADE
-- Copyright (c) 2003-2007 OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN, CEDRAT,
--                         EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class BuilderFace from BOPAlgo 
    	inherits BuilderArea from BOPAlgo 
	 
	---Purpose: The algorithm to build faces from set of edges  

uses    
    Orientation from TopAbs,
    Face from TopoDS,
    BaseAllocator from BOPCol 
--raises

is 
    Create  
    	returns BuilderFace from BOPAlgo; 
    ---C++: alias "Standard_EXPORT virtual ~BOPAlgo_BuilderFace();" 
      
    Create (theAllocator: BaseAllocator from BOPCol)  
    	returns BuilderFace from BOPAlgo;  
	
    SetFace(me:out; 
            theFace:Face from TopoDS);  
    ---Purpose: Sets the face generatix  
	 
    Face(me) 
    ---Purpose: Returns the face generatix   
    	returns Face from TopoDS; 
    ---C++:  return const &
		 
    Perform(me:out)  
    	---Purpose:  Performs the algorithm 
    	is redefined;  
	 
    PerformShapesToAvoid(me:out) 
	---Purpose:  Collect the edges that 
	--           a) are internal        	 
	--           b) are the same and have different orientation         	 
    	is redefined protected; 
	 
    PerformLoops(me:out) 
	---Purpose: Build draft wires 
        --          a)myLoops - draft wires that consist of  
        --                       boundary edges 
	--          b)myLoopsInternal - draft wires that contains 
	--                               inner edges 
    	is redefined protected;  
	 
    PerformAreas(me:out)   
    	---Purpose: Build draft faces that contains boundary edges 
    	is redefined protected;  

    PerformInternalShapes(me:out)   
    	---Purpose: Build finalized faces with internals   
    	is redefined protected;  
     
    CheckData(me:out) 
	is redefined protected;   
     
    Orientation(me) 
    	returns Orientation from TopAbs; 
 
fields  
    myFace : Face from TopoDS is protected;     
    myOrientation: Orientation from TopAbs is protected;   	      
 
end BuilderFace; 

