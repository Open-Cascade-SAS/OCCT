-- File:	StepToGeom_MakeParabola2d.cdl
-- Created:	Tue May  9 10:42:44 1995
-- Author:	Dieter THIEMANN
---Copyright:	 Matra Datavision 1994

class MakeParabola2d from StepToGeom

    ---Purpose: This class implements the mapping between classes 
    --          Parabola from StepGeom which describes a Parabola from
    --          Prostep and Parabola from Geom2d.

uses 
     Parabola from Geom2d,
     Parabola from StepGeom

is

    Convert ( myclass; SC : Parabola from StepGeom;
                       CC : out Parabola from Geom2d )
    returns Boolean from Standard;

end MakeParabola2d;
