-- Created on: 1997-07-29
-- Created by: Denis PASCAL 
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- modified     Sergey Zaritchny


class Constraint from PDataXtd inherits Attribute from PDF

	---Purpose: 

uses Integer          from Standard,
     Real             from PDataStd,
     HAttributeArray1 from PDF,
     NamedShape       from PNaming
    
is

    Create returns mutable Constraint from  PDataXtd;
    
    
    Create (Type        : Integer          from Standard;
    	    Geometries  : HAttributeArray1 from PDF;
    	    Value       : Real             from PDataStd;
    	    Plane       : NamedShape       from PNaming) 
    returns mutable Constraint from PDataXtd;
    
    
    GetValue (me) returns Real from PDataStd;
    

    GetType (me) returns Integer from Standard;
    
    
    GetGeometries (me) returns HAttributeArray1 from PDF;
    
    
    Set (me : mutable; V : Real from PDataStd);


    SetType (me : mutable; Type : Integer from Standard);
    
    
    SetGeometries (me : mutable; Geometries : HAttributeArray1 from PDF);
    
    SetPlane (me : mutable; plane : NamedShape from PNaming);
    GetPlane (me)
    returns NamedShape from PNaming;
    
    Verified(me:mutable; status : Boolean from Standard);
    Verified(me) 
    returns Boolean from Standard;    

    Inverted(me:mutable; status : Boolean from Standard);
    Inverted(me) 
    returns Boolean from Standard;    

    Reversed(me:mutable; status : Boolean from Standard);
    Reversed(me) 
    returns Boolean from Standard;    
    
fields

    myType       : Integer          from Standard;
    myGeometries : HAttributeArray1 from PDF;
    myValue      : Real             from PDataStd;
    myIsReversed : Boolean          from Standard;
    myIsInverted : Boolean          from Standard;
    myIsVerified : Boolean          from Standard;
    myPlane      : NamedShape       from PNaming;
    
end Constraint;
