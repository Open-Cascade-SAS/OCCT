-- Created on: 1995-06-12
-- Created by: Joelle CHAUVET
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Modified:	Tue Oct 15 10:12:02 1996
--              Add ChFi2d_TangencyError (PRO3529)
-- Modified:	Tue Oct 22 09:23:11 1996
--		Add ChFi2d_FirstEdgeDegenerated, ChFi2d_LastEdgeDegenerated,
--		ChFi2d_BothEdgesDegenerated (PRO4896)
-- Modified:	Fri Sep 25 09:38:04 1998
--              ChFi2d_NotAuthorized is used if the edges are not
--              lines or circles (BUC60288)

package ChFi2d 

	---Purpose: This package contains the algorithms used to build
	--          fillets or chamfers on planar wire.
	--
	-- This package provides two algorithms for 2D fillets:
	--     ChFi2d_Builder - it constructs a fillet or chamfer 
	--                      for linear and circular edges of a face.
	--     ChFi2d_FilletAPI - it encapsulates two algorithms:
	--         ChFi2d_AnaFilletAlgo - analytical constructor of the fillet.
	--                                It works only for linear and circular edges,
	--                                having a common point.
	--         ChFi2d_FilletAlgo - iteration recursive method constructing 
	--                             the fillet edge for any type of edges including
	--                             ellipses and b-splines. 
	--                             The edges may even have no common point.
	--     ChFi2d_ChamferAPI - an algoroithm for construction of chamfers 
	--                         between two linear edges of a plane.
	--
	-- The algorithms ChFi2d_AnaFilletAlgo and ChFi2d_FilletAlgo may be used directly 
	-- or via the interface class ChFi2d_FilletAPI.

uses
    TopoDS,
    TopTools,
    gp

is
    
    enumeration ConstructionError is
	---Purpose: error     that    can   occur       during   the
	--          fillet  construction on planar wire
	NotPlanar,
	    ---Purpose: the face is not planar
	NoFace,
	    ---Purpose: the face is null
    	InitialisationError,
	    ---Purpose: the two  faces used for the initialisation are
	    --          uncompatible.
	ParametersError,
	    ---Purpose: the  parameters  as  distances   or  angle for
	    --          chamfer are less or equal to zero.
    	Ready,
	    ---Purpose: the initialization has been succesfull.
	IsDone,
	ComputationError,
	    ---Purpose: the algorithm could not find a solution.
	ConnexionError,
	    ---Purpose: the vertex given  to locate the fillet  or the
	    --          chamfer  is not connected to 2 edges.
	TangencyError,
	    ---Purpose: the two edges connected to the vertex are tangent.

 
	FirstEdgeDegenerated,
	    ---Purpose: the first edge is degenerated.
	LastEdgeDegenerated,
	    ---Purpose: the last edge is degenerated.
	BothEdgesDegenerated,
	    ---Purpose: the two edges are degenerated.
    	NotAuthorized
	    ---Purpose: One or the two  edges connected to the  vertex
	    --          is a fillet or a chamfer
	    --          One or the two  edges connected to the  vertex
	    --          is not a line or a circle
	
    end ConstructionError;


    class Builder;


    CommonVertex( E1, E2 :     Edge   from TopoDS; 
    	    	  V      : out Vertex from TopoDS)
    returns Boolean
    is private;
    	---Warning: <V> has sense only if the value <True> is returned    


    FindConnectedEdges( F      :     Face   from TopoDS;
    	    	        V      :     Vertex from TopoDS;
    	    	        E1, E2 : out Edge   from TopoDS)
    returns ConstructionError from ChFi2d
    is private;

    	---Warning: <E1> and <E2> has sense only if the returned value
    	--          is <IsDone>


end ChFi2d;






