-- Created on: 1991-01-14
-- Created by: Arnaud BOUZY
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class SingleRelation from Expr

inherits GeneralRelation from Expr

uses GeneralExpression from Expr,
    NamedUnknown from Expr,
    AsciiString from TCollection

raises OutOfRange

is

    SetFirstMember(me :mutable; exp : GeneralExpression)
    ---Purpose: Defines the first member of the relation
    ---Level : Internal
    is static;
    
    SetSecondMember(me :mutable; exp : GeneralExpression)
    ---Purpose: Defines the second member of the relation
    ---Level : Internal
    is static;
    
    FirstMember(me)
    ---Purpose: Returns the first member of the relation
    ---Level : Internal
    returns GeneralExpression
    is static;

    SecondMember(me)
    ---Purpose: Returns the second member of the relation
    ---Level : Internal
    returns GeneralExpression
    is static;

    IsLinear(me)
    ---Purpose: Tests if <me> is linear between its NamedUnknowns.
    returns Boolean
    is static;

    NbOfSubRelations(me)
    ---Purpose: Returns the number of relations contained in <me>.
    returns Integer
    is static;
    
    NbOfSingleRelations(me)
    ---Purpose: Returns the number of SingleRelations contained in 
    --          <me> (Always 1).
    returns Integer
    is static;

    SubRelation(me; index : Integer)
    ---Purpose: Returns the relation denoted by <index> in <me>.
    --          An exception is raised if index is out of range.
    returns any GeneralRelation
    raises OutOfRange
    is static;

    Contains(me; exp : GeneralExpression)
    ---Purpose: Tests if <me> contains <exp>.
    returns Boolean;
    
    Replace(me : mutable ; var : NamedUnknown ; with : GeneralExpression);
    ---Purpose: Replaces all occurences of <var> with <with> in <me>.
    
fields

    myFirstMember : GeneralExpression;
    mySecondMember : GeneralExpression;

end SingleRelation;
