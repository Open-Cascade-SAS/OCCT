-- Created by: DAUTRY Philippe
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

--      	-------

---Version:	0.0
--Version	Date		Purpose
--		0.0	Mar 13 1997	Creation


package PDF 

	---Purpose: This pakage is the persistent equivalent of
	--          TDF. It describes persistent classes used to store
	--          a TDF structure into a Database.


uses

    Standard,
    PCollection,
    PColStd

is

    class Data;
    
    
    deferred class Attribute;

    class TagSource; 

    class Reference;

    -- Instantiations ---------------------------------------------------

    class HAttributeArray1 from PDF instantiates HArray1 from PCollection
    	(Attribute from PDF);

end PDF;
