-- Created on: 2000-10-05
-- Created by: Andrey BETENEV
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ActorWrite from STEPCAFControl inherits ActorWrite from STEPControl

    ---Purpose: Extends ActorWrite from STEPControl by analysis of
    --          whether shape is assembly (based on information from DECAF)

uses
    Shape from TopoDS,
    MapOfShape from TopTools

is

    Create returns ActorWrite;

    IsAssembly (me; S: in out Shape from TopoDS) returns Boolean is redefined;
    	---Purpose: Check whether shape S is assembly
	--          Returns True if shape is registered in assemblies map

    SetStdMode (me: mutable; stdmode: Boolean = Standard_True);
    	---Purpose: Set standard mode of work 
	--          In standard mode Actor (default) behaves exactly as its 
        --          ancestor, also map is cleared

    ClearMap (me: mutable);
    	---Purpose: Clears map of shapes registered as assemblies

    RegisterAssembly (me: mutable; S: Shape from TopoDS);
    	---Purpose: Registers shape to be written as assembly
	--          The shape should be TopoDS_Compound (else does nothing)

fields

    myStdMode: Boolean;
    myMap: MapOfShape from TopTools;

end ActorWrite;
