-- Created on: 1993-01-11
-- Created by: CKY / Contract Toubro-Larsen ( Anand NATRAJAN )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class PWBArtworkStackup from IGESAppli  inherits IGESEntity

        ---Purpose: defines PWBArtworkStackup, Type <406> Form <25>
        --          in package IGESAppli
        --          Used to communicate which exchange file levels are to
        --          be combined in order to create the artwork for a
        --          printed wire board (PWB). This property should be
        --          attached to the entity defining the printed wire
        --          assembly (PWA) or if no such entity exists, then the
        --          property should stand alone in the file.

uses

        HAsciiString from TCollection,
        HArray1OfInteger from TColStd

raises OutOfRange

is

        Create returns mutable PWBArtworkStackup;

        -- Specific Methods pertaining to the class

        Init (me           : mutable;
              nbPropVal    : Integer;
              anArtIdent   : HAsciiString;
              allLevelNums : HArray1OfInteger);
        ---Purpose : This method is used to set the fields of the class
        --           PWBArtworkStackup
        --       - nbPropVal    : number of property values
        --       - anArtIdent   : Artwork Stackup Identification
        --       - allLevelNums : Level Numbers

        NbPropertyValues (me) returns Integer;
        ---Purpose : returns number of property values

        Identification (me) returns HAsciiString from TCollection;
        ---Purpose : returns Artwork Stackup Identification

        NbLevelNumbers (me) returns Integer;
        ---Purpose : returns total number of Level Numbers

        LevelNumber (me; Index : Integer) returns Integer
        raises OutOfRange;
        ---Purpose : returns Level Number
        -- raises exception if Index <= 0 or Index > NbLevelNumbers

fields

--
-- Class    : IGESAppli_PWBArtworkStackup
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class PWBArtworkStackup.
--
-- Reminder : A PWBArtworkStackup instance is defined by :
--            - number of property values
--            - Artwork Stackup Identification string
--            - Level Numbers

        theNbPropertyValues    : Integer;
        theArtworkStackupIdent : HAsciiString;
        theLevelNumbers        : HArray1OfInteger;

end PWBArtworkStackup;
