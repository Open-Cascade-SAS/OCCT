-- Created on: 1991-02-21
-- Created by: Isabelle GRIGNON
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

generic class   Point from Extrema  (Pnt as any)
        inherits Storable from Standard
    	---Purpose: Definition of a point on curve.


is
    Create returns Point;
    	---Purpose: Creation of an indefinite point on curve.

    Create (U: Real; P: Pnt) returns Point;
    	---Purpose: Creation of a point on curve with a parameter 
    	--          value on the curve and a Pnt from gp.

    SetValues(me: in out; U: Real; P: Pnt)
    	---Purpose: sets the point and parameter values.
    is static;

    Value (me) returns Pnt
    	---Purpose: Returns the point.
    	---C++: return const&
    	---C++: inline
    	is static;

    Parameter (me) returns Real
    	---Purpose: Returns the parameter on the curve.
    	---C++: inline
    	is static;

fields
    myU: Real;
    myP: Pnt;

end Point;
