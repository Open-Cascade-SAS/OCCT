-- Created on: 1994-03-18
-- Created by: Yves FRICAUD
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class Curve from Bisector 

	---Purpose: 

inherits
    Curve from Geom2d

uses
    Pnt2d from gp

is
    
    Parameter ( me ; P : Pnt2d from gp) returns Real
    is deferred;
    
    IsExtendAtStart (me) returns Boolean from Standard
    is deferred;
    
    IsExtendAtEnd   (me) returns Boolean from Standard
    is deferred;

    NbIntervals (me) returns Integer
	---Purpose: If necessary,  breaks the  curve in  intervals  of
	--          continuity  <C1>.    And  returns   the number   of
	--          intervals.
    is deferred;

    IntervalFirst(me; Index : Integer from Standard) returns Real
       ---Purpose: Returns  the  first  parameter    of  the  current
       --          interval. 
    is deferred;
    
    IntervalLast(me; Index : Integer from Standard) returns Real
       ---Purpose: Returns  the  last  parameter    of  the  current
       --          interval. 
    is deferred;
    
end Curve;



