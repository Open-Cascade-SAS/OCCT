-- Created on: 1997-02-10
-- Created by: Alexander BRIVIN
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Info from Vrml 

	---Purpose:  defines a Info node of VRML specifying properties of geometry
	---          and its appearance. 
    	--  It  is  used  to  store  information  in  the  scene  graph, 
	--  Typically  for  application-specific  purposes,  copyright  messages, 
	--  or  other  strings.
uses

     AsciiString from TCollection
is
 
    Create  (  aString  :  AsciiString from TCollection  =  "<Undefined info>")    
        returns Info from Vrml; 

    SetString ( me : in out;  aString  :  AsciiString from TCollection ); 
    String ( me  )  returns  AsciiString from TCollection; 
   
    Print  ( me;  anOStream: in out OStream from Standard ) returns OStream from Standard;
    ---C++:  return  & 

fields
 
    myString  :  AsciiString from TCollection;  -- Info string

end Info;

