-- Created on: 1991-04-12
-- Created by: Michel CHAUVAT
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

--		Jean-Claude VAUTHIER January 1992


generic class VGProps from GProp (Arc as any;
                                  Face as any;  -- as FaceTool(Arc)
    	    	    	    	  Domain as any -- as DomainTool(Arc)
    	    	    	    	 )
inherits GProps

        --- Purpose :
        --  Computes the global properties of a geometric solid 
        --  (3D closed region of space) delimited with :
        --  . a surface
        --  . a point and a surface
        --  . a plane and a surface
        --  
        --  The surface can be :
        --  . a surface limited with its parametric values U-V,
        --  . a surface limited in U-V space with its curves of restriction,
        --  
        --  The surface 's requirements to evaluate the global properties
        --  are defined in the template SurfaceTool from package GProp.

uses   	Pnt      from gp,
        Pln      from gp
is

  Create returns VGProps;
  
  Create (S: Face; VLocation: Pnt from gp) returns VGProps;
        --- Purpose : 
        --  Computes the global properties of a region of 3D space
        --  delimited with the surface <S> and the point VLocation. S can be closed 
	--  The method is quick and its precision is enough for many cases of analytical 
    	--  surfaces. 
        --  Non-adaptive 2D Gauss integration with predefined numbers of Gauss points 
	--  is used. Numbers of points depend on types of surfaces and  curves.
    	--  Errror of the computation is not calculated. 
	
  Create (S: in out Face; VLocation: Pnt from gp; Eps: Real) returns VGProps; 
        --- Purpose : 
        --  Computes the global properties of a region of 3D space
        --  delimited with the surface <S> and the point VLocation. S can be closed 
	--  Adaptive 2D Gauss integration is used. 
	--  Parameter Eps sets maximal relative error of computed mass (volume) for face. 
	--  Error is calculated as Abs((M(i+1)-M(i))/M(i+1)), M(i+1) and M(i) are values 
	--  for two successive steps of adaptive integration. 

  Create (S: Face; O: Pnt from gp; VLocation: Pnt from gp) returns VGProps;
        --- Purpose :  
        --  Computes the global properties of the region of 3D space
        --  delimited with the surface <S> and the point VLocation.
	--  The method is quick and its precision is enough for many cases of analytical 
    	--  surfaces. 
        --  Non-adaptive 2D Gauss integration with predefined numbers of Gauss points 
	--  is used. Numbers of points depend on types of surfaces and  curves.
    	--  Error of the computation is not calculated. 
	
  Create (S: in out Face; O: Pnt from gp; VLocation: Pnt from gp; Eps: Real) returns VGProps;
        --- Purpose :  
        --  Computes the global properties of the region of 3D space
        --  delimited with the surface <S> and the point VLocation.
	--  Adaptive 2D Gauss integration is used. 
	--  Parameter Eps sets maximal relative error of computed mass (volume) for face. 
	--  Error is calculated as Abs((M(i+1)-M(i))/M(i+1)), M(i+1) and M(i) are values 
	--  for two successive steps of adaptive integration. 
	--          WARNING: if Eps > 0.001 algorithm performs non-adaptive integration.	  
     
  Create (S: Face; Pl: Pln from gp; VLocation: Pnt from gp) returns VGProps;
        --- Purpose :  
        --  Computes the global properties of the region of 3D space
        --  delimited with the surface <S> and the plane Pln.
	--  The method is quick and its precision is enough for many cases of analytical 
    	--  surfaces.  
        --  Non-adaptive 2D Gauss integration with predefined numbers of Gauss points 
	--  is used. Numbers of points depend on types of surfaces and  curves.
    	--  Error of the computation is not calculated. 
	
  Create (S: in out Face; Pl: Pln from gp; VLocation: Pnt from gp; Eps: Real) returns VGProps;
        --- Purpose :  
        --  Computes the global properties of the region of 3D space
        --  delimited with the surface <S> and the plane Pln.
	--  Adaptive 2D Gauss integration is used. 
	--  Parameter Eps sets maximal relative error of computed mass (volume) for face. 
	--  Error is calculated as Abs((M(i+1)-M(i))/M(i+1)), M(i+1) and M(i) are values 
	--  for two successive steps of adaptive integration. 
	--          WARNING: if Eps > 0.001 algorithm performs non-adaptive integration.	  

    	--  With  Domain  -- 

  Create (S: in out Face; D : in out Domain; VLocation: Pnt from gp) returns VGProps;
        --- Purpose : 
        --  Computes the global properties of a region of 3D space
        --  delimited with the surface <S> and the point VLocation. S can be closed 
	--  The method is quick and its precision is enough for many cases of analytical 
    	--  surfaces. 
        --  Non-adaptive 2D Gauss integration with predefined numbers of Gauss points 
	--  is used. Numbers of points depend on types of surfaces and  curves.
    	--  Errror of the computation is not calculated. 
	
  Create (S: in out Face; D : in out Domain; VLocation: Pnt from gp; Eps: Real) returns VGProps; 
        --- Purpose : 
        --  Computes the global properties of a region of 3D space
        --  delimited with the surface <S> and the point VLocation. S can be closed 
	--  Adaptive 2D Gauss integration is used. 
	--  Parameter Eps sets maximal relative error of computed mass (volume) for face. 
	--  Error is calculated as Abs((M(i+1)-M(i))/M(i+1)), M(i+1) and M(i) are values 
	--  for two successive steps of adaptive integration. 

  Create (S: in out Face; D : in out Domain; O: Pnt from gp; VLocation: Pnt from gp) returns VGProps;
        --- Purpose :  
        --  Computes the global properties of the region of 3D space
        --  delimited with the surface <S> and the point VLocation.
	--  The method is quick and its precision is enough for many cases of analytical 
    	--  surfaces. 
        --  Non-adaptive 2D Gauss integration with predefined numbers of Gauss points 
	--  is used. Numbers of points depend on types of surfaces and  curves.
    	--  Error of the computation is not calculated. 
	
  Create (S: in out Face; D : in out Domain; O: Pnt from gp; VLocation: Pnt from gp; Eps: Real) returns VGProps;
        --- Purpose :  
        --  Computes the global properties of the region of 3D space
        --  delimited with the surface <S> and the point VLocation.
	--  Adaptive 2D Gauss integration is used. 
	--  Parameter Eps sets maximal relative error of computed mass (volume) for face. 
	--  Error is calculated as Abs((M(i+1)-M(i))/M(i+1)), M(i+1) and M(i) are values 
	--  for two successive steps of adaptive integration. 
	--          WARNING: if Eps > 0.001 algorithm performs non-adaptive integration.	  
     
  Create (S: in out Face; D : in out Domain; Pl: Pln from gp; VLocation: Pnt from gp) returns VGProps;
        --- Purpose :  
        --  Computes the global properties of the region of 3D space
        --  delimited with the surface <S> and the plane Pln.
	--  The method is quick and its precision is enough for many cases of analytical 
    	--  surfaces.  
        --  Non-adaptive 2D Gauss integration with predefined numbers of Gauss points 
	--  is used. Numbers of points depend on types of surfaces and  curves.
    	--  Error of the computation is not calculated. 
	
  Create (S: in out Face; D : in out Domain; Pl: Pln from gp; VLocation: Pnt from gp; Eps: Real) returns VGProps;
        --- Purpose :  
        --  Computes the global properties of the region of 3D space
        --  delimited with the surface <S> and the plane Pln.
	--  Adaptive 2D Gauss integration is used. 
	--  Parameter Eps sets maximal relative error of computed mass (volume) for face. 
	--  Error is calculated as Abs((M(i+1)-M(i))/M(i+1)), M(i+1) and M(i) are values 
	--  for two successive steps of adaptive integration. 
	--          WARNING: if Eps > 0.001 algorithm performs non-adaptive integration.	  

  SetLocation(me: in out; VLocation: Pnt from gp);
  
  Perform(me: in out; S: Face);
  Perform(me: in out; S: in out Face; Eps: Real) returns Real;

  Perform(me: in out; S: Face; O : Pnt from gp);
  Perform(me: in out; S: in out Face; O : Pnt from gp; Eps: Real) returns Real;

  Perform(me: in out; S: Face; Pl : Pln from gp);
  Perform(me: in out; S: in out Face; Pl : Pln from gp; Eps: Real) returns Real;

  Perform(me: in out; S: in out  Face; D : in out Domain);
  Perform(me: in out; S: in out Face; D : in out Domain;  Eps: Real) returns Real;

  Perform(me: in out; S: in out Face; D : in out Domain;  O : Pnt from gp);
  Perform(me: in out; S: in out Face; D : in out Domain;  O : Pnt from gp; Eps: Real) returns Real;

  Perform(me: in out; S: in out Face; D : in out Domain;  Pl : Pln from gp);
  Perform(me: in out; S: in out Face; D : in out Domain;  Pl : Pln from gp; Eps: Real) returns Real;

  GetEpsilon(me: out) returns Real;
        --- Purpose :  
        --  If previously used methods containe Eps parameter  
    	--  gets actual relative error of the computation, else returns  1.0.
fields
 
    myEpsilon: Real from Standard;

end VGProps;


