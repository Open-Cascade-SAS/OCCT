-- Created on: 1993-03-02
-- Created by: Philippe DAUTRY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class BezierSurface from PGeom inherits BoundedSurface from PGeom

        ---Purpose :   Defines a  rational  or  non  rational   Bezier
        --         surface.  In this package the  degree of the Bezier
        --         surface is limited to MaxDegree and must be greater
        --         or equal to 1.
        --         
	---See Also : BezierSurface from Geom.

uses HArray2OfReal from PColStd,
     HArray2OfPnt  from PColgp

is


  Create returns mutable BezierSurface from PGeom;
	---Purpose: Creates a BezierSurface with default values.
    	---Level: Internal 


  Create (aURational : Boolean from Standard;
    	  aVRational : Boolean from Standard;
    	  aPoles     : HArray2OfPnt from PColgp;
    	  aWeights   : HArray2OfReal from PColStd)
     returns mutable BezierSurface from PGeom;
	---Purpose: Creates a BezierSurface with these values.
    	---Level: Internal 


  Poles (me: mutable; aPoles: HArray2OfPnt from PColgp);
	---Purpose: Set the field poles with <aPoles>.
    	---Level: Internal 



  Poles (me) returns HArray2OfPnt from PColgp;
	---Purpose: Returns the value of the field poles.
    	---Level: Internal 


  Weights (me: mutable; aWeights : HArray2OfReal from PColStd);
        ---Purpose : Set the value of the field weights with <aWeights>.
    	---Level: Internal 

  
  Weights (me) returns HArray2OfReal from PColStd;
        ---Purpose : Returns the value of the field weights.
    	---Level: Internal 

  
  URational (me: mutable; aURational: Boolean from Standard);
        ---Purpose : Set the value of the field uRational with <aURational>.
    	---Level: Internal 


  URational (me) returns Boolean from Standard;
        ---Purpose : Returns the value of the field uRational.
    	---Level: Internal 


  VRational (me: mutable; aVRational: Boolean from Standard);
        ---Purpose : Set the value of the field vRational with <aVRational>.
    	---Level: Internal 


  VRational (me) returns Boolean from Standard;
        ---Purpose : Returns the value of the field vRational.
    	---Level: Internal 



fields

   uRational : Boolean from Standard;
   vRational : Boolean from Standard;
   poles     : HArray2OfPnt from PColgp;
   weights   : HArray2OfReal from PColStd;

end;
