-- Created on: 1996-05-28
-- Created by: Denis PASCAL
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Angle from DrawDim inherits Dimension from DrawDim

	---Purpose: 

uses Face    from TopoDS,
     Display from Draw

is

    Create (plane1 : Face from TopoDS; 
            plane2 : Face from TopoDS)
    returns mutable Angle from DrawDim;
    
    Plane1 (me) returns Face from TopoDS;
	---C++: return const&

    Plane1 (me : mutable; plane : Face from TopoDS);

    Plane2  (me) returns Face from TopoDS;
	---C++: return const&

    Plane2 (me : mutable; plane : Face from TopoDS);    

    DrawOn (me; dis : in out Display);
    
fields

    myPlane1 : Face from TopoDS;
    myPlane2 : Face from TopoDS;
    
end Angle;

