-- Created on: 1996-01-22
-- Created by: Philippe MANGIN
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



deferred class DistributionOfEnergy from  FairCurve 
     inherits  FunctionSet from math

	---Purpose: Abstract class to use the Energy of an FairCurve

uses  Vector        from math, 
      FunctionSet   from math,
      HArray1OfReal  from TColStd,
      HArray1OfPnt2d from TColgp   



is

---    redefined methods

    NbVariables(me)
    	---Purpose: returns the number of variables of the function.

    returns Integer is redefined;

    
    NbEquations(me)
    	---Purpose: returns the number of equations of the function.

    returns Integer is redefined;

    
---    new methods
    Initialize( BSplOrder : Integer;
                FlatKnots :  HArray1OfReal;
		Poles     :  HArray1OfPnt2d;
    	    	DerivativeOrder : Integer;
    	    	NbValAux  : Integer = 0);
		
    SetDerivativeOrder(me :in out; DerivativeOrder : Integer); 
		    

fields

MyBSplOrder   : Integer is protected;
MyFlatKnots   : HArray1OfReal is  protected;
MyPoles       : HArray1OfPnt2d  is protected;
MyDerivativeOrder : Integer is protected;
MyNbVar       : Integer is protected;
MyNbEqua      : Integer is protected;
MyNbValAux    : Integer is protected;


end DistributionOfEnergy ;
