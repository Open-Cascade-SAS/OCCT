-- File:	Parab2d.cdl
-- Created:	Wed Aug 26 14:31:48 1992
-- Author:	Remi GILET
--		<reg@topsn3>
---Copyright:	 Matra Datavision 1992

class MakeParab2d from gce inherits Root from gce

    ---Purpose :This class implements the following algorithms used to 
    --          create Parab2d from gp.
    --  Defines an infinite parabola.
    --  An axis placement one axis defines the local cartesian
    --  coordinate system ("XAxis") of the parabola.
    --  The vertex of the parabola is the "Location" point of the 
    --  local coordinate system of the parabola. 
    --  The "XAxis" of the parabola is its axis of symmetry.
    --  The "XAxis" is oriented from the vertex of the parabola to the 
    --  Focus of the parabola.
    --  The "YAxis" is parallel to the directrix of the parabola and
    --  its "Location" point is the vertex of the parabola.
    --  The equation of the parabola in the local coordinate system is
    --  Y**2 = (2*P) * X
    --  P is the distance between the focus and the directrix of the 
    --  parabola called Parameter). 
    --  The focal length F = P/2 is the distance between the vertex 
    --  and the focus of the parabola.
    --          
    --          * Create a Parab2d from one apex  and the center.
    --          * Create a Parab2d with the directrix and the focus point.
    --          * Create a Parab2d with its vertex point and its axis 
    --            of symetry and its focus length.

uses Pnt2d   from gp,
     Ax2d    from gp,
     Ax22d   from gp,
     Parab2d from gp

raises NotDone from StdFail

is

Create (MirrorAxis : Ax2d    from gp                      ; 
    	Focal      : Real    from Standard                ;
    	Sense      : Boolean from Standard = Standard_True) 
    returns MakeParab2d;
    --- Purpose :
    --  Creates a parabola with its axis of symmetry ("MirrorAxis") 
    --  and its focal length.
    --- Warnings : It is possible to have Focal = 0.
    --  The status is "NullFocalLength" Raised if Focal < 0.0

Create (A     : Ax22d   from gp       ; 
    	Focal : Real    from Standard ) 
    returns MakeParab2d;
    --- Purpose :
    --  Creates a parabola with its local coordinate system <A> 
    --  and its focal length.
    --- Warnings : It is possible to have Focal = 0.
    --  The status is "NullFocalLength" Raised if Focal < 0.0

Create (D     : Ax2d  from gp                        ; 
    	F     : Pnt2d from gp                        ;
    	Sense : Boolean from Standard = Standard_True)  
    returns MakeParab2d;
    --- Purpose :
    --  Creates a parabola with the directrix and the focus point.
    --  The sense of parametrization is given by Sense.

Create (D     : Ax22d from gp  ; 
    	F     : Pnt2d from gp  )  
    returns MakeParab2d;
    --- Purpose :
    --  Creates a parabola with the local coordinate system and 
    --  the focus point.
    --  The sense of parametrization is given by Sense.

Create(S1     : Pnt2d   from gp                      ;
       Center : Pnt2d   from gp                      ;
    	Sense : Boolean from Standard = Standard_True) returns MakeParab2d;
    ---Purpose: Make an Parab2d with S1 as the Focal point and Center
    --          as the apex of the parabola
    --	Warning
    -- The MakeParab2d class does not prevent the
    -- construction of a parabola with a null focal distance.
    -- If an error occurs (that is, when IsDone returns
    -- false), the Status function returns:
    -- -   gce_NullFocusLength if Focal is less than 0.0, or
    -- -   gce_NullAxis if S1 and Center are coincident.
        
Value(me) returns Parab2d from gp
    raises NotDone
    is static;
    ---C++: return const&
    ---Purpose: Returns the constructed parabola.
    -- Exceptions StdFail_NotDone if no parabola is constructed.
    
Operator(me) returns Parab2d from gp
    is static;
    ---C++: return const&
    ---C++: alias "Standard_EXPORT operator gp_Parab2d() const;"

fields

    TheParab2d : Parab2d from gp;
    --The solution from gp.
    
end MakeParab2d;




