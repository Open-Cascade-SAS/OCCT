-- File:	Adaptor3d_HVertex.cdl
-- Created:	Fri Mar 25 12:31:39 1994
-- Author:	model
--		<model@topsn2>
---Copyright:	 Matra Datavision 1994


class HVertex from Adaptor3d 

	---Purpose: 


inherits TShared from MMgt

uses Pnt2d       from gp,
     Orientation from TopAbs,
     HCurve2d    from Adaptor2d

is

    Create
    
    	returns mutable HVertex from Adaptor3d;


    Create(P: Pnt2d from gp; Ori: Orientation from TopAbs;
           Resolution: Real from Standard)

    	returns mutable HVertex from Adaptor3d;


    Value(me: mutable)
    
    	returns Pnt2d from gp
    is virtual;


    Parameter(me: mutable; C: HCurve2d from Adaptor2d)
    
    	returns Real from Standard
    is virtual;


    Resolution(me: mutable; C: HCurve2d from Adaptor2d)
    
	---Purpose: Parametric resolution (2d).

    	returns Real from Standard
    is virtual;


    Orientation(me: mutable)
    
    	returns Orientation from TopAbs
    is virtual;


    IsSame(me: mutable; Other: mutable like me)
    
    	returns Boolean from Standard
    is virtual;


fields

    myPnt : Pnt2d       from gp;
    myTol : Real        from Standard;
    myOri : Orientation from TopAbs;

end HVertex;
