-- Created on: 2009-04-06
-- Created by: Sergey ZARITCHNY
-- Copyright (c) 2009-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class Pattern from TDataXtd inherits Attribute from TDF

	---Purpose: a general pattern model

uses 
     Array1OfTrsf from TDataXtd,
     LabelList    from TDF,
     GUID         from Standard

is

    GetID (myclass)   
    ---C++: return const &  
    returns GUID from Standard;    
   
    ID(me)
    	returns GUID from Standard
	is redefined static;
	---Purpose: Returns the ID of the attribute.
	--          
	---C++: return const &

    PatternID(me)
    	returns GUID from Standard
	is deferred;
	---Purpose: Returns the ID of the attribute.
	--          
	---C++: return const &

    NbTrsfs(me)
    returns Integer from Standard
    is deferred;
        ---Purpose: Give the number of transformation

    ComputeTrsfs(me; Trsfs : in out Array1OfTrsf from TDataXtd)
    is deferred;
        ---Purpose: Give the transformations

end Pattern;


