-- Created on: 2000-06-07
-- Created by: Galina KULIKOVA
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class FixSmallBezierCurves from ShapeUpgrade inherits FixSmallCurves from ShapeUpgrade

	---Purpose: 

uses

    --HArray1OfCurve from TColGeom,
    --HArray1OfCurve from TColGeom2d,
    --HSequenceOfReal from TColStd,
    Edge from TopoDS,
    Face from TopoDS,
    Curve from Geom,
    Curve from Geom2d,
    Status from ShapeExtend
is

    Create returns FixSmallBezierCurves from ShapeUpgrade;
    ---Purpose :
    
    Approx(me : mutable; Curve3d :  out Curve from Geom;
    	   	    	 Curve2d :  out Curve from Geom2d;
    	    	    	 Curve2dR : out Curve from Geom2d;
    	    	    	 First, Last : in out Real) returns Boolean is redefined;
    --Perform(me : mutable; theSegments3d :in out HArray1OfCurve from TColGeom;
    --	    	    	 theKnots3d : in out HSequenceOfReal from TColStd;
    --	    	    	 theSegments2d :in out HArray1OfCurve from TColGeom2d;
    --	    	    	 theKnots2d : in out HSequenceOfReal from TColStd) returns Boolean is redefined;
    ---Purpose :
    


end FixSmallBezierCurves;
