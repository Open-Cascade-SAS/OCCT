-- Created on: 1993-05-28
-- Created by: Modelistation
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class FaceClassifier from BRepClass inherits FClassifier from BRepClass

	---Purpose: Provides Constructors with a Face.

uses
    FaceExplorer from BRepClass,
    Face         from TopoDS,
    Pnt2d        from gp,
    Pnt          from gp

is
    Create returns FaceClassifier from BRepClass;
	---Purpose: Empty constructor, undefined algorithm.
	
	
	
      
    Create(F : in out FaceExplorer from BRepClass; 
    	   P : Pnt2d from gp; Tol : Real)
    returns FaceClassifier from BRepClass;
	---Purpose: Creates an algorithm to classify the Point  P with
	--          Tolerance <T> on the face described by <F>.
	
    Create(F : Face from TopoDS; 
    	   P : Pnt2d from gp; Tol : Real)
    returns FaceClassifier from BRepClass;
	---Purpose: Creates an algorithm to classify the Point  P with
	--          Tolerance <T> on the face <F>.
	
    Perform(me : in out;
    	    F : Face from TopoDS; 
    	    P : Pnt2d from gp; Tol : Real)
	---Purpose: Classify  the Point  P  with  Tolerance <T> on the
	--          face described by <F>.
    is static;

    
    Create(F : Face from TopoDS; 
    	   P : Pnt from gp; Tol : Real)
    returns FaceClassifier from BRepClass;
	---Purpose: Creates an algorithm to classify the Point  P with
	--          Tolerance <T> on the face <F>.
	
    Perform(me : in out;
    	    F : Face from TopoDS; 
    	    P : Pnt from gp; Tol : Real)
	---Purpose: Classify  the Point  P  with  Tolerance <T> on the
	--          face described by <F>.
    is static;   


end FaceClassifier;
