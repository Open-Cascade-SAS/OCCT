-- Created on: 2002-12-10
-- Created by: data exchange team
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V2.0

class VolumeElementPurpose from StepElement
inherits SelectType from StepData

    ---Purpose: Representation of STEP SELECT type VolumeElementPurpose

uses
    SelectMember from StepData,
    EnumeratedVolumeElementPurpose from StepElement,
    HAsciiString from TCollection

is
    Create returns VolumeElementPurpose from StepElement;
	---Purpose: Empty constructor

    CaseNum (me; ent: Transient) returns Integer;
	---Purpose: Recognizes a kind of VolumeElementPurpose select type
	--          return 0 

    CaseMem (me; ent: SelectMember from StepData) returns Integer is redefined;
	---Purpose: Recognizes a items of select member VolumeElementPurposeMember
	--          1 -> EnumeratedVolumeElementPurpose
	--          2 -> ApplicationDefinedElementPurpose
	--          0 else


     NewMember(me) returns SelectMember from StepData is redefined;
	---Purpose: Returns a new select member the type VolumeElementPurposeMember

    SetEnumeratedVolumeElementPurpose(me: in out; aVal :EnumeratedVolumeElementPurpose from StepElement);
	---Purpose: Set Value for EnumeratedVolumeElementPurpose

    EnumeratedVolumeElementPurpose (me) returns EnumeratedVolumeElementPurpose from StepElement;
	---Purpose: Returns Value as EnumeratedVolumeElementPurpose (or Null if another type)

    SetApplicationDefinedElementPurpose(me: in out; aVal :HAsciiString from TCollection);
	---Purpose: Set Value for ApplicationDefinedElementPurpose

    ApplicationDefinedElementPurpose (me) returns HAsciiString from TCollection;
	---Purpose: Returns Value as ApplicationDefinedElementPurpose (or Null if another type)

end VolumeElementPurpose;
