-- Created by: Peter KURNEV
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement. 

 
class Section from BOPAlgo  
    inherits Builder from BOPAlgo
 
    ---Purpose: 
    -- The algorithm to build a Secton between the arguments. 
    -- The Section consists of vertices and edges. 
    -- The Section contains:
    -- 1. new vertices that are subjects of V/V, E/E, E/F, F/F interferences
    -- 2. vertices that are subjects of V/E, V/F interferences
    -- 3. new edges that are subjects of F/F interferences
    -- 4. edges that are Common Blocks

    -- The vertex is included in Section only when it is not shared 
    -- between the edges above

uses 
    ShapeEnum from TopAbs,
    Shape from TopoDS,   
    ListOfShape from TopTools, 
    BaseAllocator from BOPCol,  
    PaveFiller from BOPAlgo 

--raises

is
    Create  
        returns Section from BOPAlgo;  
    ---C++: alias "Standard_EXPORT virtual ~BOPAlgo_Section();"  
    ---Purpose:  Empty constructor    
 
    Create (theAllocator: BaseAllocator from BOPCol)
        returns Section from BOPAlgo; 
    ---Purpose:  Empty constructor    
    --
    --  protected methods 
    -- 
    CheckData(me:out) 
        is redefined protected; 
    ---Purpose:  
    
    PerformInternal1(me:out; 
        thePF:PaveFiller from BOPAlgo) 
        is redefined protected;   
    ---Purpose:  Performs calculations using prepared Filler 
    --           object <thePF>          	 
     
    BuildSection(me:out) 
        is virtual; 
    --
    --  History 
    -- 
    Generated (me:out;  
            theS : Shape from TopoDS) 
        returns ListOfShape from TopTools
        is redefined; 
    ---C++: return const & 
    ---Purpose: Returns the  list of shapes generated from the
    --          shape theS. 
    
end Section;
