-- Created on: 1996-12-05
-- Created by: Jacques MINOT/Odile Olivier/Serguei ZARITCHNY
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Modified     Mon 12-january-98
--		<odl@sacadox.paris1.matra-dtv.fr>, 


class DiameterDimension from AIS inherits Relation from AIS


	---Purpose: A framework to display diameter dimensions.
    	-- A diameter is displayed with arrows and text. The
    	-- text gives the length of the diameter.
    	-- The algorithm takes a length along a face and
    	-- analyzes it as an arc. It then reconstructs the circle
    	-- corresponding to the arc and calculates the
    	-- diameter of this circle. This diameter serves as a
    	-- relational reference in 3d presentations of the surface.
	
uses

     Shape                 from TopoDS,
     Circ                  from gp,
     Pnt                   from gp, 
     Pln                   from gp, 
     Plane                 from Geom, 
     Surface               from Geom,
     Presentation          from Prs3d,
     PresentationManager3d from PrsMgr,
     Selection             from SelectMgr,
     Projector             from Prs3d,
     Transformation        from Geom,
     ExtendedString        from TCollection,    
     ArrowSide             from DsgPrs, 
     KindOfSurface         from AIS,
     KindOfDimension       from AIS 

raises ConstructionError from Standard     
      
is
    Create (aShape      : Shape          from TopoDS;
	    aVal        : Real           from Standard;
	    aText       : ExtendedString from TCollection)    
	---Purpose: Constructs a diameter display object defined by the
    	-- shape aFShape, the dimension aVal and the text aText.
    returns mutable DiameterDimension from AIS;

    Create (aShape      : Shape          from TopoDS;
	    aVal        : Real           from Standard;
	    aText       : ExtendedString from TCollection;	    
	    aPosition   : Pnt            from gp;
	    aSymbolPrs  : ArrowSide      from DsgPrs;    
	    aDiamSymbol : Boolean        from Standard;    
    	    anArrowSize : Real           from Standard = 0.0)
	---Purpose: Constructs a diameter display object defined by the
    	-- shape aFShape, the dimension aVal and the text
    	-- aText, the point of origin of the diameter aPosition,
    	-- and the type of arrow aSymbolPrs with the size anArrowSize.
    	-- If the Boolean aDiamSymbol is true.
    returns mutable DiameterDimension from AIS;

    KindOfDimension(me) returns KindOfDimension from AIS 
        ---C++: inline
    	---Purpose:
    	-- Indicates that we are concerned with a length.
    is redefined;

    IsMovable(me) returns Boolean from Standard 
        ---C++: inline    
    	---Purpose:
    	-- Returns true if the diameter dimension is movable
    is redefined;        

    DiamSymbol(me: mutable) returns Boolean from Standard 
	---C++: inline
	---Purpose:
    	-- Returns the symbol for diameter dimension. This will
    	-- be either arrow, text, or a combination of both.
    is static;

    SetDiamSymbol(me: mutable;aDiamSymbol: Boolean from Standard) 
        ---C++: inline
    	---Purpose:
    	-- Sets the symbol for diameter dimension aDiamSymbol.
    	-- This can be an arrow, a text or both.
    is static;
 
--    SetPlane(me: mutable; aPlane : Plane from Geom)
--    is static;
--    ---C++: inline
    
--    Plane(me) returns any Plane  from Geom 
--    is static;
--    ---C++: inline
--    ---C++: return  const  & 

          
-- Methods from PresentableObject

    Compute(me                  : mutable;
    	    aPresentationManager: PresentationManager3d from PrsMgr;
    	    aPresentation       : mutable Presentation from Prs3d;
    	    aMode               : Integer from Standard= 0) 
    is redefined private;
    
    Compute(me:mutable;
    	        aProjector: Projector from Prs3d;
                aPresentation: mutable Presentation from Prs3d)
    is redefined static private;     
    
    Compute(me            : mutable;
    	    aProjector    : Projector from Prs3d;
    	    aTrsf         : Transformation from Geom;
	    aPresentation : mutable Presentation from Prs3d)
    is redefined;
    ---Purpose: computes the presentation according to a point of view
    --          given by <aProjector>. 
    --          To be Used when the associated degenerated Presentations 
    --          have been transformed by <aTrsf> which is not a Pure
    --          Translation. The HLR Prs can't be deducted automatically
    --          WARNING :<aTrsf> must be applied
    --           to the object to display before computation  !!!

-- Methods from SelectableObject

    ComputeSelection(me         : mutable;
    	    	     aSelection : mutable Selection from SelectMgr;
    	    	     aMode      : Integer from Standard)
    is redefined private;

--
--     Computation private methods
--

    ComputeOneFaceDiameter(me: mutable;
    	    	     	aPresentation : mutable Presentation from Prs3d)
    is private; 
     
    ComputeOneCylFaceDiameter(me: mutable;
    	    	     	aPresentation : mutable Presentation from Prs3d; 
    	    	     	aSurfType     : KindOfSurface  from  AIS; 
    	    	    	aSurf         : Surface  from  Geom  )
    is private; 
     
    ComputeOnePlanarFaceDiameter(me: mutable;
    	    	     	aPresentation : mutable Presentation from Prs3d  )
    is private; 
    
    ComputeOneEdgeDiameter(me: mutable;
    	    	     	aPresentation : mutable Presentation from Prs3d)
    is private;
    
    ComputeCircleDiameter(me: mutable;
    	    	     	  aPresentation : mutable Presentation from Prs3d)
    is private;
    
    ComputeArcDiameter(me: mutable;
    	    	       aPresentation : mutable Presentation from Prs3d; 
    	    	       ptFirst : Pnt from gp;
    	    	       ptend   : Pnt from gp)
    is private;
    
    ComputeArcSelection(me      : mutable;
    	    	     aSelection : mutable Selection from SelectMgr)
    is private;
    
fields
     
    myCircle       : Circ    from gp;
    myIsAnArc      : Boolean from Standard;
    myDiamSymbol   : Boolean from Standard; 
    myFirstPar     : Real    from Standard;      
    myLastPar      : Real    from Standard;   

end DiameterDimension;
