-- Created on: 1995-03-31
-- Created by: Jean-Louis Krenkel
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Update:      Thu Mar 24 16:05:00 1998
--              Adds <useMFT> parameter in the SetFontMap() method
--              and adds the new method UseMFT()
--              for using MDTV fonts instead system fonts.


class Viewer from V2d inherits Viewer from Viewer
---Purpose:
-- This class defines a 2D viewer which manages one
-- 2D view at least and the attributes of this view (ex: ColorMap, etc.).
uses
    ColorMap,TypeMap,WidthMap,FontMap,MarkMap from Aspect,
    GraphicDevice from Aspect,
    ExtendedString,AsciiString from TCollection,
    View from V2d,
    View from Graphic2d,
    RectangularGrid from V2d,CircularGrid from V2d,
    Grid from Aspect,
    GridType from Aspect,GridDrawMode from Aspect,
    NameOfColor from Quantity,Length from Quantity,
    Color from Quantity,
    PlaneAngle from Quantity,
    ListOfTransient from TColStd,
    ListIteratorOfListOfTransient from TColStd
is

    Create(aGraphicDevice: GraphicDevice from Aspect;
	   aName: ExtString from Standard;
	   aDomain: CString from Standard = "")
    returns mutable Viewer from V2d;
---Purpose:
-- Constructs a viewer object defined by the graphic
-- device aGraphicDevice that determines the screen
-- attributes, a default view and the name aName.
        
    Create(aGraphicDevice: GraphicDevice from Aspect;
    	   aView: View from Graphic2d;
	   aName: ExtString from Standard;
	   aDomain: CString from Standard = "")
    returns mutable Viewer from V2d;
---Purpose:
-- Constructs a viewer object defined by the graphic
-- device aGraphicDevice that determines the screen
-- attributes, the first view aView and the name aName.
        
    AddView(me: mutable; aView: View from V2d)
    is static;
---Purpose: Adds another 2D view to the viewer.    
    RemoveView(me: mutable; aView: View from V2d)
    is static;
---Purpose: Removes the view aView from the viewer.
    Update(me: mutable)
    is redefined static;
---Purpose: Updates the display of all views of the viewer.
    UpdateNew(me: mutable)
    is static;
---Purpose: Updates the most recent changes in all the active views of the viewer.
    SetColorMap(me: mutable; aColorMap: ColorMap from Aspect) 
    is static;
---Purpose:
-- Replaces the default color map of the viewer with the
-- new color map aColorMap.    
    SetTypeMap(me: mutable; aTypeMap: TypeMap from Aspect) 
    is static;
---Purpose:
-- Replaces the default type map of the viewer with the
-- new type map aTypeMap.    
    SetWidthMap(me: mutable; aWidthMap: WidthMap from Aspect) 
    is static;
---Purpose:
-- Replaces the default width map of the viewer with the
-- new width map aWidthMap.    
    SetFontMap(me: mutable; aFontMap: FontMap from Aspect;
			    useMFT: Boolean from Standard = Standard_True) 
    is static;
---Purpose:
-- Replaces the default font map of the viewer with the
-- new font map aFontMap. When useMFT is equal to
-- Standard_True, MDTV fonts are used instead of system fonts.
    SetMarkMap(me: mutable; aMarkMap: MarkMap from Aspect) 
    is static;
---Purpose:
-- Replaces the default mark map of the viewer with the
-- new mark map aMarkMap.    
    ColorMap(me) returns ColorMap from Aspect
    is static;
 --- Purpose: Returns the active color map of the viewer.  
    TypeMap(me) returns  TypeMap from Aspect 
    is static;
--- Purpose: Returns the active type map of the viewer.   
    WidthMap(me) returns WidthMap from Aspect
    is static;
---Purpose: Returns the active width map of the viewer.    
    FontMap(me) returns  FontMap from Aspect 
    is static;
---Purpose: Returns the active font map for the viewer.
    MarkMap(me) returns MarkMap from Aspect
    is static;
---Purpose: Returns the active mark map of the viewer.
    UseMFT ( me ) returns Boolean from Standard 
    is static;
---Purpose: Returns True when the viewer uses MFT fonts
-- instead of system fonts.    
    View(me) returns View from Graphic2d;
  ---Purpose: Returns the first view of the viewer.  
    InitializeColor(me: mutable; aColor: NameOfColor from Quantity)
    ---Purpose: Creates a color in the color map of the driver if 
    --          the color does not yes exist.
    --          Returns the index of the color in the modified color map.
    returns Integer from Standard;

    InitActiveViews(me: mutable) 
    ---Purpose: initializes an iteration on the active views.
    is static;
	
    MoreActiveViews (me)
    returns Boolean from Standard
    ---Purpose: returns true if there are more active view(s) to return.
    is static;
	
    NextActiveViews (me: mutable)
    ---Purpose : Go to the next active view
    --           (if there is not, ActiveView will raise an exception)
    is static;
	
    ActiveView(me)
    returns mutable View from V2d is static;

 ---Purpose:
-- Returns the current view from the activated views.
    
    IsEmpty(me) returns Boolean from Standard;

---Purpose:
-- Returns True when no more secondary views exist in the viewer.
    Grid(me) returns mutable Grid from Aspect
    is static private;
    
    GridType(me) returns GridType from Aspect
    ---Purpose: returns the current grid type.
    is static;
    
    Hit(me; X,Y: Length from Quantity;
    	    gx,gy: out Length from Quantity)
    ---Purpose: returns the point (gx,gy) according to the grid.
    is static;

    ActivateGrid(me: mutable; aGridType: GridType from Aspect;
    	                      aGridDrawMode: GridDrawMode from Aspect)
    is static;

    DeactivateGrid(me: mutable)
    is static;

    IsActive(me) 
    returns Boolean from Standard
    is static;
---Purpose: Returns True when a grid is active in the viewer.    
    RectangularGridValues(me; 
          XOrigin, YOrigin, XStep, YStep: out Length from Quantity;
    	  RotationAngle: out PlaneAngle from Quantity)
    is static;
---Purpose: Returns the parameters of the current rectangular grid.
    SetRectangularGridValues(me: mutable; 
          XOrigin, YOrigin, XStep, YStep: Length from Quantity;
    	  RotationAngle: PlaneAngle from Quantity)
    is static;
 ---Purpose:
-- Sets the rectangular grid:
-- -   XOrigin, YOrigin define the point of origin of the grid,
-- -   XStep defines the interval between two vertical lines,
-- -   YStep defines the interval between two horizontal lines,
-- -   RotationAngle defines the rotation angle of the grid. 
    
    CircularGridValues(me; 
          XOrigin, YOrigin, RadiusStep: out Length from Quantity;
	  DivisionNumber: out Integer from Standard;
    	  RotationAngle: out PlaneAngle from Quantity)
    is static;
---Purpose: Returns the parameters of the current circular grid.
    SetCircularGridValues(me: mutable; 
          XOrigin, YOrigin, RadiusStep: Length from Quantity;
	  DivisionNumber: Integer from Standard;
    	  RotationAngle: PlaneAngle from Quantity)
    is static;
---Purpose:
-- Sets the circular grid:
-- -   XOrigin, YOrigin specify the origin of the grid,
-- -   RadiusStep defines the interval between two circles,
-- -   DivisionNumber determines the section number of half a circle,
-- -   RotationAngle defines the rotation angle of the grid.    

    SetGridColor(me: mutable; color1, color2 : Color from Quantity)
    is static;
    
    HitPointMarkerIndex(me) returns Integer from Standard
    is static private;
    
    HitPointColor(me) returns Integer from Standard
    is static private;
    
    CoordinatesColor(me) returns Integer from Standard
    is static private;
    
    Init(me:mutable) 
    is static private;
    
    
    
fields

    myColorMap: ColorMap from Aspect;
    myTypeMap: TypeMap from Aspect;
    myWidthMap: WidthMap from Aspect;
    myFontMap: FontMap from Aspect;
    myMarkMap: MarkMap from Aspect;
    myGraphicView: View from Graphic2d;
    myViews: ListOfTransient from TColStd;
    myViewsIterator:ListIteratorOfListOfTransient from TColStd;

    myRGrid: RectangularGrid from V2d;
    myCGrid: CircularGrid from V2d;
    myHitPointMarkerIndex: Integer from Standard;
    myHitPointColorIndex: Integer from Standard;
    myCoordinatesColorIndex: Integer from Standard;
    myGridType: GridType from Aspect;    
    myUseMFT: Boolean from Standard;
friends
    class View from V2d
end Viewer from V2d;
