-- Created on: 1997-04-01
-- Created by: Christian CAILLET
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class FieldList1  from StepData    inherits FieldList  from StepData

    ---Purpose : Describes a list of ONE field

uses Field from StepData

raises OutOfRange

is

    Create returns FieldList1;
    ---Purpose : Creates a FieldList of 1 Field

    NbFields (me) returns Integer  is redefined;
    ---Purpose : Returns the count of fields. Here, returns 1

    Field  (me; num : Integer) returns Field
    ---Purpose : Returns the field n0 <num> between 1 and NbFields (read only)
	raises OutOfRange
    --           Error if <num> out of range
    	is redefined;
    ---C++ : return const &

    CField (me : in out; num : Integer) returns Field
    ---Purpose : Returns the field n0 <num> between 1 and NbFields, in order to
    --           modify its content
	raises OutOfRange
    --           Error if <num> out of range
    	is redefined;
    ---C++ : return &

    Destroy (me: in out) is virtual;
    ---C++ : alias "Standard_EXPORT virtual ~StepData_FieldList1() { Destroy(); }"

fields

    thefield : Field from StepData;

end FieldList1;
