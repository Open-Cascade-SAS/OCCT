-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class AutoDesignOrganizationAssignment from StepAP214 

inherits OrganizationAssignment from StepBasic 

uses

	HArray1OfAutoDesignGeneralOrgItem from StepAP214, 
	AutoDesignGeneralOrgItem from StepAP214, 
	Organization from StepBasic, 
	OrganizationRole from StepBasic
is

	Create returns AutoDesignOrganizationAssignment;
	---Purpose: Returns a AutoDesignOrganizationAssignment


	Init (me : mutable;
	      aAssignedOrganization : Organization from StepBasic;
	      aRole : OrganizationRole from StepBasic) is redefined;

	Init (me : mutable;
	      aAssignedOrganization : Organization from StepBasic;
	      aRole : OrganizationRole from StepBasic;
	      aItems : HArray1OfAutoDesignGeneralOrgItem from StepAP214) is virtual;

	-- Specific Methods for Field Data Access --

	SetItems(me : mutable; aItems : HArray1OfAutoDesignGeneralOrgItem);
	Items (me) returns HArray1OfAutoDesignGeneralOrgItem;
	ItemsValue (me; num : Integer) returns AutoDesignGeneralOrgItem;
	NbItems (me) returns Integer;

fields

	items : HArray1OfAutoDesignGeneralOrgItem from StepAP214; -- a SelectType

end AutoDesignOrganizationAssignment;
