-- Created on: 1992-11-18
-- Created by: Christian CAILLET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



deferred class SelectAnyType  from IFSelect  inherits SelectExtract

    ---Purpose : A SelectAnyType sorts the Entities of which the Type is Kind
    --           of a given Type : this Type for Match is specific of each
    --           class of SelectAnyType

uses Type, InterfaceModel

is

    TypeForMatch (me) returns Type  is deferred;
    ---Purpose : Returns the Type which has to be matched for select

    Sort (me; rank : Integer; ent : Transient; model : InterfaceModel)
    	returns Boolean;
    ---Purpose : Returns True for an Entity (model->Value(num)) which is kind
    --           of the choosen type, given by the method TypeForMatch.
    --           Criterium is IsKind.

end SelectAnyType;
