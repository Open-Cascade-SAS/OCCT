-- Created on: 1994-06-17
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class FacetedBrepAndBrepWithVoids from StepShape 

inherits ManifoldSolidBrep from StepShape 


	--- This class is an implementation of EXPRESS
	--  ANDOR Subtype Declaration.
uses

	FacetedBrep from StepShape, 
	BrepWithVoids from StepShape, 
	ClosedShell from StepShape, 
	HArray1OfOrientedClosedShell from StepShape, 
	OrientedClosedShell from StepShape,
	HAsciiString from TCollection
is

	Create returns mutable FacetedBrepAndBrepWithVoids;
	---Purpose: Returns a FacetedBrepAndBrepWithVoids


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aOuter : mutable ClosedShell from StepShape) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aOuter : mutable ClosedShell from StepShape;
	      aFacetedBrep : mutable FacetedBrep from StepShape;
	      aBrepWithVoids : mutable BrepWithVoids from StepShape);

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aOuter : mutable ClosedShell from StepShape;
	      aVoids : mutable HArray1OfOrientedClosedShell from StepShape);

	-- Specific Methods for Field Data Access --

	SetFacetedBrep(me : mutable; aFacetedBrep : mutable FacetedBrep);
	FacetedBrep (me) returns mutable FacetedBrep;
	SetBrepWithVoids(me : mutable; aBrepWithVoids : mutable BrepWithVoids);
	BrepWithVoids (me) returns mutable BrepWithVoids;

	-- Specific Methods for ANDOR Field Data Access --

	SetVoids(me : mutable; aVoids : mutable HArray1OfOrientedClosedShell);
	Voids (me) returns mutable HArray1OfOrientedClosedShell;
	VoidsValue (me; num : Integer) returns mutable OrientedClosedShell;
	NbVoids (me) returns Integer;

	-- Specific Methods for ANDOR Field Data Access --


fields

	facetedBrep : FacetedBrep from StepShape;
	brepWithVoids : BrepWithVoids from StepShape;

end FacetedBrepAndBrepWithVoids;
