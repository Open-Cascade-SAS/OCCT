-- Created on: 1997-04-21
-- Created by: Denis PASCAL
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



deferred class Dimension from DrawDim inherits Drawable3D from Draw

	---Purpose: 

uses 
    Real       from Standard,
    Pnt        from gp,
    Color      from Draw,
    Display    from Draw

is

    Initialize;

    SetValue (me : mutable; avalue : Real from Standard);
    
    GetValue (me)
    returns Real from Standard;
    
    IsValued (me)
    returns Boolean from Standard;
    
    TextColor(me : mutable; C : Color from Draw);
    
    TextColor(me) returns Color from Draw;
    
    DrawText(me; Pos : Pnt from gp; D : in out Display from Draw);
    
fields

    is_valued     : Boolean from Standard is protected;
    myValue       : Real    from Standard is protected;
    myTextColor   : Color   from Draw     is protected;
    
end Dimension;
