-- Created on: 2001-07-25
-- Created by: Julia DOROVSKIKH
-- Copyright (c) 2001-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DocumentRetrievalDriver from XmlDrivers inherits DocumentRetrievalDriver from XmlLDrivers

uses

    ADriverTable		from XmlMDF, 
    ADriver                     from XmlMDF, 
    Element                     from XmlObjMgt,
    MessageDriver               from CDM

is
    Create returns mutable DocumentRetrievalDriver from XmlDrivers;
    -- Constructor

    AttributeDrivers	(me : mutable; theMsgDriver: MessageDriver from CDM)
	returns ADriverTable from XmlMDF
	is redefined virtual; 
	 
    ReadShapeSection (me:mutable; thePDoc  :  Element from XmlObjMgt; 
                                  theMsgDriver : MessageDriver from CDM) 
        returns ADriver from XmlMDF
        is redefined virtual; 
	 
    ShapeSetCleaning(me:mutable; theDriver : ADriver from XmlMDF) 
        is redefined virtual;
	
    PropagateDocumentVersion(me:mutable; theDocVersion : Integer from Standard) 
        is redefined virtual;  
	 
end DocumentRetrievalDriver;
