-- Created on: 1996-06-04
-- Created by: Stagiaire Xuan Trang PHAMPHU
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Corde from BlendFunc

	---Purpose: This function calculates point (pts) on the curve of
 	--          intersection between the normal to a curve (guide)
 	--          in a chosen parameter and a surface  (surf), so
 	--          that pts was at a given distance from the guide.
	--          X(1),X(2) are the parameters U,V of pts on surf.

 
uses Vector   from math,
     Matrix   from math,
     Gauss    from math,	
     Vec      from gp,
     Vec2d    from gp,	     	    
     Pnt      from gp,
     Pnt2d    from gp,
     HCurve   from Adaptor3d,
     HSurface from Adaptor3d

raises  
    DomainError from Standard
    	
     
is

    Create(S: HSurface from Adaptor3d; CGuide: HCurve from Adaptor3d)     
    	returns Corde from BlendFunc;
	
	
    SetParam(me: in out; Param: Real from Standard);


    SetDist(me: in out; Dist: Real from Standard);
       
		
    Value(me: in out; X: Vector; F: out Vector)
    	---Purpose: computes the values <F> of the Function for the 
    	--          variable <X>.
    	--          Returns True if the computation was done successfully, 
    	--          False otherwise.

    	returns Boolean from Standard;    	

	
    Derivatives(me: in out; X: Vector; D: out Matrix)
    	---Purpose: returns the values <D> of the derivatives for the 
    	--          variable <X>.
    	--          Returns True if the computation was done successfully, 
    	--          False otherwise.	

    returns Boolean from Standard;
    
 
    PointOnS(me)
    
    	returns Pnt from gp
	---C++: return const&
	;


    PointOnGuide(me)
    
    	returns Pnt from gp
	---Purpose: returns the point of parameter <Param> on CGuide
	---C++: return const&
	;
	
    NPlan(me)
    
    	returns Vec from gp
	---Purpose: returns the normal to CGuide at Ptgui.
	---C++: return const&           
	;
	
    IsTangencyPoint(me)
    
	---Purpose: Returns True when it is not possible to compute
	--          the tangent vectors at PointOnS.
    
    	returns Boolean from Standard;
	
	
    TangentOnS(me)
    
	---Purpose: Returns the tangent vector at PointOnS, in 3d space.

    	returns Vec from gp
	---C++: return const&
    	raises DomainError from Standard;
	--- The exception is raised when IsTangencyPoint
	--  returns Standard_True.	
	
	    
    Tangent2dOnS(me)
    
	---Purpose: Returns the tangent vector at PointOnS, in the
	--          parametric space of the first surface.

    	returns Vec2d from gp
	---C++: return const&
    	raises DomainError from Standard;
	--- The exception is raised when IsTangencyPoint
	--  returns Standard_True.	

	    
    DerFguide(me: in out; Sol : Vector from math; DerF : out Vec2d from gp);
	---Purpose: Derived of the function compared to the parameter
	-- of the guideline
			
			
    IsSolution(me : in out;
    	       Sol: Vector from math; Tol: Real from Standard)  
	  
	---Purpose: Returns False if Sol is not solution else returns
	--          True and updates the fields tgs and tg2d  
      
      returns Boolean from Standard;  
    
fields

    surf       : HSurface from Adaptor3d;    
    guide      : HCurve from Adaptor3d;	
    pts        : Pnt     from gp;
    pt2d       : Pnt2d   from gp;
    dis        : Real    from Standard;
    normtg     : Real    from Standard;	
    theD       : Real    from Standard;     
    ptgui      : Pnt     from gp;
    nplan      : Vec     from gp;	
    d1gui      : Vec     from gp;
    d2gui      : Vec     from gp;
    tgs        : Vec     from gp;
    tg2d       : Vec2d   from gp; 
    istangent  : Boolean from Standard;	

end Corde;    
