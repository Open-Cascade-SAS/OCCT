-- File:	TopOpeBRepBuild_SolidAreaBuilder.cdl
-- Created:	Thu Dec 21 17:07:40 1995
-- Author:	Jean Yves LEBEY
--		<jyl@meteox>
---Copyright:	 Matra Datavision 1995

class SolidAreaBuilder from TopOpeBRepBuild 
    inherits Area3dBuilder from TopOpeBRepBuild

---Purpose: 
-- The SolidAreaBuilder algorithm is used to construct Solids from a LoopSet,
-- where the Loop is the composite topological object of the boundary,
-- here wire or block of edges.
-- The LoopSet gives an iteration on Loops.
-- For each Loop  it indicates if it is on the boundary (wire) or if it
-- results from  an interference (block of edges).
-- The result of the SolidAreaBuilder is an iteration on areas.
-- An area is described by a set of Loops.

uses

    LoopSet from TopOpeBRepBuild,
    LoopClassifier from TopOpeBRepBuild
    
is

    Create returns SolidAreaBuilder;

    Create(LS : in out LoopSet; LC : in out LoopClassifier;
    	   ForceClass : Boolean = Standard_False) returns SolidAreaBuilder;
    ---Purpose: Creates a SolidAreaBuilder to build Solids on
    -- the (shells,blocks of face) of <LS>, using the classifier <LC>.
    
    InitSolidAreaBuilder(me: in out;
    	    	         LS : in out LoopSet; LC : in out LoopClassifier;
    	    	         ForceClass : Boolean = Standard_False) is static;
		    
end SolidAreaBuilder from TopOpeBRepBuild;
