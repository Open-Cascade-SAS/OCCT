-- Created on: 1995-12-08
-- Created by: Jean-Pierre COMBE
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class SymbPresentation from DsgPrs
    	---Purpose: A framework to define display of symbols.
uses
    Presentation from Prs3d,
    Pnt from gp,
    Drawer from Prs3d,
    ExtendedString from TCollection
    	
is  
    Add( myclass; aPresentation: Presentation from Prs3d;
    	    	  aDrawer: Drawer from Prs3d;
		  aText: ExtendedString from TCollection;
		  OffsetPoint: Pnt from gp);
    	---Purpose: Adds the text aText and the point OffsetPoint to the
    	-- presentation object aPresentation.
    	-- The display attributes of the shaded plane are
    	-- defined by the attribute manager aDrawer.

end SymbPresentation;
