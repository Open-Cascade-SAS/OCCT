-- Created on: 1994-06-01
-- Created by: Christian CAILLET
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class SelectFromDrawing  from IGESSelect  inherits SelectDeduct

    ---Purpose : This selection gets in all the model, the entities which are
    --           attached to the drawing(s) given as input. This includes :
    --           - Drawing Frame (Annotations directky referenced by Drawings)
    --           - Entities attached to the single Views referenced by Drawings

uses AsciiString from TCollection, EntityIterator, Graph

raises InterfaceError

is

    Create returns mutable SelectFromDrawing;
    ---Purpose : Creates a SelectFromDrawing

    RootResult (me; G : Graph) returns EntityIterator  raises InterfaceError;
    ---Purpose : Selects the Entities which are attached to the Drawing(s)
    --           present in the Input

    Label (me) returns AsciiString from TCollection;
    ---Purpose : Returns the label, with is "Entities attached to Drawing"

end SelectFromDrawing;
