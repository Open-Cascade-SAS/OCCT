-- File:        RepresentationMap.cdl
-- Created:     Mon Dec  4 12:02:31 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWRepresentationMap from RWStepRepr

	---Purpose : Read & Write Module for RepresentationMap

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     RepresentationMap from StepRepr,
     EntityIterator from Interface

is

	Create returns RWRepresentationMap;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable RepresentationMap from StepRepr);

	WriteStep (me; SW : in out StepWriter; ent : RepresentationMap from StepRepr);

	Share(me; ent : RepresentationMap from StepRepr; iter : in out EntityIterator);

end RWRepresentationMap;
