-- Created by: DAUTRY Philippe
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

--      	----------------

---Version:	0.0
--Version	Date		Purpose
--		0.0	Apr  4 1997	Creation


deferred class ASDriver from MDF
    inherits TShared from MMgt

	---Purpose: Attribute Storage Driver.

uses

    Attribute from TDF,
    Attribute from PDF,
    SRelocationTable from MDF, 
    MessageDriver from CDM, 
    ExtendedString from TCollection

-- raises

is
    Initialize (theMessageDriver : MessageDriver from CDM); 
    
    VersionNumber(me) returns Integer from Standard
    	is deferred;
	---Purpose: Returns the version number from which the driver
	--          is available.

    SourceType(me) returns Type from Standard
    	is deferred;
	---Purpose: Returns the type of source object, inheriting from
	--          Attribute from TDF.

    NewEmpty(me)
    	returns mutable Attribute from PDF
    	is deferred;
	---Purpose: Creates a new attribute from PDF.

    Paste(me;
    	  aSource     :         Attribute from TDF;
    	  aTarget     : mutable Attribute from PDF;
    	  aRelocTable : SRelocationTable from MDF)
    	is deferred;
	---Purpose: Translate the contents of <aSource> and put it
	--          into <aTarget>, using the relocation table
	--          <aRelocTable> to keep the sharings. 
	
    WriteMessage (me; theMessage : ExtendedString from TCollection);
        ---Purpose: To send message to Application (if MessageDriver defined) 
	
fields 

    myMessageDriver : MessageDriver from CDM;  
    
end ASDriver;
