-- File:        ExtrudedAreaSolid.cdl
-- Created:     Fri Dec  1 11:11:20 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class ExtrudedAreaSolid from StepShape 

inherits SweptAreaSolid from StepShape 

uses

	Direction from StepGeom, 
	Real from Standard, 
	HAsciiString from TCollection, 
	CurveBoundedSurface from StepGeom
is

	Create returns mutable ExtrudedAreaSolid;
	---Purpose: Returns a ExtrudedAreaSolid


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aSweptArea : mutable CurveBoundedSurface from StepGeom) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aSweptArea : mutable CurveBoundedSurface from StepGeom;
	      aExtrudedDirection : mutable Direction from StepGeom;
	      aDepth : Real from Standard) is virtual;

	-- Specific Methods for Field Data Access --

	SetExtrudedDirection(me : mutable; aExtrudedDirection : mutable Direction);
	ExtrudedDirection (me) returns mutable Direction;
	SetDepth(me : mutable; aDepth : Real);
	Depth (me) returns Real;

fields

	extrudedDirection : Direction from StepGeom;
	depth : Real from Standard;

end ExtrudedAreaSolid;
