-- Created on: 1992-04-23
-- Created by: Modelistation
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Marker3D from Draw inherits Drawable3D from Draw

	---Purpose: 

uses
    Pnt from gp,
    Color from Draw,
    MarkerShape from Draw,
    Display from Draw

is
    Create(P : Pnt from gp; T : MarkerShape from Draw; C : Color from Draw; 
    	ISize : Integer = 5) returns mutable Marker3D from Draw;
	
    Create(P : Pnt from gp; T : MarkerShape from Draw; C : Color from Draw; 
    	RSize : Real) returns mutable Marker3D from Draw;

    ChangePos(me : mutable) returns Pnt from gp;
    ---C++: return &
    ---Purpose: myPos field

    DrawOn(me; dis : in out Display from Draw);

    PickReject(me; X,Y,Prec : Real) returns Boolean
    ---Purpose: Returs always false
    is redefined;

fields

    myPos : Pnt from gp;
    myCol : Color from Draw;
    myTyp : MarkerShape from Draw;
    mySiz : Integer;
    myRSiz : Real; 
    myIsRSiz : Boolean;

end Marker3D;
