-- Created on: 1994-06-27
-- Created by: Design
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class VoidBinder  from Transfer  inherits Binder

    ---Purpose : a VoidBinder is used to bind a starting item with a status,
    --           error or warning messages, but no result
    --           It is interpreted by TransferProcess, which admits a
    --           VoidBinder to be over-written, and copies its check to the
    --           new Binder

uses CString, Type

is

    Create returns mutable VoidBinder;

--    IsMultiple (me) returns Boolean;
    ---Purpose : a VoidBinder is not Multiple (Remark : it is not Simple too)
    --           But it can bring next results ...

    ResultType (me) returns Type;
    ---Purpose : while a VoidBinder admits no Result, its ResultType returns
    --           the type of <me>

    ResultTypeName (me) returns CString;
    ---Purpose : Returns "(void)"

end VoidBinder;
