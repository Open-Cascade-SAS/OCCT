-- File:	StepVisual_MarkerMember.cdl
-- Created:	Tue Apr  1 18:01:43 1997
-- Author:	Christian CAILLET
--		<cky@heliox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1997


class MarkerMember  from StepVisual    inherits SelectInt  from StepData

    ---Purpose : Defines MarkerType as unique member of MarkerSelect
    --           Works with an EnumTool

uses CString, MarkerType from StepVisual

is

    Create returns mutable MarkerMember;

    HasName (me) returns Boolean  is redefined;
    -- returns True

    Name    (me) returns CString  is redefined;
    -- returns MARKER_TYPE

    SetName (me : mutable; name : CString)  returns Boolean  is redefined;
    -- does nothing and returns True

    EnumText (me) returns CString  is redefined;
    -- returns the string counterpart of a value

    SetEnumText (me : mutable; val : Integer; text : CString)  is redefined;
    -- considers text and interprets it to set val

    SetValue  (me : mutable; val : MarkerType from StepVisual);
    -- Sets directly the good value as enum

    Value     (me) returns MarkerType from StepVisual;

end MarkerMember;
