-- Created on: 1994-03-28
-- Created by: Remi LEQUETTE
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Point from DrawTrSurf inherits Drawable3D from Draw

	---Purpose: A drawable point.

uses
    	Pnt from gp,
    	Pnt2d from gp,
	MarkerShape from Draw,
     	Color from Draw,
     	Display from Draw,
     	Drawable3D from Draw,
	Interpretor from Draw

is

    Create( P : Pnt from gp; 
    	    Shape : MarkerShape from Draw;
	    Col   : Color from Draw) 
    returns mutable Point from DrawTrSurf;
    
    Create( P : Pnt2d from gp; 
    	    Shape : MarkerShape from Draw;
	    Col   : Color from Draw) 
    returns mutable Point from DrawTrSurf;
    
    DrawOn (me; dis : in out Display from Draw);
     
    Is3D(me) returns Boolean
	---Purpose: Is a 3D object. (Default True).
    is redefined;
    
    Point(me) returns Pnt from gp
    is static;
    
    Point(me : mutable; P : Pnt from gp)
    is static;

    Point2d(me) returns Pnt2d from gp
    is static;
    
    Point2d(me : mutable; P : Pnt2d from gp)
    is static;

  Color(me : mutable; aColor : Color from Draw)
     is static;

  Color (me)  returns Color from Draw
     is static;
     
  Shape(me : mutable; S : MarkerShape from Draw)
  is static;
  
  Shape(me) returns MarkerShape from Draw
  is  static;
     
  Copy(me) returns mutable Drawable3D from Draw
	---Purpose: For variable copy.
  is redefined;
  
  Dump(me; S : in out OStream)
	---Purpose: For variable dump.
  is redefined;

  Whatis(me; I : in out Interpretor from Draw)
	---Purpose: For variable whatis command.
  is redefined;

fields

    myPoint : Pnt from gp;
    is3D    : Boolean;
    myShape : MarkerShape from Draw;
    myColor : Color from Draw;

end Point;


