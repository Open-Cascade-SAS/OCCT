-- Created on: 1995-03-06
-- Created by: Laurent PAINNOT
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




package Poly

        ---Purpose: This  package  provides  classes  and services  to
        --          handle :
        --
        --          * 3D triangular polyhedrons.
        --
        --          * 3D polygons.
        --
        --          * 2D polygon.
        --
        --          * Tools to dump, save and restore those objects.

uses

    MMgt,
    TCollection,
    TColStd,
    gp,
    TColgp,
    TShort

is

    class Triangle;
        ---Purpose: A triangle is  a triplet  of integers (indices  of
        --          the nodes).

    class Array1OfTriangle
    instantiates Array1 from TCollection(Triangle from Poly);

    class HArray1OfTriangle
    instantiates HArray1 from TCollection(Triangle         from Poly,
                                          Array1OfTriangle from Poly);

    class Triangulation;
        ---Purpose: A   Triangulation  is  a   3D  polyhedron made  of
        --          triangles.  It   is  made  of  a nodes  which  are
        --          indexed. Nodes  have a 3d  value  and a  2d value.
        --          Triangles are triplet of node indices.
        --
        --          This is a Transient class.


    class Polygon3D;
        ---Purpose: A Polygon3D is  made of  indexed nodes.
        --          Nodes have a 3d value.

    class Polygon2D;
        ---Purpose: A Polygon2D is made of  indexed nodes.
        --          Nodes have a 2d value.

    class PolygonOnTriangulation;
        ---Purpose: A polygonOnTriangulation is made of node indices
        --          referencing a triangulation.


    --
    -- Tools to use triangulations
    --

    class Connect;
        ---Purpose: Computes and  stores  the    link from   nodes  to
        --          triangles     and from triangles to   neighbouring
        --          triangles.
        -- This tool is obsolete, replaced by Poly_CoherentTriangulation

    --
    --     Data types for the Coherent Triangulation data model
    --
    imported CogerentTriangulation;
    imported CoherentTriangle;
    imported CoherentNode;
    imported CoherentLink;
    imported CoherentTriPtr;
    imported ListOfTriangulation;

    imported MakeLoops;
        ---Purpose: Algorithm to make minimal loops in a graph

    --
    --  Package methods
    --

    Catenate (lstTri: ListOfTriangulation from Poly)
        returns Triangulation from Poly;
        ---Purpose: Join several triangulations to one new triangulation object.
        --          The new triangulation is just a mechanical sum of input
        --          triangulations, without node sharing. UV coordinates are
        --          dropped in the result.

    Write(T       : Triangulation from Poly;
          OS      : in out OStream;
          Compact : Boolean = Standard_True);

        ---Purpose: Writes the content of the triangulation <T> on the
        --          stream <OS>. If <Compact> is true this is a "save"
        --          format  intended  to  be read back   with the Read
        --          method. If compact is False  it is a "Dump" format
        --          intended to be informative.

    Write(P       : Polygon3D from Poly;
          OS      : in out OStream;
          Compact : Boolean = Standard_True);

        ---Purpose: Writes  the  content  of the 3D polygon <P> on the
        --          stream <OS>. If <Compact> is true this is a "save"
        --          format  intended  to  be read back   with the Read
        --          method. If compact is False  it is a "Dump" format
        --          intended to be informative.

    Write(P       : Polygon2D from Poly;
          OS      : in out OStream;
          Compact : Boolean = Standard_True);

        ---Purpose: Writes the  content  of the 2D polygon  <P> on the
        --          stream <OS>. If <Compact> is true this is a "save"
        --          format  intended  to  be read back   with the Read
        --          method. If compact is False  it is a "Dump" format
        --          intended to be informative.


    Dump(T       : Triangulation from Poly;
         OS      : in out OStream);
       ---Purpose: Dumps  the triangulation.  This   is a call to  the
       --          previous method with Comapct set to False.

    Dump(P       : Polygon3D from Poly;
         OS      : in out OStream);
       ---Purpose: Dumps  the  3D  polygon.  This   is a call to  the
       --          previous method with Comapct set to False.

    Dump(P       : Polygon2D from Poly;
         OS      : in out OStream);
       ---Purpose: Dumps  the  2D  polygon.  This   is a call to  the
       --          previous method with Comapct set to False.


    ReadTriangulation(IS : in out IStream)
    returns Triangulation from Poly;
        ---Purpose: Reads a triangulation from the stream <IS>.

    ReadPolygon3D(IS : in out IStream)
    returns Polygon3D from Poly;
        ---Purpose: Reads a 3d polygon from the stream <IS>.

    ReadPolygon2D(IS : in out IStream)
    returns Polygon2D from Poly;
        ---Purpose: Reads a 2D polygon from the stream <IS>.

    ComputeNormals(Tri : Triangulation from Poly);
        ---Purpose: Compute node normals for face triangulation
        --  as mean normal of surrounding triangles

    PointOnTriangle(P1, P2, P3, P: XY from gp; UV: out XY from gp)
    returns Real;
        ---Purpose: Computes parameters of the point P on triangle
        --          defined by points P1, P2, and P3, in 2d.
        --          The parameters U and V are defined so that
        --          P = P1 + U * (P2 - P1) + V * (P3 - P1),
        --          with U >= 0, V >= 0, U + V <= 1.
        --          If P is located outside of triangle, or triangle
        --          is degenerated, the returned parameters correspond
        --          to closest point, and returned value is square of
        --          the distance from original point to triangle (0 if
        --          point is inside).

end Poly;
