-- Created on: 1992-01-09
-- Created by: Remi GILET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


generic class FunctionTanObl from GccIter (
    TheCurve     as any;
    TheCurveTool as any) -- as CurvePGTool from GccInt (TheCurve)

inherits FunctionWithDerivative from math
    ---Purpose: This class describe a function of a single variable.

uses Dir2d from gp     

     
is

Create (Curve : TheCurve      ;
    	Dir   : Dir2d from gp ) returns FunctionTanObl from GccIter;

Value (me : in out      ;
       X  :        Real ;
       F  :    out Real ) returns Boolean;
    ---Purpose: Computes the value of the function F for the variable X.
    --          It returns True if the computation is successfully done,
    --          False otherwise.

Derivative (me    : in out      ;
            X     :        Real ;
            Deriv :    out Real ) returns Boolean;
    ---Purpose: Computes the derivative of the function F for the variable X.
    --          It returns True if the computation is successfully done,
    --          False otherwise.

Values (me    : in out      ;
        X     :        Real ;
        F     : out    Real ;
        Deriv : out    Real ) returns Boolean;
    ---Purpose: Computes the value and the derivative of the function F 
    --          for the variable X.
    --          It returns True if the computation is successfully done,
    --          False otherwise.

fields

TheCurv      : TheCurve        ;
TheDirection : Dir2d    from gp;

end FunctionTanObl;






