-- Created on: 1993-05-12
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred generic class ArcTool from Contap
    (TheArc as any )


    ---Purpose: Template class for a tool on the restriction of
    --          a surface.
    -- It is possible to implement this class with an instantiation
    -- of the class CurveTool from Adaptor3d.


uses Pnt2d from gp,
     Vec2d from gp

is

    Value(myclass; A: TheArc; X: Real from Standard)
    
	---Purpose: Returns the value in the parametric space
	--          of the surface S, of the point of parameter X
	--          on the arc A.

    	returns Pnt2d from gp;


    D1(myclass; A: TheArc; X: Real from Standard;
                P      : out Pnt2d from gp;
                D2D    : out Vec2d from gp);
    
	---Purpose: Returns the value and the first derivatives in
	--          the parametric space of the surface S of the point
	--          at parameter X on the arc A.


    Resolution(myclass; A: TheArc; Tol3d: Real from Standard)

        ---Purpose :  Returns the parametric resolution corresponding
        --         to the space resolution Tol3d.

    	returns Real from Standard;


end ArcTool;
