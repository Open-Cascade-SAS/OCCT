-- Created on: 1993-12-03
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




package BlendFunc

    ---Purpose: This package provides a set of generic functions, that can
    --          instantiated to compute blendings between two surfaces
    --          (Constant radius, Evolutive radius, Ruled surface).


uses Blend, Adaptor2d, Adaptor3d, math, gp, Convert, TColgp, TColStd, GeomAbs, Law

is

    class ConstRad;

    class ConstRadInv;

    class Ruled;

    class RuledInv;

    class EvolRad;

    class EvolRadInv;
    
    class CSConstRad;

    class CSCircular;

    class Corde;

    class Chamfer;

    class ChamfInv;
    
    class ChAsym;
    
    class ChAsymInv;
    
    class Tensor;

    enumeration SectionShape is
    	Rational,         -- default in algoritmes
	QuasiAngular,
	Polynomial,
	Linear            -- for chamfers ??
    end SectionShape;


    GetShape(SectShape: SectionShape from BlendFunc; 
             MaxAng:    Real         from  Standard;
	     NbPoles,NbKnots,Degree : out Integer from Standard;
             TypeConv : out ParameterisationType from Convert);

    Knots(SectShape: SectionShape from BlendFunc; 
    	  TKnots: out Array1OfReal from TColStd);

    Mults(SectShape: SectionShape from BlendFunc; 
    	  TMults: out Array1OfInteger from TColStd);

    GetMinimalWeights(SectShape: SectionShape from BlendFunc;
    	              TConv      : ParameterisationType from Convert;
    	              AngleMin   : Real;
		      AngleMax   : Real;
		      Weigths    : out Array1OfReal  from TColStd);	      
	      
    NextShape(S : Shape from GeomAbs)
	      ---Purpose: Used  to obtain the next level of continuity.
	      ---Level: Internal
	      returns Shape from GeomAbs;

    ComputeNormal(Surf : HSurface from Adaptor3d;
                  p2d : Pnt2d from gp;
                  Normal : out Vec from gp)
    returns Boolean from Standard;

    ComputeDNormal(Surf : HSurface from Adaptor3d;
                   p2d : Pnt2d from gp;
                   Normal, DNu, DNv : out Vec from gp)
    returns Boolean from Standard;
	      
end BlendFunc;
