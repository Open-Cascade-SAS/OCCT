-- Created on: 1991-05-14
-- Created by: Laurent PAINNOT
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class BrentMinimum from math
     ---Purpose:
     -- This class implements the Brent's method to find the minimum of
     -- a function of a single variable.
     -- No knowledge of the derivative is required.

uses Matrix from math, 
     Vector from math,
     Function from math,
     OStream from Standard

raises NotDone from StdFail

is

   Create(TolX: Real; 
          NbIterations: Integer = 100; 
          ZEPS: Real = 1.0e-12)
       ---Purpose:
       -- This constructor should be used in a sub-class to initialize
       -- correctly all the fields of this class. 
   returns BrentMinimum;


   Create(TolX: Real; Fbx: Real;
          NbIterations: Integer = 100; 
          ZEPS: Real = 1.0e-12)
       ---Purpose:
       -- This constructor should be used in a sub-class to initialize
       -- correctly all the fields of this class. 
       -- It has to be used if F(Bx) is known.
   returns BrentMinimum;


   Delete(me) is static;
    ---Purpose: Destructor alias.
    ---C++: inline
    ---C++: alias "  Standard_EXPORT virtual ~math_BrentMinimum();"


    Perform(me: in out; F: in out Function;
            Ax, Bx, Cx: Real)
        ---Purpose:
        -- Brent minimization is performed on function F from a given
        -- bracketing triplet of abscissas Ax, Bx, Cx (such that Bx is
        -- between Ax and Cx, F(Bx) is less than both F(Bx) and F(Cx))
        -- The solution is found when: abs(Xi - Xi-1) <= TolX * abs(Xi) + ZEPS;
    is static;


    IsSolutionReached(me: in out; theFunction: in out Function)
        ---Purpose:
        -- This method is called at the end of each iteration to check if the
        -- solution is found.
        -- It can be redefined in a sub-class to implement a specific test to
        -- stop the iterations.
    ---C++:inline
    returns Boolean is virtual;


    IsDone(me)
    	---Purpose: Returns true if the computations are successful, otherwise returns false.
    	---C++: inline

    returns Boolean
    is static;
    
    
    Location(me)
        ---Purpose: returns the location value of the minimum.
        -- Exception NotDone is raised if the minimum was not found.
    	---C++: inline
    returns Real
    raises NotDone
    is static;
    
    
    Minimum(me)
    	---Purpose: returns the value of the minimum.
        -- Exception NotDone is raised if the minimum was not found.
        ---C++: inline

    returns Real
    raises NotDone
    is static;
    

    NbIterations(me)
    	---Purpose: returns the number of iterations really done during the
        -- computation of the minimum.
        -- Exception NotDone is raised if the minimum was not found.
    	---C++: inline

    returns Integer
    raises NotDone
    is static;


    Dump(me; o: in out OStream)
	---Purpose: Prints on the stream o information on the current state 
    	--          of the object.
    	--          Is used to redefine the operator <<.

    is static;


fields

Done:      Boolean;
a:         Real is protected;
b:         Real is protected;
x:         Real is protected;
fx:        Real is protected;
fv:        Real is protected;
fw:        Real is protected;
iter:      Integer;
XTol:      Real is protected;
EPSZ:      Real is protected;
Itermax:   Integer;
myF:       Boolean;

end BrentMinimum;
