-- Created on: 1994-11-14
-- Created by: Jean Claude VAUTHIER 
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



package StlTransfer 

	---Purpose: The  package   Algorithm  for Meshing   implements
	--          facilities to compute  the Mesh data-structure, as
	--          defined in package StlMesh, from a shape of package
	--          TopoDS.  The triangulation  is  computed  with the
	--          Delaunay      algorithm   implemented in   package
	--          BRepMesh.  The  result   is  stored  in  the  mesh
	--          data-structure Mesh from package StlMesh.
	--          

uses  

    StlMesh,
    TopoDS

is
    BuildIncrementalMesh (Shape      : in      Shape from TopoDS; 
    	       	    	  Deflection : in      Real  from Standard;
    	       	    	  InParallel : in      Boolean from Standard;
    	       	          Mesh       : Mesh  from StlMesh)
     raises ConstructionError;
end StlTransfer;






