-- Created on: 1996-01-05
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class CompositeClassifier from TopOpeBRepBuild
    inherits LoopClassifier from TopOpeBRepBuild

---Purpose: 
-- classify composite Loops, i.e, loops that can be either a Shape, or
-- a block of Elements.

uses
    
    ShapeEnum from TopAbs,
    Shape from TopoDS,
    State from TopAbs,
    Loop from TopOpeBRepBuild,
    BlockBuilder from TopOpeBRepBuild
    
is

    Initialize(BB : BlockBuilder);

    Compare(me : in out; L1,L2 : Loop) returns State from TopAbs
    is redefined;

    CompareShapes(me : in out; B1,B2 : Shape from TopoDS)
    ---Purpose: classify shape <B1> with shape <B2>
    returns State from TopAbs is deferred;
    
    CompareElementToShape(me : in out; E,B : Shape from TopoDS)
    ---Purpose: classify element <E> with shape <B>
    returns State from TopAbs is deferred;
    
    ResetShape(me : in out; B : Shape from TopoDS) is deferred;
    ---Purpose: prepare classification involving shape <B>
    -- calls ResetElement on first element of <B>
    
    ResetElement(me : in out; E : Shape from TopoDS) is deferred;
    ---Purpose: prepare classification involving element <E>.
    
    CompareElement(me : in out; E : Shape from TopoDS)  
    returns Boolean from Standard 
    is deferred;
    ---Purpose: Add element <E> in the set of elements used in classification.  
    --  Returns FALSE if the element <E> has been already added to the set of elements, 
    --  otherwise returns TRUE.
     
    State(me : in out) returns State from TopAbs is deferred;
    ---Purpose: Returns state of classification of 2D point, defined by 
    -- ResetElement, with the current set of elements, defined by Compare.

fields

    myBlockBuilder : Address is protected; -- (TopOpeBRepBuild_BlockBuilder*)

end CompositeClassifier from TopOpeBRepBuild;
