-- Created on: 1993-09-06
-- Created by: Christian CAILLET
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class ReadWriteModule  from IGESBasic   inherits ReadWriteModule from IGESData

    ---Purpose : Defines basic File Access Module for IGESBasic (specific parts)
    --           Specific actions concern : Read and Write Own Parameters of
    --           an IGESEntity.

uses Transient, FileReaderData,
     IGESEntity, DirPart, IGESReaderData, ParamReader, IGESWriter

raises DomainError

is

    Create returns mutable ReadWriteModule from IGESBasic;
    ---Purpose : Creates a ReadWriteModule & puts it into ReaderLib & WriterLib

    CaseIGES (me; typenum, formnum : Integer) returns Integer;
    ---Purpose : Defines Case Numbers for Entities of IGESBasic

    ReadOwnParams (me; CN : Integer; ent : mutable IGESEntity;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError;
    ---Purpose : Reads own parameters from file for an Entity of IGESBasic

    WriteOwnParams (me; CN : Integer;  ent : IGESEntity;
    	    	    IW : in out IGESWriter);
    ---Purpose : Writes own parameters to IGESWriter

end ReadWriteModule;
