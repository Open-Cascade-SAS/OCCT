-- Created on: 1996-02-06
-- Created by: Robert COUBLANC
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SensitiveCircle from Select3D 
inherits SensitivePoly from Select3D

    ---Purpose: A framework to define sensitive 3D arcs and circles. 
    -- In some cases this class can raise Standard_ConstructionError and 
    -- Standard_OutOfRange exceptions. For more details see Select3D_SensitivePoly.
uses
    Pnt             from gp,
    Pnt2d           from gp,
    Projector       from Select3D,
    Lin             from gp,
    EntityOwner     from SelectBasics,
    ListOfBox2d     from SelectBasics,
    PickArgs        from SelectBasics,
    Circle          from Geom,
    Array1OfPnt     from TColgp,
    HArray1OfPnt    from TColgp,
    Array1OfPnt2d   from TColgp,
    Box2d           from Bnd,
    Location        from TopLoc,
    Pnt             from Select3D, 
    Pnt2d           from Select3D, 
    Projector       from Select3D,
    SensitiveEntity from Select3D, 
    Circle          from Geom

raises
    ConstructionError from Standard,
    OutOfRange from Standard

is
    Create (OwnerId      : EntityOwner from SelectBasics;
            TheCircle    : Circle from Geom;
            FilledCircle : Boolean = Standard_False;
            NbOfPoints   : Integer = 6)
     returns mutable SensitiveCircle;
        ---Level: Public 
        ---Purpose: Constructs the sensitive circle object defined by the
        -- owner OwnerId, the circle Circle, the Boolean
        -- FilledCircle and the number of points NbOfPoints.

    Create (OwnerId      : EntityOwner from SelectBasics;
            TheCircle    : Circle from Geom;
            u1           : Real ;   
            u2           : Real;
            FilledCircle : Boolean = Standard_False;
            NbOfPoints   : Integer = 6)
     returns mutable SensitiveCircle;
        ---Level: Public 
        ---Purpose: Constructs the sensitive arc object defined by the
        -- owner OwnerId, the circle Circle, the parameters u1
        -- and u2, the Boolean FilledCircle and the number of points NbOfPoints.
        -- u1 and u2 define the first and last points of the arc on Circle.

    Create(OwnerId  : EntityOwner from SelectBasics;
           apolyg3d : HArray1OfPnt   from TColgp;
       FilledCircle : Boolean from Standard = Standard_False)
    returns mutable SensitiveCircle;
        ---Level: Internal 
        ---Purpose: Constructs the sensitive circle object defined by the
        -- owner OwnerId, the array of triangles apolyg3d, and the Boolean FilledCircle.
        -- apolyg3d is an array of consecutive triangles on the
        -- circle. The triangle i+1 lies on the intersection of the
        -- tangents to the circle of i and i+2. Note, that the first point of apolyg3d 
        -- must be equal to the last point of apolyg3d. 

    Create(OwnerId  : EntityOwner from SelectBasics;
           apolyg3d : Array1OfPnt   from TColgp;
       FilledCircle : Boolean from Standard = Standard_False)
    returns mutable SensitiveCircle;
        ---Purpose: Constructs the sensitive circle object defined by the
        -- owner OwnerId, the array of points apolyg3d, and the Boolean FilledCircle. 
        -- If the length of apolyg3d is more then 1, the first point of apolyg3d 
        -- must be equal to the last point of apolyg3d. 

    Matches (me : mutable;
             thePickArgs : PickArgs from SelectBasics;
             theMatchDMin, theMatchDepth : out Real from Standard)
    returns Boolean is redefined static;
    ---Level: Public
    ---Purpose: Checks whether the sensitive entity matches the picking
    -- detection area (close to the picking line).
    -- For details please refer to base class declaration.

    Matches (me  :mutable; 
             XMin,YMin,XMax,YMax : Real from Standard;
             aTol: Real from Standard)
    returns Boolean
    is redefined static;
     
    Matches (me  :mutable; 
             Polyline:Array1OfPnt2d from TColgp;
             aBox:Box2d from Bnd;
             aTol: Real from Standard) 
    returns Boolean
    is redefined virtual;
        ---Level: Public 
    

    ComputeDepth (me;
                  thePickLine : Lin from gp;
                  theDetectedIndex : Integer from Standard)
    returns Real from Standard;
    ---Level: Public
    ---Purpose: Compute depth of sensitive circle for the detected sub-part.
    -- @param thePickLine [in] the picking line.
    -- @param theDetectedIndex [in] index of the detected sub-part.
    -- @return depth on the picking line.

    ArrayBounds(me;Low,Up:in out Integer);
    
    GetPoint3d(me;rank:Integer) returns Pnt from gp;
        ---Level: Internal 

    Dump(me; S: in out OStream;FullDump : Boolean from Standard = Standard_True) is redefined virtual; 

    GetConnected(me: mutable; theLocation : Location from TopLoc) 
    returns SensitiveEntity from Select3D 
    is redefined virtual; 
        ---Level: Public 
        ---Purpose: Returns the copy of this. 

    Project(me: mutable;aProjector: Projector from Select3D) is redefined virtual;

    ComputeCenter3D(me: mutable) is private; 
        ---Level: Internal 
        ---Purpose: Computes myCenter3D as the barycenter of points from mypolyg3d

fields

    myFillStatus    : Boolean;
    myCenter2D      : Pnt2d from Select3D; -- used for Matches()
    myCenter3D      : Pnt from Select3D; -- used for Matches()
    myCircle        : Circle from Geom;
    mystart         : Real from Standard; -- used for GetConnected() 
    myend           : Real from Standard; -- used for GetConnected()
    
end SensitiveCircle;

