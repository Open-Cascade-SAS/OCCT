-- Created on: 1992-08-26
-- Created by: Remi GILET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MakeTranslation

from gce

    ---Purpose: This class implements elementary construction algorithms for a
    -- translation in 3D space. The result is a gp_Trsf transformation.
    -- A MakeTranslation object provides a framework for:
    -- -   defining the construction of the transformation,
    -- -   implementing the construction algorithm, and
    -- -   consulting the result.

uses Pnt  from gp,
     Trsf from gp,
     Vec  from gp,
     Real from Standard
     
is

Create(Vect : Vec from gp) returns MakeTranslation;
    --- Purpose: Constructs a translation along the vector " Vect"
    
Create(Point1 : Pnt from gp;
       Point2 : Pnt from gp) returns MakeTranslation;
    ---Purpose: Constructs a translation along the vector
    --   (Point1,Point2) defined from the point Point1 to the point Point2.
        
Value(me) returns Trsf from gp
    is static;
    ---C++: return const&
    ---Purpose:
    -- Returns the constructed transformation.

Operator(me) returns Trsf from gp
    is static;
    ---C++: return const&
    ---C++: alias "Standard_EXPORT operator gp_Trsf() const;"

fields

    TheTranslation : Trsf from gp;

end MakeTranslation;

