-- Created on: 1993-07-22
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MakeSphere from BRepPrimAPI  inherits MakeOneAxis from BRepPrimAPI 

	---Purpose: Describes functions to build spheres or portions of spheres.
    	-- A MakeSphere object provides a framework for:
    	-- -   defining the construction of a sphere,
    	-- -   implementing the construction algorithm, and
    	-- -   consulting the result.

uses
    Pnt      from gp,
    Ax2      from gp,
    Sphere   from BRepPrim,
    OneAxis  from BRepPrim

raises
    DomainError from Standard

is
    Create(R : Real)
    returns MakeSphere from BRepPrimAPI
	---Purpose: Make a sphere of radius R.
	---Level: Public

    raises
    	DomainError from Standard; -- if R  <= Precision::Confusion()

    Create(R, angle : Real)
    returns MakeSphere from BRepPrimAPI
	---Purpose: Make a sphere of radius R.
	---Level: Public
    raises
    	DomainError from Standard; -- if R  <= Precision::Confusion()

    Create(R, angle1, angle2 : Real)
    returns MakeSphere from BRepPrimAPI
	---Purpose: Make a sphere of radius R.
	---Level: Public
    raises
    	DomainError from Standard; -- if R  <= Precision::Confusion()

    Create(R, angle1, angle2, angle3 : Real)
    returns MakeSphere from BRepPrimAPI
	---Purpose: Make a sphere of radius R.
	---Level: Public
    raises
    	DomainError from Standard; -- if R  <= Precision::Confusion()

    Create(Center : Pnt from gp; R : Real)
    returns MakeSphere from BRepPrimAPI
	---Purpose: Make a sphere of radius R.
	---Level: Public
    raises
    	DomainError from Standard; -- if R  <= Precision::Confusion()

    Create(Center : Pnt from gp; R, angle : Real)
    returns MakeSphere from BRepPrimAPI
	---Purpose: Make a sphere of radius R.
	---Level: Public
    raises
    	DomainError from Standard; -- if R  <= Precision::Confusion()

    Create(Center : Pnt from gp; R, angle1, angle2 : Real)
    returns MakeSphere from BRepPrimAPI
	---Purpose: Make a sphere of radius R.
	---Level: Public
    raises
    	DomainError from Standard; -- if R  <= Precision::Confusion()

    Create(Center : Pnt from gp; R, angle1, angle2, angle3 : Real)
    returns MakeSphere from BRepPrimAPI
	---Purpose: Make a sphere of radius R.
	---Level: Public
    raises
    	DomainError from Standard; -- if R  <= Precision::Confusion()

    Create(Axis : Ax2 from gp; R : Real)
    returns MakeSphere from BRepPrimAPI
	---Purpose: Make a sphere of radius R.
	---Level: Public
    raises
    	DomainError from Standard; -- if R  <= Precision::Confusion()

    Create(Axis : Ax2 from gp; R, angle : Real)
    returns MakeSphere from BRepPrimAPI
	---Purpose: Make a sphere of radius R.
	---Level: Public
    raises
    	DomainError from Standard; -- if R  <= Precision::Confusion()

    Create(Axis : Ax2 from gp; R, angle1, angle2 : Real)
    returns MakeSphere from BRepPrimAPI
	---Purpose: Make a sphere of radius R.
	---Level: Public
    raises
    	DomainError from Standard; -- if R  <= Precision::Confusion()

    Create(Axis : Ax2 from gp; R, angle1, angle2, angle3 : Real)
    returns MakeSphere from BRepPrimAPI
	---Purpose: Make a sphere of radius R.
	---Level: Public
    raises
    	DomainError from Standard; -- if R  <= Precision::Confusion()
    
    	---Purpose: For all algorithms The resulting shape is composed of
    	-- -   a lateral spherical face,
    	-- -   two planar faces parallel to the plane z = 0 if the
    	--   sphere is truncated in the v parametric direction, or
    	--   only one planar face if angle1 is equal to -p/2 or if
    	--     angle2 is equal to p/2 (these faces are circles in
    	--   case of a complete truncated sphere),
    	-- -   and in case of a portion of sphere, two planar faces
    	--   to shut the shape.(in the planes u = 0 and u = angle).   

    OneAxis(me : in out) returns Address;
	---Purpose: Returns the algorithm.
	---Level: Advanced

    Sphere(me : in out) returns Sphere from BRepPrim
	---Purpose: Returns the algorithm.
	--          
	---C++: return &
	---Level: Public 
    is static;

fields

    mySphere : Sphere from BRepPrim;

end MakeSphere;
