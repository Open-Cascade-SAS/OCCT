-- Created on: 1995-05-10
-- Created by: Denis PASCAL
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package PDataStd 

	---Purpose: 


uses Standard,
     PDF,
     PCollection,
     PColStd,
     TColStd


is


    ---Purpose: General Data
    --          ============

    class Name;
    
    class Comment;
    
    ---Purpose: Basic Data for Modeling
    --          =======================

    class Integer; 
    
    class IntegerArray; 
     
    class IntegerArray_1; 
    
    class Real;

    class RealArray; 
    
    class RealArray_1;     
    
    class ExtStringArray; 
     
    class ExtStringArray_1;

    class TreeNode;	    
    
    class Expression;
    
    class Relation;
    
    class Variable;
    
    ---Purpose: Document Data for Modeling
    --          ==========================
    
    class NoteBook; 
 
    class UAttribute;
        
    class Directory;

     
    -- Extension    
    class Tick;
    
    -- Lists:
    class IntegerList;
    class RealList;
    class ExtStringList;
    class BooleanList;
    class ReferenceList;

    -- Arrays:
    class BooleanArray;
    class ReferenceArray;
    class ByteArray;
    class ByteArray_1; 
    
    class NamedData; 
    class AsciiString; 
    class IntPackedMap;  
    class IntPackedMap_1;
     

    class HArray1OfHAsciiString instantiates
    	    	    HArray1 from PCollection (HAsciiString from PCollection);

        class HArray1OfHArray1OfInteger instantiates HArray1 from  PCollection( 
		HArray1OfInteger  from  PColStd); 
		 
	class HArray1OfHArray1OfReal instantiates HArray1 from  PCollection( 
		HArray1OfReal  from  PColStd); 
		 
	class HArray1OfByte instantiates HArray1 from  PCollection( 
		Byte  from  Standard);   
		
end PDataStd;
