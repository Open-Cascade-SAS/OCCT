-- Created on: 2003-02-04
-- Created by: data exchange team
-- Copyright (c) 2003-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class ElementGeometricRelationship from StepFEA
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity ElementGeometricRelationship

uses
    ElementOrElementGroup from StepFEA,
    AnalysisItemWithinRepresentation from StepElement,
    ElementAspect from StepElement

is
    Create returns ElementGeometricRelationship from StepFEA;
	---Purpose: Empty constructor

    Init (me: mutable; aElementRef: ElementOrElementGroup from StepFEA;
                       aItem: AnalysisItemWithinRepresentation from StepElement;
                       aAspect: ElementAspect from StepElement);
	---Purpose: Initialize all fields (own and inherited)

    ElementRef (me) returns ElementOrElementGroup from StepFEA;
	---Purpose: Returns field ElementRef
    SetElementRef (me: mutable; ElementRef: ElementOrElementGroup from StepFEA);
	---Purpose: Set field ElementRef

    Item (me) returns AnalysisItemWithinRepresentation from StepElement;
	---Purpose: Returns field Item
    SetItem (me: mutable; Item: AnalysisItemWithinRepresentation from StepElement);
	---Purpose: Set field Item

    Aspect (me) returns ElementAspect from StepElement;
	---Purpose: Returns field Aspect
    SetAspect (me: mutable; Aspect: ElementAspect from StepElement);
	---Purpose: Set field Aspect

fields
    theElementRef: ElementOrElementGroup from StepFEA;
    theItem: AnalysisItemWithinRepresentation from StepElement;
    theAspect: ElementAspect from StepElement;

end ElementGeometricRelationship;
