-- File:	IGESDraw_ToolDrawing.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolDrawing  from IGESDraw

    ---Purpose : Tool to work on a Drawing. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses Drawing from IGESDraw,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolDrawing;
    ---Purpose : Returns a ToolDrawing, ready to work


    ReadOwnParams (me; ent : mutable Drawing;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : Drawing;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : Drawing;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a Drawing <ent>, from
    --           its specific (own) parameters

    OwnCorrect (me; ent : mutable Drawing) returns Boolean  is static;
    ---Purpose : Sets automatic unambiguous Correction on a Drawing
    --           (Null Views are removed from list)

    DirChecker (me; ent : Drawing) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : Drawing;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : Drawing; entto : mutable Drawing;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : Drawing;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolDrawing;
