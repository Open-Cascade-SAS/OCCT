-- Created on: 1994-05-31
-- Created by: Christian CAILLET
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class SelectName  from IGESSelect  inherits  SelectExtract

    ---Purpose : Selects Entities which have a given name.
    --           Consider Property Name if present, else Short Label, but
    --           not the Subscript Number
    --           First version : keeps exact name
    --           Later : regular expression

uses AsciiString from TCollection, HAsciiString from TCollection,
     Transient, InterfaceModel

is

    Create returns mutable SelectName;
    ---Purpose : Creates an empty SelectName : every entity is considered
    --           good (no filter active)

    Sort (me; rank : Integer; ent : Transient; model : InterfaceModel)
    	returns Boolean;
    ---Purpose : Returns True if Name of Entity complies with Name Filter

    SetName (me : mutable; name : HAsciiString from TCollection);
    ---Purpose : Sets a Name as a criterium : IGES Entities which have this name
    --           are kept (without regular expression, there should be at most
    --           one). <name> can be regarded as a Text Parameter

    Name (me) returns HAsciiString from TCollection;
    ---Purpose : Returns the Name used as Filter

    ExtractLabel (me) returns AsciiString from TCollection;
    ---Purpose : Returns the Selection criterium : "IGES Entity, Name : <name>"

fields

    thename : HAsciiString from TCollection;

end SelectName;
