-- File:	IGESSolid_ToolConicalSurface.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolConicalSurface  from IGESSolid

    ---Purpose : Tool to work on a ConicalSurface. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses ConicalSurface from IGESSolid,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolConicalSurface;
    ---Purpose : Returns a ToolConicalSurface, ready to work


    ReadOwnParams (me; ent : mutable ConicalSurface;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : ConicalSurface;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : ConicalSurface;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a ConicalSurface <ent>, from
    --           its specific (own) parameters

    DirChecker (me; ent : ConicalSurface) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : ConicalSurface;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : ConicalSurface; entto : mutable ConicalSurface;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : ConicalSurface;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolConicalSurface;
