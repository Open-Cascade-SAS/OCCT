-- Created on: 1993-03-23
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class LoopSet from TopOpeBRepBuild

uses

    Loop                     from TopOpeBRepBuild,
    ListOfLoop               from TopOpeBRepBuild,
    ListIteratorOfListOfLoop from TopOpeBRepBuild

is
    
    Create returns LoopSet;
    
    Delete(me:out) is virtual;
    ---C++: alias "Standard_EXPORT virtual ~TopOpeBRepBuild_LoopSet(){Delete() ; }"
    
    -- filling : append loops (shapes,blocks) in list
    ChangeListOfLoop(me : in out) returns ListOfLoop is static;
    ---C++: return &

    -- exploration of the loops
    InitLoop(me : in out) is virtual;
    MoreLoop(me) returns Boolean is virtual;
    NextLoop(me : in out) is virtual;
    Loop(me) returns Loop from TopOpeBRepBuild is virtual;
    ---C++: return const &
    
fields

    myListOfLoop : ListOfLoop;
    myLoopIterator : ListIteratorOfListOfLoop;
    myLoopIndex : Integer from Standard;
    myNbLoop : Integer from Standard;
    
end LoopSet from TopOpeBRepBuild;
