-- Created on: 1997-01-20
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


package TestTopOpeDraw

uses 

    TopoDS,
    Draw,
    DrawTrSurf,
    DBRep,
    TCollection,
    Geom2d,
    Geom,
    gp,
    TestTopOpeTools,
    Standard,
    TColgp
        
is
    
    class ListOfPnt2d instantiates List from TCollection(Pnt2d from gp);
    class DrawableSHA;
    class DrawableSUR;
    class DrawableC3D;
    class DrawableC2D;
    class DrawableP3D;
    class Array1OfDrawableP3D instantiates Array1 from TCollection
    (DrawableP3D from TestTopOpeDraw);
    class HArray1OfDrawableP3D instantiates HArray1 from TCollection
    (DrawableP3D from TestTopOpeDraw,Array1OfDrawableP3D from TestTopOpeDraw);
    class DrawableP2D;

    class DrawableMesure;
    class Array1OfDrawableMesure instantiates Array1 from TCollection
    (DrawableMesure from TestTopOpeDraw);
    class HArray1OfDrawableMesure instantiates HArray1 from TCollection
    (DrawableMesure from TestTopOpeDraw,
     Array1OfDrawableMesure from TestTopOpeDraw);

    AllCommands(I : in out Interpretor from Draw);
    OtherCommands(I : in out Interpretor from Draw);

end TestTopOpeDraw;
