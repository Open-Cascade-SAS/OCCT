-- Created on: 1999-03-24
-- Created by: data exchange team
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class AssemblyLink from STEPSelections inherits TShared from MMgt

	---Purpose: 

uses
    
    NextAssemblyUsageOccurrence from StepRepr,
    ContextDependentShapeRepresentation from StepShape,
    AssemblyComponent from STEPSelections

is

    Create returns mutable AssemblyLink from STEPSelections;
    
    Create(nauo: NextAssemblyUsageOccurrence from StepRepr;
    	   item: Transient from Standard;
	   part: AssemblyComponent from STEPSelections)
    returns mutable AssemblyLink from STEPSelections;
    
    --Methods for setting and obtaining fields
    
    GetNAUO(me) returns NextAssemblyUsageOccurrence from StepRepr;
    	---Purpose:
	---C++: inline
	
    GetItem(me) returns Transient from Standard;
    	---Purpose:
	---C++: inline
	
    GetComponent(me) returns AssemblyComponent from STEPSelections;
    	---Purpose:
	---C++: inline
    
    SetNAUO(me: mutable; nauo: NextAssemblyUsageOccurrence from StepRepr);
    	---Purpose:
	---C++: inline
	
    SetItem(me: mutable; item: Transient from Standard);
    	---Purpose:
	---C++: inline
    
    SetComponent(me: mutable; part: AssemblyComponent from STEPSelections);
	---Purpose:
	---C++: inline

fields

    myNAUO     : NextAssemblyUsageOccurrence from StepRepr;
    myItem     : Transient from Standard;
    myComponent: AssemblyComponent from STEPSelections;

end AssemblyLink;
