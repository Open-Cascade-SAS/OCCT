-- Created on: 1998-03-04
-- Created by: Julia Gerasimova
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class BadEdgeFilter from AIS inherits Filter from SelectMgr

	---Purpose: A Class

uses

    EntityOwner                    from SelectMgr,
    Edge                           from TopoDS,
    DataMapOfIntegerListOfShape    from TopTools,    
    ShapeEnum                      from TopAbs
    
is
    Create
    returns mutable BadEdgeFilter from AIS;
    	--- Purpose: Constructs an empty filter object for bad edges.   
    ActsOn( me; aType : ShapeEnum from TopAbs )
    returns Boolean from Standard
    is redefined;
    
    IsOk( me; EO : EntityOwner from SelectMgr )
    returns Boolean from Standard is redefined virtual;

    SetContour( me : mutable ; Index : Integer from Standard );
    	---Purpose: sets  <myContour> with  current  contour. used  by
    	--          IsOk.

    AddEdge( me: mutable ; anEdge : Edge from TopoDS;
    	    	    	   Index : Integer from Standard );
    	---Purpose:  Adds an  edge  to the list  of non-selectionnable
    	--          edges.

    RemoveEdges( me: mutable ; Index : Integer from Standard );
    	---Purpose: removes from the  list of non-selectionnable edges
    	--          all edges in the contour <Index>.

fields

    myBadEdges : DataMapOfIntegerListOfShape from TopTools;
    myContour  : Integer                     from Standard;

end BadEdgeFilter;
