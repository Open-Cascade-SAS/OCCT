-- File:	BndLib_Add3dCurve.cdl
-- Created:	Thu Jul  8 17:29:02 1993
-- Author:	Isabelle GRIGNON
--		<isg@sdsun2>
---Copyright:	 Matra Datavision 1993


class Add3dCurve from BndLib 
    	---Purpose: Computes the bounding box for a curve in 3d.
    	-- Functions to add a 3D curve to a bounding box.
    	-- The 3D curve is defined from a Geom curve.
        
uses Box   from Bnd,
     Curve from Adaptor3d

is
    Add(myclass; C   :        Curve from Adaptor3d;
    	    	 Tol :        Real  from Standard; 
    	    	 B   : in out Box   from Bnd);
    	---Purpose: Adds to the bounding box B the curve C
    	-- B is then enlarged by the tolerance value Tol.
    	-- Note: depending on the type of curve, one of the following
    	-- representations of the curve C is used to include it in the bounding box B:
    	-- -   an exact representation if C is built from a line, a circle   or a conic curve,
    	-- -   the poles of the curve if C is built from a Bezier curve or   a BSpline curve,
    	---   if not, the points of an approximation of the curve C.
    	-- Warning
    	-- C is an adapted curve, that is, an object which is an interface between:
    	-- -   the services provided by a 3D curve from the package   Geom
    	-- -   and those required of the curve by the computation algorithm.
    	--  The adapted curve is created in the following way:
    	--    Handle(Geom_Curve) mycurve = ... ;
    	--    GeomAdaptor_Curve C(mycurve);
    	-- The bounding box B is then enlarged by adding it:
    	--    Bnd_Box B;
    	-- // ...
    	--    Standard_Real Tol = ... ;
    	--    Add3dCurve::Add ( C, Tol, B );
    	-- Exceptions
    	-- Standard_Failure if the curve is built from:
    	-- -   a Geom_Line, or
    	-- -   a Geom_Parabola, or
    	-- -   a Geom_Hyperbola,
    	-- and P1 and P2 are either two negative infinite real
    	-- numbers, or two positive infinite real numbers.
    
    
    
    Add(myclass; C     :        Curve from Adaptor3d; 
    	    	 U1,U2 :        Real  from Standard;
    	         Tol   :        Real  from Standard;
    	         B     : in out Box   from Bnd);
    	---Purpose: Adds to the bounding box B the curve C
    	-- the arc of the curve C limited by the two parameter values P1 and P2.
 	-- Note: depending on the type of curve, one of the following
    	-- representations of the curve C is used to include it in the bounding box B:
    	-- -   an exact representation if C is built from a line, a circle   or a conic curve,
    	-- -   the poles of the curve if C is built from a Bezier curve or   a BSpline curve,
    	---   if not, the points of an approximation of the curve C.
    	-- Warning
    	-- C is an adapted curve, that is, an object which is an interface between:
    	-- -   the services provided by a 3D curve from the package   Geom
    	-- -   and those required of the curve by the computation algorithm.
    	--  The adapted curve is created in the following way:
    	--    Handle(Geom_Curve) mycurve = ... ;
    	--    GeomAdaptor_Curve C(mycurve);
    	-- The bounding box B is then enlarged by adding it:
    	--    Bnd_Box B;
    	-- // ...
    	--    Standard_Real Tol = ... ;
    	--    Add3dCurve::Add ( C, Tol, B );
    	-- Exceptions
    	-- Standard_Failure if the curve is built from:
    	-- -   a Geom_Line, or
    	-- -   a Geom_Parabola, or
    	-- -   a Geom_Hyperbola,
    	-- and P1 and P2 are either two negative infinite real
    	-- numbers, or two positive infinite real numbers.
  
end Add3dCurve;
