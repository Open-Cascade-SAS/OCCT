-- Created on: 1992-08-27
-- Created by: Christophe MARION
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class DrawableEdgeTool from HLRTest inherits Drawable3D from Draw

	---Purpose: 

uses
    Boolean  from Standard,
    Integer  from Standard,
    Display  from Draw,
    Algo     from HLRBRep,
    Data     from HLRBRep,
    EdgeData from HLRBRep

is
    Create(Alg     : Algo    from HLRBRep;
           Visible : Boolean from Standard;
           IsoLine : Boolean from Standard;
           Rg1Line : Boolean from Standard;
           RgNLine : Boolean from Standard;
           ViewId  : Integer from Standard)
    returns mutable DrawableEdgeTool from HLRTest;
    
    DrawOn(me; D : in out Display from Draw);
    
    InternalDraw(me; D   :in out Display from Draw;
                     typ :       Integer from Standard)
    is static private;
    
    DrawFace(me; D      : in out Display from Draw;
                 typ    :        Integer from Standard;
                 nCB    :        Integer from Standard;
                 iface  :        Integer from Standard;
		 e2,iCB : in out Integer from Standard;
                 DS     : in out Data    from HLRBRep)
    is static private;
    
    DrawEdge(me; D      : in out Display  from Draw;
                 inFace :        Boolean  from Standard;
                 typ    :        Integer  from Standard;
                 nCB    :        Integer  from Standard;
                 ie     :        Integer  from Standard;
		 e2,iCB : in out Integer  from Standard;
                 ed     : in out EdgeData from HLRBRep)
    is static private;
    
fields
    myAlgo    : Algo    from HLRBRep;
    myVisible : Boolean from Standard;
    myIsoLine : Boolean from Standard;
    myRg1Line : Boolean from Standard;
    myRgNLine : Boolean from Standard;
    myViewId  : Integer from Standard;

end DrawableEdgeTool;
