-- File:	QARina.cdl
-- Created:	Tue Mar 19 09:16:47 2002
-- Author:	QA Admin
--		<qa@umnox.nnov.matra-dtv.fr>
---Copyright:	 Matra Datavision 2002

package QARina
     uses Draw
is
    Commands(DI : in out Interpretor from Draw);
end;
    
