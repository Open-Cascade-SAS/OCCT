-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class EdgeLoop from StepShape 

inherits Loop from StepShape 
-- WARNING : Multiple EXPRESS inheritance
-- Not yet automaticly managed
-- inherits Path from StepShape 


-- Hand made changes : All the attributes theoricly inherited from the Path
-- entity are explicitly declared in the EdgeLoop entity.
-- The path is not directly referenced by any other entities. As far as
-- Path supertype, topological representation item, is also a 
-- supertype of Edge, this mapping is equivalent.

uses

    	HAsciiString          from TCollection,
	HArray1OfOrientedEdge from StepShape, 
	OrientedEdge          from StepShape

is

	Create returns mutable EdgeLoop;
	---Purpose: Returns a EdgeLoop

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aEdgeList : mutable HArray1OfOrientedEdge from StepShape);

	-- Specific Methods for Field Data Access --

	SetEdgeList(me : mutable; aEdgeList : mutable HArray1OfOrientedEdge);
	EdgeList (me) returns mutable HArray1OfOrientedEdge;
	EdgeListValue (me; num : Integer) returns mutable OrientedEdge;
	NbEdgeList (me) returns Integer;

fields

	edgeList : HArray1OfOrientedEdge from StepShape;

end EdgeLoop;
