-- File:	StepToGeom_MakeConic.cdl
-- Created:	Mon Jun 21 11:18:38 1993
-- Author:	Martine LANGLOIS
---Copyright:	 Matra Datavision 1993

class MakeConic from StepToGeom

    ---Purpose: This class implements the mapping between classes 
    --          Conic from StepGeom
    --          which describes a Conic from prostep and Conic from Geom .
    --          As Conic is an abstract class
    --          this class is an access to the sub-class required.

uses Conic from Geom,
     Conic from StepGeom

is 

    Convert ( myclass; SC : Conic from StepGeom;
                       CC : out Conic from Geom )
    returns Boolean from Standard;

end MakeConic;
