-- Created on: 1997-03-27
-- Created by: Denis PASCAL
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package DDataStd 

	---Purpose: commands for Standard Attributes.
	--          =================================


uses Draw,
     TDF,
     TDataStd,     
     TDataXtd,
     TopoDS,
     MMgt,
     Standard,
     TNaming, 
     TCollection

is 

    class DrawPresentation;
    
    class DrawDriver;

    class TreeBrowser;
    ---Purpose: Used to browse tree nodes.

    ---Purpose: commands
    --          ========

    AllCommands (I : in out Interpretor from Draw);
    ---Purpose: command to set and get modeling attributes

    NamedShapeCommands (I : in out Interpretor from Draw);
    ---Purpose: to set and get NamedShape

    BasicCommands  (I : in out Interpretor from Draw);
    ---Purpose: to set and get Integer, Real,  Reference, Geometry

    DatumCommands (I : in out Interpretor from Draw);
    ---Purpose: to set and get Datum attributes

    ConstraintCommands (I : in out Interpretor from Draw);
    ---Purpose: to set and get Constraint and Constraint  attributes    

    ObjectCommands (I : in out Interpretor from Draw);
    ---Purpose: to set and get Objects attributes

    DrawDisplayCommands  (I : in out Interpretor from Draw);
    ---Purpose: to display standard attributes

    NameCommands (I: in out Interpretor from Draw);
    ---Purpose: to set and get Name attribute    
    
    TreeCommands (I: in out Interpretor from Draw);    
    ---Purpose: to build, edit and browse an explicit tree of labels
    
    ---Purpose: package methods
    --          ===============

    DumpConstraint (C : Constraint from TDataXtd; S : in out OStream);


end DDataStd;

