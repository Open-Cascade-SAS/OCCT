-- Created on: 1993-06-11
-- Created by: Martine LANGLOIS
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


package GeomToStep

--- Purpose: Creation des entites geometriques du schema PmsAp2Demo3d a 
--  partir des entites de Geom ou de gp.
--  Update : mise a jour pour traiter le schema StepGeom, pour demo de 94

uses gp, Geom, Geom2d, StepGeom, StdFail, TColgp

is

private deferred class Root;
class MakeCartesianPoint;
class MakeAxis1Placement;
class MakeAxis2Placement2d;
class MakeAxis2Placement3d;
class MakeDirection;
class MakeVector;
class MakeCurve;
class MakeConic;
class MakeBoundedCurve;
class MakeCircle;
class MakeEllipse;
class MakeHyperbola;
class MakeParabola;
class MakeBSplineCurveWithKnots;
class MakeBSplineCurveWithKnotsAndRationalBSplineCurve;
class MakeLine;
class MakePolyline;
class MakePlane;
class MakeSurface;
class MakeBoundedSurface;
class MakeElementarySurface;
class MakeSweptSurface;
class MakeConicalSurface;
class MakeCylindricalSurface;
class MakeRectangularTrimmedSurface;
class MakeSphericalSurface;
class MakeSurfaceOfLinearExtrusion;
class MakeSurfaceOfRevolution;
class MakeToroidalSurface;
class MakeBSplineSurfaceWithKnots;
class MakeBSplineSurfaceWithKnotsAndRationalBSplineSurface;

end GeomToStep;
