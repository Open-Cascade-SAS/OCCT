-- Created on: 1998-03-12
-- Created by: Pierre BARRAS
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class SplitCurve from ShapeUpgrade inherits TShared from MMgt

    	---Purpose: Splits a  curve with a  criterion.
    
uses     
    Curve          from Geom,
    HArray1OfCurve from TColGeom,
    HSequenceOfReal  from TColStd,
    Shape          from GeomAbs,
    Status         from  ShapeExtend
is 
 
    Create returns mutable SplitCurve from ShapeUpgrade;
    	---Purpose: Empty constructor.

    Init (me: mutable; First, Last: Real);
    	---Purpose: Initializes with curve first and last parameters.
	
    SetSplitValues (me: mutable; SplitValues: HSequenceOfReal from TColStd);
    	---Purpose: Sets the parameters where splitting has to be done.
	
    Build (me: mutable; Segment: Boolean) is virtual;
       ---Purpose: If Segment is True, the result is composed with
       --  segments of the curve bounded by the SplitValues.  If
       --  Segment is False, the result is composed with trimmed
       --  Curves all based on the same complete curve.
       --  

    SplitValues(me) returns HSequenceOfReal from TColStd;
       ---C++: return const &
       --- Purpose : returns all the splitting values including the  
       --  First and Last parameters of the input curve

       
    ---Level: Internal
    
    --PrepareKnots (me: mutable) is protected;
    	---Purpose: Merges input split values and new ones into myGlobalKnots
    
    Compute(me: mutable) is virtual;
    	---Purpose: Calculates points for correction/splitting of the curve
    
    Perform(me: mutable; Segment: Boolean = Standard_True);
    	---Purpose: Performs correction/splitting of the curve.
	---         First defines splitting values by method Compute(), then calls method Build().   
	
    Status (me; status: Status from ShapeExtend) returns Boolean;
    	---Purpose: Returns the status 
	-- OK    - no splitting is needed
	-- DONE1 - splitting required and gives more than one segment
	-- DONE2 - splitting is required, but gives only one segment (initial)
	-- DONE3 - geometric form of the curve or parametrisation is modified
fields 
 
    mySplitValues     : HSequenceOfReal from TColStd is protected;  
    myNbCurves        : Integer is protected;
    myStatus : Integer is protected; 
end;
    
