-- Created on: 1997-02-12
-- Created by: Alexander BRIVIN
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Scale from Vrml 

	---Purpose: defines a Scale node of VRML specifying transform
	---          properties.
    	--  This  node  defines  a  3D  scaling  about  the  origin. 
    	--  By  default  : 
	--    myRotation  =  (1 1 1)

uses
 
    Vec  from  gp 

is
    Create returns Scale from Vrml;
 
    Create  (  aScaleFactor  :  Vec  from  gp ) 
    	returns Scale from Vrml;

    SetScaleFactor ( me : in out; aScaleFactor : Vec  from  gp );
    ScaleFactor ( me )  returns   Vec  from  gp;

    Print  ( me;  anOStream: in out OStream from Standard) returns OStream from Standard;
    ---C++:  return  & 

fields
 
    myScaleFactor  :  Vec  from  gp;  -- Scale factors in x, y, and z

end Scale;
