-- Created on: 1993-06-23
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class Surface from TopOpeBRepDS

    ---Purpose: A Geom poimt and a tolerance.

uses

    Surface from Geom

is

    Create returns Surface from TopOpeBRepDS; 
    
    Create(P : Surface from Geom; T : Real from Standard)
    returns Surface from TopOpeBRepDS; 
     
--modified by NIZNHY-PKV Tue Oct 30 09:27:32 2001  f    
    Create  (Other :Surface from TopOpeBRepDS) 
    	returns Surface from TopOpeBRepDS; 
	 
    Assign(me :out;  
    	    Other: Surface from TopOpeBRepDS);  
    ---C++: alias operator=
--modified by NIZNHY-PKV Tue Oct 30 09:27:25 2001  t     

    Surface(me) returns Surface from Geom
	---C++: return const &
    is static;
    
    Tolerance(me) returns Real from Standard
    is static;

    Tolerance(me : in out; tol : Real)
    ---Purpose: Update the tolerance
    is static;
	
    Keep(me) returns Boolean from Standard
    is static;
    ChangeKeep(me : in out; B : Boolean from Standard)
    is static;

fields

    mySurface   : Surface from Geom;
    myTolerance : Real from Standard;
    myKeep      : Boolean from Standard;

end Surface from TopOpeBRepDS;
