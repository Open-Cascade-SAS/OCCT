-- File:	RWStepRepr_RWPropertyDefinitionRepresentation.cdl
-- Created:	Thu Dec 12 17:15:59 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWPropertyDefinitionRepresentation from RWStepRepr

    ---Purpose: Read & Write tool for PropertyDefinitionRepresentation

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    PropertyDefinitionRepresentation from StepRepr

is
    Create returns RWPropertyDefinitionRepresentation from RWStepRepr;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : PropertyDefinitionRepresentation from StepRepr);
	---Purpose: Reads PropertyDefinitionRepresentation

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: PropertyDefinitionRepresentation from StepRepr);
	---Purpose: Writes PropertyDefinitionRepresentation

    Share (me; ent : PropertyDefinitionRepresentation from StepRepr;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWPropertyDefinitionRepresentation;
