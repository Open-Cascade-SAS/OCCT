-- Created on: 1997-10-07
-- Created by: Laurent BUCHARD
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class Tool from BRepTopAdaptor 

uses 
    Face       from TopoDS,
    TopolTool  from BRepTopAdaptor,
    HSurface   from Adaptor3d


is 

  Create
     returns Tool from BRepTopAdaptor;

  Create(F     : Face from TopoDS;
    	 Tol2d : Real from Standard)
     returns Tool from BRepTopAdaptor;
     
  Create(Surface: HSurface from Adaptor3d;
         Tol2d  : Real from Standard)
     returns Tool from BRepTopAdaptor;
 
 
  Init(me    : in out;
       F     : Face from TopoDS;
       Tol2d : Real from Standard);
       
  Init(me     : in out;
       Surface: HSurface from Adaptor3d;
       Tol2d  : Real from Standard);       
	  
  ---- 

  GetTopolTool(me: in out) 
     returns mutable TopolTool from BRepTopAdaptor;
     
  SetTopolTool(me: in out ; 
               TT: TopolTool from BRepTopAdaptor);
	
  GetSurface(me: in out)
    returns mutable HSurface from Adaptor3d;
    
	
  ---
	
  Destroy(me: in out) ;
    ---C++: alias ~
    
fields

  myloaded    : Boolean   from Standard;
  myTopolTool : TopolTool from BRepTopAdaptor; 
  myHSurface  : HSurface  from Adaptor3d;

end Tool;
