-- Created on: 1996-04-10
-- Created by: Joelle CHAUVET
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Modified:	Mon Dec  9 10:30:56 1996
--    by:	Joelle CHAUVET
--		G1135 : Empty constructor

class Framework from AdvApp2Var

uses

    Boolean,Real,NoSuchObject from Standard,
    HArray1OfReal from TColStd,
    IsoType from GeomAbs,
    SequenceOfNode,SequenceOfStrip,Iso,Node from AdvApp2Var

raises NoSuchObject from Standard

is

    Create returns Framework;
    Create(Frame : SequenceOfNode; 
           UFrontier, VFrontier : SequenceOfStrip)  
    returns Framework;
    
    FirstNotApprox(me; IndexIso,IndexStrip : out Integer; 
                       anIso : out Iso) 
    ---Purpose: search the Index of the first Iso not approximated,
    --          if all Isos are approximated Standard_False is returned.
    returns Boolean; 

    FirstNode(me; Type : IsoType; IndexIso,IndexStrip : Integer) 
    returns Integer;
    
    LastNode(me; Type : IsoType; IndexIso,IndexStrip : Integer) returns Integer; 
    
    ChangeIso(me: in out; IndexIso,IndexStrip : Integer; anIso : Iso);
    
    Node(me; IndexNode : Integer)
    ---C++: return const&
    ---C++: inline    
    returns Node
    raises NoSuchObject from Standard;
	
    Node(me; U,V : Real) 
    ---C++: return const&
    returns Node
    raises NoSuchObject from Standard;
	
    IsoU(me; U,V0,V1 : Real) 
    ---C++: return const&
    returns Iso
    raises NoSuchObject from Standard;
	
    IsoV(me; U0,U1,V : Real) 
    ---C++: return const&    
    returns Iso
    raises NoSuchObject from Standard;
	
    ChangeNode(me: in out; IndexNode : Integer)
    ---C++: return &
    ---C++: inline    
    returns Node;

    
    UpdateInU(me: in out; CuttingValue : Real);
    
    UpdateInV(me: in out; CuttingValue : Real);
    
    UEquation(me; IndexIso,IndexStrip : Integer) 
    ---C++: return const &
    returns HArray1OfReal; 
    
    VEquation(me; IndexIso,IndexStrip : Integer)
    ---C++: return const & 
     returns HArray1OfReal;
 

fields

    myNodeConstraints    : SequenceOfNode;
    myUConstraints       : SequenceOfStrip;
    myVConstraints       : SequenceOfStrip;

end Framework;

