-- Created on: 1992-05-27
-- Created by: Remi LEQUETTE
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.





class TVertex from BRep inherits TVertex from TopoDS

	---Purpose: The TVertex from  BRep inherits  from  the TVertex
	--          from TopoDS. It contains the geometric data.
	--          
	--          The  TVertex contains a 3d point and a tolerance.
	--            
uses
    Pnt    from gp,
    TShape from TopoDS,
    ListOfPointRepresentation from BRep

is
    Create returns mutable TVertex from BRep;

    Tolerance(me) returns Real
	---C++: inline
    is static;
    
    Tolerance(me : mutable; T : Real)
	---C++: inline
    is static;
    
    UpdateTolerance(me : mutable; T : Real)
	---Purpose: Sets the tolerance  to the   max  of <T>  and  the
	--          current  tolerance.
	--          
	---C++: inline
    is static;

    Pnt(me) returns Pnt from gp
	---C++: inline
	---C++: return const &
    is static;
    
    Pnt(me : mutable; P : Pnt from gp)
	---C++: inline
    is static;
    
    Points(me) returns ListOfPointRepresentation from BRep
	---C++: inline
	---C++: return const &
    is static;
    
    ChangePoints(me : mutable) returns ListOfPointRepresentation from BRep
	---C++: inline
	---C++: return &
    is static;
    
    EmptyCopy(me) returns mutable TShape from TopoDS;
	---Purpose: Returns a copy  of the  TShape  with no sub-shapes.
    
fields

    myPnt       : Pnt from gp;
    myTolerance : Real;
    myPoints    : ListOfPointRepresentation from BRep;

end TVertex;
