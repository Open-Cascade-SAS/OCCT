-- Created on: 1997-10-28
-- Created by: Roman BORISOV
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Curve2d from Approx 

	---Purpose: Makes  an  approximation  for  HCurve2d  from  Adaptor3d

uses
    HCurve2d    from  Adaptor2d, 
    Shape  from  GeomAbs, 
    BSplineCurve  from  Geom2d 
    
is
  Create(C2D  :  HCurve2d    from  Adaptor2d; 
    	 First, 
	 Last, 		      
         TolU,  TolV  :  Real; 
	 Continuity  :  Shape  from  GeomAbs; 
         MaxDegree  :  Integer  ; 
         MaxSegments  :  Integer) 
	      
     returns  Curve2d;	 
      
    IsDone(me) returns Boolean from Standard;
    
    HasResult(me) returns  Boolean from Standard;
   
    Curve(me) 
    returns  BSplineCurve  from  Geom2d; 
     
    MaxError2dU(me) returns  Real;  
    MaxError2dV(me) returns  Real;
    
fields
   
  myCurve            : BSplineCurve  from  Geom2d; 
  myIsDone           : Boolean       from  Standard;   
  myHasResult        : Boolean       from  Standard; 
  myMaxError2dU      : Real          from  Standard; 
  myMaxError2dV      : Real          from  Standard; 
  
end Curve2d;
