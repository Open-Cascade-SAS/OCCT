-- Created on: 1997-10-29
-- Created by: Roman BORISOV
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Assembly from FEmTool

	---Purpose: Assemble and solve system from (one dimensional) Finite Elements  

uses 
    Array2OfInteger  from  TColStd, 
    HAssemblyTable  from  FEmTool, 
    Matrix  from  math, 
    Vector  from  math,	     
    ProfileMatrix  from  FEmTool, 
    SeqOfLinConstr  from  FEmTool, 
    SequenceOfReal  from  TColStd 
    
raises   
        NotDone  from  StdFail, 
        DimensionError, 
	DomainError
is 
    Create(Dependence :  Array2OfInteger  from  TColStd; 
           Table      :  HAssemblyTable  from  FEmTool)   
    returns  Assembly from FEmTool; 
     
    NullifyMatrix(me : in  out); 
    ---Purpose: Nullify all Matrix 's Coefficient
           
    AddMatrix(me  : in  out;   
              Element    :  Integer; 
	      Dimension1 :  Integer; 
	      Dimension2 :  Integer; 
              Mat  :  Matrix  from  math)
    ---Purpose: Add an elementary Matrix in the assembly Matrix 
    	raises  DomainError; --  if  Dependence(Dimension1,Dimension2)  is  False
              
    NullifyVector(me : in  out);                
    ---Purpose:  Nullify  all  Coordinate of  assembly  Vector (second member)
     
    AddVector(me  :  in  out; 
              Element    :  Integer; 
	      Dimension  :  Integer; 
              Vec  :  Vector  from  math);  
    ---Purpose: Add an elementary Vector in the assembly Vector (second member)     

    ResetConstraint(me : in  out);                
    ---Purpose: Delete all Constraints.
    
    NullifyConstraint(me : in  out);                
    ---Purpose: Nullify all Constraints.   
     
    AddConstraint(me : in  out; 
            IndexofConstraint :  Integer;
            Element           :  Integer; 
            Dimension         :  Integer;	     
            LinearForm        :  Vector  from  math;
            Value             :  Real); 
	         
     
    Solve(me  :  in  out)  returns  Boolean; 
    ---Purpose: Solve the assembly system         
    --          Returns Standard_False if the computation failed.
     
    Solution(me;  Solution : out  Vector  from  math) 
    raises  NotDone  from  StdFail;  -- if the system is not solved.  
     
    NbGlobVar(me) 
    returns  Integer; 
     
    GetAssemblyTable(me;  AssTable  :  out  HAssemblyTable  from  FEmTool);
	      
fields  
    myDepTable  :  Array2OfInteger;
    myRefTable  :  HAssemblyTable; 
    IsSolved    :  Boolean;
    H           :  ProfileMatrix  from  FEmTool;  
    B	        :  Vector  from  math;
    GHGt        :  ProfileMatrix  from  FEmTool; 
    G	        :  SeqOfLinConstr  from  FEmTool; 
    C           :  SequenceOfReal  from  TColStd;     
end Assembly;

