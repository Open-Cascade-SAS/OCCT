-- Created on: 2002-01-04
-- Created by: data exchange team
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1

class SeamEdge from StepShape
inherits OrientedEdge from StepShape

    ---Purpose: Representation of STEP entity SeamEdge

uses
    HAsciiString from TCollection,
    Vertex from StepShape,
    Edge from StepShape,
    Pcurve from StepGeom

is
    Create returns SeamEdge from StepShape;
	---Purpose: Empty constructor

    
		       
    Init (me: mutable; aRepresentationItem_Name: HAsciiString from TCollection;	       
                       aOrientedEdge_EdgeElement: Edge from StepShape;
                       aOrientedEdge_Orientation: Boolean;
                       aPcurveReference: Pcurve from StepGeom);
	---Purpose: Initialize all fields (own and inherited)

    PcurveReference (me) returns Pcurve from StepGeom;
	---Purpose: Returns field PcurveReference
    SetPcurveReference (me: mutable; PcurveReference: Pcurve from StepGeom);
	---Purpose: Set field PcurveReference

fields
    thePcurveReference: Pcurve from StepGeom;

end SeamEdge;
