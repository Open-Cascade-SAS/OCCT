-- Created on: 2002-04-09
-- Created by: QA Admin
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PresentableObject from QABugs inherits InteractiveObject from AIS
uses
    Selection from SelectMgr,
    PresentationManager3d from PrsMgr,
    Presentation from Prs3d,
    TypeOfPresentation3d from PrsMgr
is
    
    Create(aTypeOfPresentation3d: TypeOfPresentation3d from PrsMgr = PrsMgr_TOP_AllView) returns PresentableObject from QABugs;
    
    ComputeSelection(me:mutable; aSelection : Selection from SelectMgr;
                                 aMode      : Integer) is redefined virtual protected;

    Compute(me:mutable;
    	    aPresentationManager: PresentationManager3d from PrsMgr;
            aPresentation: Presentation from Prs3d;
            aMode: Integer from Standard = 0)
    is redefined virtual protected;
	    
end PresentableObject;
    
