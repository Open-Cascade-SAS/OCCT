-- Created on: 1997-05-21
-- Created by: Christian CAILLET
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DescrGeneral  from StepData    inherits GeneralModule  from StepData

    ---Purpose : Works with a Protocol by considering its entity descriptions


uses Transient,
     EntityIterator from Interface,
     ShareTool      from Interface,
     Check          from Interface,
     CopyTool       from Interface,
     Protocol  from StepData

is

    Create (proto : Protocol from StepData) returns DescrGeneral;

    FillSharedCase (me; CN : Integer; ent : Transient;
        iter : in out EntityIterator);

    CheckCase (me; CN : Integer; ent : Transient; shares : ShareTool;
    	ach : in out Check);

    CopyCase (me; CN : Integer; entfrom : Transient; entto : mutable Transient;
    	TC : in out CopyTool);

    NewVoid (me; CN : Integer; ent : out mutable Transient) returns Boolean;

fields

    theproto : Protocol from StepData;

end DescrGeneral;
