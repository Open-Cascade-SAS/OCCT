-- Created on: 2002-12-12
-- Created by: data exchange team
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class FeaGroup from StepFEA
inherits Group from StepBasic

    ---Purpose: Representation of STEP entity FeaGroup

uses
    HAsciiString from TCollection,
    FeaModel from StepFEA

is
    Create returns FeaGroup from StepFEA;
	---Purpose: Empty constructor

    Init (me: mutable; aGroup_Name: HAsciiString from TCollection;
                       aGroup_Description: HAsciiString from TCollection;
                       aModelRef: FeaModel from StepFEA);
	---Purpose: Initialize all fields (own and inherited)

    ModelRef (me) returns FeaModel from StepFEA;
	---Purpose: Returns field ModelRef
    SetModelRef (me: mutable; ModelRef: FeaModel from StepFEA);
	---Purpose: Set field ModelRef

fields
    theModelRef: FeaModel from StepFEA;

end FeaGroup;
