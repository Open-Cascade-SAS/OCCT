-- File:        Product.cdl
-- Created:     Mon Dec  4 12:02:29 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWProduct from RWStepBasic

	---Purpose : Read & Write Module for Product

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     Product from StepBasic,
     EntityIterator from Interface

is

	Create returns RWProduct;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable Product from StepBasic);

	WriteStep (me; SW : in out StepWriter; ent : Product from StepBasic);

	Share(me; ent : Product from StepBasic; iter : in out EntityIterator);

end RWProduct;
