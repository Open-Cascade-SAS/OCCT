-- File:	MDataStd_RealStorageDriver.cdl
-- Created:	Wed Apr  9 16:56:00 1997
-- Author:	VAUTHIER Jean-Claude
---Copyright:	 Matra Datavision 1997


class RealStorageDriver from MDataStd inherits ASDriver from MDF

	---Purpose: 

uses SRelocationTable from MDF,
     Attribute        from TDF,
     Attribute        from PDF, 
     MessageDriver    from CDM
is

    Create(theMessageDriver : MessageDriver from CDM) -- Version 0
    returns mutable RealStorageDriver from MDataStd;


    VersionNumber(me) returns Integer from Standard;
	---Purpose: Returns the version number from which the driver
	--          is available: 0.

    SourceType(me) returns Type from Standard;
	---Purpose: Returns the type: Real from TDataStd.

    NewEmpty (me) returns mutable Attribute from PDF;


    Paste(me;
    	  Source     :         Attribute from TDF;
    	  Target     : mutable Attribute from PDF;
    	  RelocTable : SRelocationTable from MDF);


end RealStorageDriver;

