-- File:	StepData_ReadWriteModule.cdl
-- Created:	Mon Jan 25 18:44:05 1993
-- Author:	Christian CAILLET
--		<cky@sdsun2>
---Copyright:	 Matra Datavision 1993


deferred class ReadWriteModule  from StepData  inherits
    	       ReaderModule     from Interface

    ---Purpose : Defines basic File Access Module (Recognize, Read, Write)
    --           That is : ReaderModule (Recognize & Read) + Write for
    --           StepWriter (for a more centralized description)
    --  Warning : A sub-class of ReadWriteModule, which belongs to a particular
    --           Protocol, must use the same definition for Case Numbers (give
    --           the same Value for a StepType defined as a String from a File
    --           as the Protocol does for the corresponding Entity)

uses Transient,  AsciiString from TCollection,
     SequenceOfAsciiString from TColStd,
     Check, FileReaderData,   StepReaderData,  StepWriter

raises DomainError

is

    CaseNum (me; data : FileReaderData; num : Integer) returns Integer;
    ---Purpose : Translate the Type of record <num> in <data> to a positive
    --           Case Number, or 0 if failed.
    --           Works with a StepReaderData, in which the Type of an Entity
    --           is defined as a String : Reads the RecordType <num> then calls
    --           CaseNum (this type)
    --  Warning : The methods CaseStep, StepType and Recognize,
    --           must be in phase (triplets CaseNum-StepType-Type of Object)

    CaseStep (me; atype : AsciiString from TCollection) returns Integer
        is deferred;
    ---Purpose : Defines Case Numbers corresponding to the recognized Types
    --           Called by CaseNum (data,num) above for a Simple Type Entity
    --  Warning : CaseStep must give the same Value as Protocol does for the
    --           Entity type which corresponds to this Type given as a String

    CaseStep (me; types : SequenceOfAsciiString from TColStd) returns Integer
    	is virtual;
    ---Purpose : Same a above but for a Complex Type Entity ("Plex")
    --           The provided Default recognizes nothing


    IsComplex (me; CN : Integer) returns Boolean  is virtual;
    ---Purpose : Returns True if the Case Number corresponds to a Complex Type
    --           ("Plex"). Remember that all possible combinations must be
    --           aknowledged to be processed
    --           Default is False for all cases. For a Protocol which defines
    --           possible Plexes, this method must be redefined.

    StepType (me; CN : Integer) returns AsciiString from TCollection
        is deferred;
    ---Purpose : Function specific to STEP, which delivers the StepType as it
    --           is recorded in and read from a File compliant with STEP.
    --           This method is symmetric to the method CaseStep.
    --           StepType can be different from Dynamic Type's name, but
    --           belongs to the same class of Object.
    --           Returns an empty String if <CN> is zero.
    --  Warning : For a Complex Type Entity, returns an Empty String
    --           (Complex Type must be managed by users)
    ---C++ : return const &

    ShortType (me; CN : Integer) returns AsciiString from TCollection
    	is virtual;
    ---Purpose : Function specific to STEP. Some STEP Types have a short form
    --           This method can be redefined to fill it
    --           By default, returns an empty string, which is then interpreted
    --           to take normal form from StepType

    ComplexType (me; CN : Integer;
    	    	 types : in out SequenceOfAsciiString from TColStd)
    	returns Boolean  is virtual;
    ---Purpose : Function specific to STEP, which delivers the list of types
    --           which corresponds to a complex type. If <CN> is not for a
    --           complex type, this method returns False. Else it returns True
    --           and fills the list in alphabetic order.
    --           The default returns False. To be redefined as required.

    Read (me; CN : Integer; data : FileReaderData; num : Integer;
    	ach : in out Check; ent : mutable Transient)
    	raises DomainError;
    ---Purpose : General Read Function, calls ReadStep

    ReadStep (me; CN : Integer; data : StepReaderData; num : Integer;
    	ach : in out Check; ent : mutable Transient)
    	raises DomainError  is deferred;
    ---Purpose : Specific Read Function. Works with StepReaderData

    WriteStep (me; CN : Integer; SW : in out StepWriter; ent : Transient)
    	is deferred;
    ---Purpose : Write Function, switched by CaseNum

end ReadWriteModule;
