-- Created on: 1993-03-24
-- Created by: Philippe DAUTRY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Circle from Geom2d inherits Conic from Geom2d

        --- Purpose : Describes a circle in the plane (2D space).
    	-- A circle is defined by its radius and, as with any conic
    	-- curve, is positioned in the plane with a coordinate
    	-- system (gp_Ax22d object) where the origin is the
    	-- center of the circle.
    	-- The coordinate system is the local coordinate
    	-- system of the circle.
    	-- The orientation (direct or indirect) of the local
    	-- coordinate system gives an explicit orientation to the
    	-- circle, determining the direction in which the
    	-- parameter increases along the circle.
    	-- The Geom2d_Circle circle is parameterized by an angle:
    	-- P(U) = O + R*Cos(U)*XDir + R*Sin(U)*YDir
    	-- where:
    	-- - P is the point of parameter U,
    	-- - O, XDir and YDir are respectively the origin, "X
    	--   Direction" and "Y Direction" of its local coordinate system,
    	-- - R is the radius of the circle.
    	-- The "X Axis" of the local coordinate system therefore
 	-- defines the origin of the parameter of the circle. The
    	-- parameter is the angle with this "X Direction".
    	-- A circle is a closed and periodic curve. The period is
    	-- 2.*Pi and the parameter range is [ 0,2.*Pi [.
    	-- See Also
    	-- GCE2d_MakeCircle which provides functions for
    	-- more complex circle constructions
    	-- gp_Ax22d and  gp_Circ2d for an equivalent, non-parameterized data structure.

uses Ax2d     from gp, 
     Ax22d    from gp,
     Circ2d   from gp,
     Pnt2d    from gp,
     Trsf2d   from gp, 
     Vec2d    from gp,
     Geometry from Geom2d


raises ConstructionError from Standard,
       RangeError        from Standard

is


  Create (C : Circ2d)   returns mutable Circle;
	--- Purpose :  Constructs a circle by conversion of the gp_Circ2d circle C.


  Create (A : Ax2d; Radius : Real;
          Sense: Boolean from Standard = Standard_True)  
  returns mutable Circle
        --- Purpose : Constructs a circle of radius Radius, whose center is the origin of axis
    	--   A; A is the "X Axis" of the local coordinate system
    	--   of the circle; this coordinate system is direct if
    	--   Sense is true (default value) or indirect if Sense is false.
    	-- Note: It is possible to create a circle where Radius is equal to 0.0.
    	-- Exceptions Standard_ConstructionError if Radius is negative.
     raises ConstructionError;


  Create (A : Ax22d; Radius : Real)  returns mutable Circle
        --- Purpose : Constructs a circle
	-- of radius Radius, where the coordinate system A
    	--   locates the circle and defines its orientation in the plane such that:
    	--   - the center of the circle is the origin of A,
    	--   - the orientation (direct or indirect) of A gives the
    	--    orientation of the circle.
     raises ConstructionError;


  SetCirc2d (me : mutable; C : Circ2d);
        --- Purpose :
        --  Converts the gp_Circ2d circle C into this circle.

  SetRadius (me : mutable; R : Real)
        --- Warnings : Assigns the value R to the radius of this circle.
    	-- Note: It is possible to have a circle with a radius equal to 0.0.
    	-- Exceptions Standard_ConstructionError if R is negative.
     raises ConstructionError;


  Circ2d (me)   returns Circ2d;
        --- Purpose :
        --  Returns the non persistent circle from gp with the same 
        --  geometric properties as <me>.

  Radius(me) returns Real
  is static;
    	---Purpose: Returns the radius of this circle.
        
  ReversedParameter(me; U : Real) returns Real is redefined static;
  	---Purpose: Computes the parameter on the reversed circle for
    	-- the point of parameter U on this circle.
    	-- For a circle, the returned value is: 2.*Pi - U.


  Eccentricity (me)   returns Real is redefined static;
        --- Purpose :  Returns 0., which is the eccentricity of any circle.


  FirstParameter (me)   returns Real is redefined static;
        --- Purpose : Returns 0.0


  LastParameter (me)   returns Real is redefined static;
        --- Purpose : Returns 2*PI.


  IsClosed (me)   returns Boolean is redefined static;
        --- Purpose : returns True.


  IsPeriodic (me)  returns Boolean is redefined static;
        --- Purpose : returns True. The period of a circle is 2.*Pi.


  D0(me; U : Real; P : out Pnt2d) is redefined static;
	---Purpose: Returns in P the point of parameter U.
        --  P = C + R * Cos (U) * XDir + R * Sin (U) * YDir
        --  where C is the center of the circle , XDir the XDirection and
        --  YDir the YDirection of the circle's local coordinate system.


  D1 (me; U : Real; P : out Pnt2d; V1 : out Vec2d) is redefined static;
        --- Purpose :
        --  Returns the point P of parameter U and the first derivative V1.


  D2 (me; U : Real; P : out Pnt2d; V1, V2 : out Vec2d) is redefined static;
        --- Purpose :
        --  Returns the point P of parameter U, the first and second 
        --  derivatives V1 and V2.


  D3 (me; U : Real; P : out Pnt2d; V1, V2, V3 : out Vec2d) is redefined static;
        --- Purpose :
        --  Returns the point P of parameter u, the first second and third
        --  derivatives V1 V2 and V3.
        

  DN (me; U : Real; N : Integer)   returns Vec2d
        --- Purpose : For the point of parameter U of this circle, computes
    	-- the vector corresponding to the Nth derivative.
    	-- Exceptions: Standard_RangeError if N is less than 1.
            raises RangeError
     is redefined static;



  Transform (me : mutable; T : Trsf2d) is redefined static;
---Purpose: Applies the transformation T to this circle.

       
  Copy (me)  returns mutable like me
     is redefined static;
---Purpose: Creates a new object which is a copy of this circle.
    
fields

  radius : Real;

end;

