-- Created on: 1993-06-14
-- Created by: Martine LANGLOIS
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MakeLine from GeomToStep inherits Root from GeomToStep

    ---Purpose: This class implements the mapping between classes 
    --          Line from Geom and Lin from gp, and the class
    --          Line from StepGeom which describes a line from
    --          Prostep. 
  
uses Lin  from gp,
     Lin2d from gp,
     Line from Geom,
     Line from Geom2d,
     Line from StepGeom
     
raises NotDone from StdFail
     
is 

Create ( L : Lin from gp ) returns MakeLine;

Create ( L : Lin2d from gp ) returns MakeLine;

Create ( C : Line from Geom ) returns MakeLine;

Create ( C : Line from Geom2d ) returns MakeLine;

Value (me) returns Line from StepGeom
    raises NotDone
    is static;
    ---C++: return const&
 
fields

    theLine : Line from StepGeom;
    	-- The solution from StepGeom
    	
end MakeLine;


