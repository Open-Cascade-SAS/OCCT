-- Created on: 1992-08-26
-- Created by: Jean Louis FRENKEL
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


package StdPrs
    	---Purpose: The StdPrs package provides standard display tools
	-- for specific geometries and topologies whereas
	-- Prs3d provides those for generic objects. Among
	-- these classes are definitions of the display of the
	-- specific geometry or topology in various display
	-- modes such as wireframe, shading or hidden line removal mode.
    	       
uses
        Prs3d,
	Geom,
	Geom2d,
	Adaptor3d,
	Adaptor2d,
        GeomAdaptor,
	Geom2dAdaptor,
        BRepAdaptor,
	TopTools,
	TopoDS,
	TopExp,
        TopAbs,
	BRepTools,
	Bnd,
        TColStd,
        HLRAlgo,
    	HLRBRep,
        Quantity,
	BRepMesh,
	gp,
	TColgp,
	Poly,
	TopLoc, 
	Graphic3d

is
   class ToolPoint;
   class ToolVertex;
   class ToolRFace;
   class HLRToolShape;
   --class ToolSectionShape;
   class ToolShadedShape;
   class ShadedShape;
   
   
   class Point 
   instantiates Point from Prs3d(Point from Geom, ToolPoint from StdPrs); 
   
   class Vertex 
   instantiates Point from Prs3d(Vertex from TopoDS, ToolVertex from StdPrs); 
   
   class PoleCurve;
	---Purpose: computes the presentation of curves by drawing
	--          a broken line linking the poles of the curve.

   class Plane;
   	---Purpose: computes the presentation of a infinite plane.

   class WFPoleSurface;
   	---Purpose: computes the presentation of surfaces by drawing a
	--          double network of lines linking the poles of the surface
	--          in the two parametric direction.
	

   class DeflectionCurve;		      
	---Purpose: computes the presentation of objects to be
	--          seen as curves. The computation will be made
	--          according to a maximal chordial deviation.
	          
	---Category: Wireframe algorithms
   
   class WFDeflectionSurface;
	---Purpose: computes the wireframe presentation of surfaces 
	--          by displaying a given number of U and/or V isoparametric
	---         curves. The isoparametric curves are drawn with respect
	--          to a given maximal chordial deviation.

   class ShadedSurface;
   	---Purpose: computes the shading presentation of surfaces.

   -----------------------------------------------
   --- deflection drawing classes :
   -----------------------------------------------

   class WFDeflectionRestrictedFace;


   class WFDeflectionShape instantiates WFShape from Prs3d
	 (WFDeflectionRestrictedFace from StdPrs,
	  DeflectionCurve            from StdPrs,
    	  Vertex                     from StdPrs);
		      
		      
   -----------------------------------------------
   --- Instantiations whith no deflection drawing.
   -----------------------------------------------

   class Curve;
   	---Purpose: computes the presentation of objects to be
	--          seen as curves. The computation will be made
	--          whith a constant number of points.


   class WFSurface;
   	---Purpose: computes the wireframe presentation of surfaces 
	--          by displaying a given number of U and/or V isoparametric
	---         curves. The isoparametric curves are drawn with respect
	--          to a given number of points.


   class WFRestrictedFace instantiates WFRestrictedFace from Prs3d  
    	 (Curve     from StdPrs,
    	  ToolRFace from StdPrs);


   class WFShape instantiates WFShape from Prs3d
	 (WFRestrictedFace  from StdPrs,
	  Curve             from StdPrs,
    	  Vertex            from StdPrs);

    class HLRShape instantiates HLRShape from Prs3d 
    	  (Shape           from TopoDS,
           HLRToolShape    from StdPrs,
	   Curve           from BRepAdaptor,
	   DeflectionCurve from StdPrs);
			
    class HLRPolyShape; 
     
    imported NListOfSequenceOfPnt from Prs3d; 
    imported NListIteratorOfListOfSequenceOfPnt from Prs3d;
    
			
end StdPrs;



