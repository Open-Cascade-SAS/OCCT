-- Created on: 1994-09-05
-- Created by: Gilles DEBARBOUILLE
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class VariableInstance from Dynamic

inherits

    AbstractVariableInstance from Dynamic
    
	---Purpose: This    class  is set   in     the fields of   the
	--          MethodInstance  class.  When   a MethodInstance is
	--          done each  variable of   the definition   must  be
	--          defined in the instance by a VariableInstance with
	--          the same name as in the definition.  If the method
	--          instance is directly  used  by an application  the
	--          user    value    is   directly    set   into   the
	--          VariableInstance. If now the MethodInstance enters
	--          in  the   definition of    a CompositMethod It  is
	--          necessary to define the correspondance between the
	--          variables of the CompositMethod definition and the
	--          use throughout the MethodInstance.

uses

    Variable from Dynamic


is

    Create returns mutable VariableInstance from Dynamic;
    
    ---Level: Public 
    
    ---Purpose: Returns a new empty instance of this class.
    
    Variable(me : mutable ; avariable : Variable from Dynamic)
    
    ---Level: Public 
    
    ---Purpose: Sets    the    variable  <avariable>     into      the
    --          VariableInstance <me>.
    
    is redefined;
    
    Variable(me) returns Variable from Dynamic
    
    ---Level: Public 
    
    ---Purpose: Returns       the      variable contained     into the
    --          VariableInstance <me>.
    
    is static;

fields

    thevariable : Variable from Dynamic;

end VariableInstance;
