-- Created on: 1993-03-23
-- Created by: BBL
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class AidaAlienData from AlienImage inherits AlienImageData from AlienImage

	---Version: 0.0

	---Level: Public
	---Purpose: This class defines an Aida Alien image.


uses
	File 			from OSD,
	ColorImage 		from Image,
	PseudoColorImage 	from Image,
	ColorMap 		from Aspect,
	HArray2OfInteger 	from TColStd,
	DitheringMethod 	from Image,
	Image			from Image

raises
	OutOfRange 	from Standard,
	TypeMismatch 	from Standard

is
	Create returns mutable AidaAlienData from AlienImage ;

	Clear( me : in out mutable ) ;
	---Level: Public
	---Purpose: Frees memory allocated by AidaAlienData
	---C++: alias ~

	Read ( me : in out mutable ; afile : in out File from OSD )
	  returns Boolean from Standard ;
	---Level: Public
	  ---Purpose: Read content of a  AidaAlienData object from a file .
	  --          Returns True if file is a Aida file .

	Write( me : in immutable; afile : in out File from OSD )
	  returns Boolean from Standard ;
	---Level: Public
	  ---Purpose: Write content of a  AidaAlienData object to a file .

	ToImage( me : in  immutable) 
	  returns mutable Image from Image 
          raises TypeMismatch from Standard ;
	  ---Purpose : Converts a AidaAlienData object to a Image object.

	FromImage( me : in out mutable ; anImage : in Image from Image )
          raises TypeMismatch from Standard ;
	  ---Purpose : Converts a Image object to a AidaAlienData object.

	SetColorImageDitheringMethod( me : in out mutable ; 
				      aMethod : DitheringMethod from Image;
				      aColorMap : ColorMap from Aspect ) ;

	---Level: Public
	  ---Purpose: Set the ImageDitheringMethod and the ColorMap when
	  --          FromImage is called with a ColorImage .
	  --	      Aida BYTEMAPS file handle only PseudoColorImage .
	  --          Default value is DM_NearestColor,
	  --		ColorCubeColorMap( 40, 5,1, 8,6, 3,54 )


        AllocData( me : in out mutable ; DX,DY : in Integer from Standard ) 
		is private;
	---Level: Internal
	   ---Purpose : Allocate HArray2 to store Image data

    	Pixel   ( me : in immutable ;     X,Y : in Integer from Standard ) 
			returns Integer from Standard
    			raises OutOfRange from Standard is private ;
	---Level: Internal

    	SetPixel( me : in out mutable; X,Y   : in Integer from Standard ;
			Value : in Integer from Standard )
    			raises OutOfRange from Standard is private ;
	---Level: Internal

	FromPseudoColorImage( me      : in out mutable; 
			      anImage : in PseudoColorImage from Image )
		is private ;
	---Level: Internal
	  ---Purpose : convert a Image object to a AidaAlienData object.

	FromColorImage( me : in out mutable;
			anImage : in ColorImage from Image)
		is private ;
	---Level: Internal
	  ---Purpose : convert a Image object to a AidaAlienData object.

fields
	myDitheringMethod   : DitheringMethod from Image is protected ;

	myDitheringColorMap : ColorMap from Aspect  is protected ;

	myColors : ColorMap from Aspect  is protected ;
	myColorsIsDef : Boolean from Standard  is protected ;

			-- AidaColors definition
	myData	 : HArray2OfInteger from TColStd ;
	myDataIsDef : Boolean from Standard  is protected ;

end ;
 
