-- Created on: 1997-05-21
-- Created by: Christian CAILLET
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DescrProtocol  from StepData    inherits FileProtocol  from StepData

    ---Purpose : A DescrProtocol is a protocol dynamically (at execution time)
    --           defined with :
    --           - a list of resources (inherits FileProtocol)
    --           - a list of entity descriptions
    --           i.e. it can be defined with only C++ writing to initialize it
    --           Its initialization must :
    --           - set its schema name
    --           - define its resources (which can also be other DescrProtocol)
    --           - define its entity descriptions
    --           - record it in the system by calling RecordLib

uses CString, AsciiString from TCollection

is

    Create returns mutable DescrProtocol;

    SetSchemaName (me : mutable; name : CString);
    ---Purpose : Defines a specific Schema Name for this Protocol

    LibRecord     (me);
    ---Purpose : Records this Protocol in the service libraries, with a
    --           DescrGeneral and a DescrReadWrite
    --           Does nothing if the Protocol brings no proper description

    SchemaName (me) returns CString  is redefined;
    ---Purpose : Returns the Schema Name attached to each class of Protocol
    --           here, returns the SchemaName set by SetSchemaName
    -- was C++ : return const

fields

    thename : AsciiString;

end DescrProtocol;
