-- File:	RWStepRepr_RWReprItemAndLengthMeasureWithUnit.cdl
-- Created:	Thu Aug 21 11:55:04 2003
-- Author:	Sergey KUUL
--		<skl@petrox.nnov.matra-dtv.fr>
---Copyright:	 Matra Datavision 2003

class RWReprItemAndLengthMeasureWithUnit from RWStepRepr

	---Purpose : Read & Write Module for ReprItemAndLengthMeasureWithUni

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     ReprItemAndLengthMeasureWithUnit from StepRepr

is

	Create returns RWReprItemAndLengthMeasureWithUnit;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable ReprItemAndLengthMeasureWithUnit from StepRepr);

	WriteStep (me; SW : in out StepWriter; ent : ReprItemAndLengthMeasureWithUnit from StepRepr);

end RWReprItemAndLengthMeasureWithUnit;
