-- Created by: TCL
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class ToleranceFrame from Prs2d inherits Line from Graphic2d

uses

	GraphicObject     from Graphic2d,
	Drawer            from Graphic2d,
	Length	          from Quantity,
	ExtendedString    from TCollection,
	TypeOfTolerance   from Prs2d,
	Tolerance         from Prs2d,
        Array1OfShortReal from TShort,
        FStream           from Aspect,
	Pnt2d             from gp,
	HArray1OfPnt2d    from TColgp
is
	-------------------------
	-- Category: Constructors
	-------------------------

	Create( aGO                   : GraphicObject   from Graphic2d;
        	aX, aY                : Length          from Quantity;
		aHeight               : Length          from Quantity;
            	aTolType              : TypeOfTolerance from Prs2d = Prs2d_TOT_NONE;
            	aTolTxt               : CString         from Standard = "";
		aTxt1                 : CString         from Standard = "";
		aTxt2                 : CString         from Standard = "";
            	anAngle               : Real            from Standard = 0.0;
     	    	aScale                : Real            from Standard = 1.0 );

	---Level: Public
	---Purpose: Creates a frame with a type of tolerance <aTolType>, 
	--          tolerance <aTolTxt>, the reference point is <aXPosition>, <aYPosition
	--          <aX>, <aY> - the center of left vertical edge of this frame
	---Category: Constructor

	--------------------------
	-- Category: Draw and Pick
	--------------------------

	Draw( me : mutable; aDrawer: Drawer from Graphic2d )
    	is static protected;
	---Level: Internal
	---Purpose: Draws the angle <me>.

	Pick( me : mutable; X, Y: ShortReal from Standard;
		  aPrecision: ShortReal from Standard;
		  aDrawer: Drawer from Graphic2d)
	    returns Boolean from Standard
	is static protected;
	---Level: Internal
	---Purpose: Returns Standard_True if the tolerance frame <me> is picked,
	--	    Standard_False if not.
	
	SetHeight( me: mutable; aHSize: Real from Standard );
	---Level: Public
	---Purpose: Defines the height of the frame 

	Height( me ) returns Real from Standard;
	---Level: Public
	---Purpose: Indicates the current height of the frame

 	---------------------------------------------------

	Save( me; aFStream: in out FStream from Aspect ) is virtual;

	ArrayOfPnt2d( me ) returns HArray1OfPnt2d from TColgp;
	---Level: Public
    	---C++: return const
	---Purpose: Returns array of 2d points, which produce frame for tolerance
	--          Size of array == 4

	SetTolText( me: mutable; aText: CString from Standard );
   	---Level: Public
	---Purpose: Sets the text to this tolerance

	SetText1( me: mutable; aText: CString from Standard );
   	---Level: Public

	SetText2( me: mutable; aText: CString from Standard );
   	---Level: Public


	TolText( me ) returns ExtendedString from TCollection;
	---Level: Public
	---Purpose: Returns text and array, which contain points of cell 
        --          which separates the text from other parameters

	Text1( me ) returns ExtendedString from TCollection;
	---Level: Public

	Text2( me ) returns ExtendedString from TCollection;
	---Level: Public

	TextScale( me ) returns Real from Standard;
        ---Level: Public
	

fields

	myX          : ShortReal         from Standard;
    	myY          : ShortReal         from Standard;
    	myTolTxt     : ExtendedString    from TCollection; 
  	myTxt1       : ExtendedString    from TCollection;
	myTxt2       : ExtendedString    from TCollection;
    	myHeight     : ShortReal         from Standard;
    	myAngle      : ShortReal         from Standard;
    	myScale      : ShortReal         from Standard;
	myHTol       : Tolerance         from Prs2d;

  	myXVert      : Array1OfShortReal from TShort;
	myYVert      : Array1OfShortReal from TShort;
	
    
end ToleranceFrame from Prs2d;
