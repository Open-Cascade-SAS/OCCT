-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Block from StepShape 

inherits GeometricRepresentationItem from StepGeom

uses

	Axis2Placement3d from StepGeom, 
	Real from Standard, 
	HAsciiString from TCollection
is

	Create returns mutable Block;
	---Purpose: Returns a Block


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aPosition : mutable Axis2Placement3d from StepGeom;
	      aX : Real from Standard;
	      aY : Real from Standard;
	      aZ : Real from Standard) is virtual;

	-- Specific Methods for Field Data Access --

	SetPosition(me : mutable; aPosition : mutable Axis2Placement3d);
	Position (me) returns mutable Axis2Placement3d;
	SetX(me : mutable; aX : Real);
	X (me) returns Real;
	SetY(me : mutable; aY : Real);
	Y (me) returns Real;
	SetZ(me : mutable; aZ : Real);
	Z (me) returns Real;

fields

	position : Axis2Placement3d from StepGeom;
	x : Real from Standard;
	y : Real from Standard;
	z : Real from Standard;

end Block;
