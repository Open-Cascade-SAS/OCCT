-- Created on: 2008-12-10
-- Created by: Pavel TELKOV
-- Copyright (c) 2008-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MaterialToolDriver from XmlMXCAFDoc  inherits ADriver from XmlMDF

        ---Purpose: Attribute Driver.

uses
    SRelocationTable from XmlObjMgt,
    RRelocationTable from XmlObjMgt,
    Persistent       from XmlObjMgt,
    MessageDriver    from CDM,
    Attribute        from TDF

is
    Create (theMsgDriver:MessageDriver from CDM)
    returns MaterialToolDriver from XmlMXCAFDoc;

    NewEmpty (me)  
    returns Attribute from TDF
    is redefined;

    Paste(me; theSource     : Persistent from XmlObjMgt;
              theTarget     : Attribute from TDF;
              theRelocTable : out RRelocationTable from XmlObjMgt)
    returns Boolean from Standard
    is redefined;

    Paste(me; theSource     : Attribute from TDF;
              theTarget     : in out Persistent from XmlObjMgt;
              theRelocTable : out SRelocationTable from XmlObjMgt)
    is redefined;

end;
