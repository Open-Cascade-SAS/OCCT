-- Created on: 2007-08-17
-- Created by: Sergey ZARITCHNY
-- Copyright (c) 2007-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class HDataMapOfStringByte from TDataStd inherits TShared from MMgt 

	---Purpose: Extension of TDataStd_DataMapOfStringByte class  
    	--          to be manipulated by handle.

uses
    DataMapOfStringByte from TDataStd 
    
is
    Create( NbBuckets: Integer from Standard = 1 )  
    returns mutable HDataMapOfStringByte from TDataStd;    
     
    Create( theOther:  DataMapOfStringByte from TDataStd)  
    returns mutable HDataMapOfStringByte from TDataStd;
     
    Map( me ) returns DataMapOfStringByte from TDataStd
	---C++: return const &
        ---C++: inline      
    is static;	    	
	  
    ChangeMap( me: mutable ) returns DataMapOfStringByte from TDataStd 
    	---C++: return &
        ---C++: inline 
    is static; 	    	
 
fields
    
    myMap : DataMapOfStringByte from TDataStd ;  
   
end HDataMapOfStringByte;
