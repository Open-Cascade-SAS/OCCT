-- Created on: 1993-03-09
-- Created by: Jean-Louis Frenkel
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class HLRToolShape from StdPrs

uses 
    Shape          from TopoDS,
    Curve          from BRepAdaptor,
    Data           from HLRBRep,
    EdgeIterator   from HLRAlgo,
    Projector      from HLRAlgo

is
    Create (TheShape    : Shape     from TopoDS;
            TheProjector: Projector from HLRAlgo) 
    	    returns HLRToolShape from StdPrs;
    NbEdges(me) returns Integer from Standard;
    InitVisible(me: in out; EdgeNumber: Integer from Standard);
    MoreVisible(me) returns Boolean from Standard;
    NextVisible(me: in out);
    Visible(me: in out ; TheEdge : out Curve from BRepAdaptor;
                U1,U2   : out Real from Standard);
    InitHidden(me:in out; EdgeNumber: Integer from Standard);
    MoreHidden(me) returns Boolean from Standard;
    NextHidden(me: in out);
    Hidden(me: in out; TheEdge : out Curve from BRepAdaptor; 
                U1,U2  : out Real from Standard);

fields
    MyData              : Data         from HLRBRep;
    myEdgeIterator      : EdgeIterator from HLRAlgo;
    MyCurrentEdgeNumber : Integer      from Standard;

end HLRToolShape from StdPrs;
