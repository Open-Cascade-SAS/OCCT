-- Created on: 1993-06-23
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class CurvePointInterference from TopOpeBRepDS 
    inherits Interference from TopOpeBRepDS

    ---Purpose: An interference with a parameter.

uses

    Transition  from TopOpeBRepDS,
    Kind        from TopOpeBRepDS,
    OStream     from Standard    
    
is

    Create(T  : Transition from TopOpeBRepDS;
	   ST : Kind from TopOpeBRepDS;
	   S  : Integer from Standard;
	   GT : Kind from TopOpeBRepDS;
	   G  : Integer from Standard;
	   P  : Real from Standard) 
    returns mutable CurvePointInterference from TopOpeBRepDS; 
	    
    Parameter(me) returns Real from Standard
    is static;
    
    Parameter(me : mutable; P : Real from Standard)
    is static;

    Dump(me; OS : in out OStream from Standard) returns OStream
    is redefined;
    ---C++: return &
    
fields

    myParam : Real from Standard;

end CurvePointInterference from TopOpeBRepDS;
