-- Created on: 1993-06-23
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PointData from TopOpeBRepDS
    inherits GeometryData from TopOpeBRepDS

uses

    Point from TopOpeBRepDS

is  

    Create returns PointData;
    Create(P : Point from TopOpeBRepDS) returns PointData;
    Create(P : Point from TopOpeBRepDS; I1,I2 : Integer) returns PointData;
    SetShapes(me:out;I1,I2:Integer);
    GetShapes(me;I1,I2:out Integer);
    
fields 
    
    myPoint : Point from TopOpeBRepDS;
    myS1,myS2 : Integer;
    
friends 

    class DataStructure from TopOpeBRepDS
    
end PointData from TopOpeBRepDS; 
