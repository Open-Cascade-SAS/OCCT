-- Created on: 1993-03-10
-- Created by: JCV
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class Point from Geom inherits Geometry from Geom



    	---Purpose : The abstract class Point describes the common
    	-- behavior of geometric points in 3D space.
    	-- The Geom package also provides the concrete class
    	-- Geom_CartesianPoint.

uses Pnt from gp

is


  Coord (me; X, Y, Z : out Real) 
        ---Purpose : returns the Coordinates of <me>.
     is deferred;


  Pnt (me)  returns Pnt
        ---Purpose : returns a non transient copy of <me>
     is deferred;


  X (me)  returns Real
        ---Purpose : returns the X coordinate of <me>.
     is deferred;


  Y (me)  returns Real
        ---Purpose : returns  the Y coordinate of <me>.
     is deferred;


  Z (me)   returns Real
        ---Purpose : returns the Z coordinate of <me>.
     is deferred;


  Distance (me; Other : Point)  returns Real;
        ---Purpose : Computes the distance between <me> and <Other>.

  
  SquareDistance (me; Other : Point)  returns Real;
        ---Purpose : Computes the square distance between <me> and <Other>.

end;

