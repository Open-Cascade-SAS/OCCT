-- Created on: 1997-10-22
-- Created by: Philippe MANGIN / Sergey SOKOLOV
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class Base from PLib inherits TShared from MMgt 

---Purpose: To work with different polynomial's Bases 

uses 
    Array1OfReal from TColStd
  
is  
    ToCoefficients (me ; Dimension, Degree : Integer;
                    CoeffinBase  : Array1OfReal from TColStd ;
                    Coefficients : out Array1OfReal from TColStd) 
---Purpose:
--   Convert the polynomial P(t) in the canonical base.
    is deferred;

    D0 (me : mutable; U : Real;  
    	BasisValue : out Array1OfReal from TColStd) 
---Purpose: Compute the values of the basis functions in u
--     
    is deferred;
 
    D1 (me : mutable; U : Real;  
      	BasisValue : out Array1OfReal from TColStd; 
     	BasisD1    : out Array1OfReal from TColStd)
---Purpose: Compute the values and the derivatives values of
--          the basis functions in u
    is deferred;
  
    D2 (me : mutable; U : Real;  
    	BasisValue : out Array1OfReal from TColStd; 
	BasisD1    : out Array1OfReal from TColStd; 
    	BasisD2    : out Array1OfReal from TColStd) 
---Purpose: Compute the values and the derivatives values of
--          the basis functions in u
    is deferred;

    D3 (me : mutable; U : Real;  
    	BasisValue : out Array1OfReal from TColStd; 
	BasisD1    : out Array1OfReal from TColStd; 
    	BasisD2    : out Array1OfReal from TColStd; 
        BasisD3    : out Array1OfReal from TColStd)
---Purpose: Compute the values and the derivatives values of
--          the basis functions in u
    is deferred; 

    WorkDegree (me)  returns Integer    
    --- Purpose: returns WorkDegree   
    is  deferred; 

    ReduceDegree ( me ; Dimension ,  MaxDegree  : Integer ;  Tol : Real ; 
                   BaseCoeff :  in  out  Real;
                   NewDegree : out Integer ;
                   MaxError  : out Real)
                            
---Purpose:
--   Compute NewDegree <= MaxDegree so that MaxError is lower
--   than Tol. 
--   MaxError can be greater than Tol if it is not possible
--   to find a NewDegree <= MaxDegree.
--   In this case NewDegree = MaxDegree
-- 

    is  deferred;

end Base;
