-- Created on: 2002-12-12
-- Created by: data exchange team
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class PropertyDefinitionRelationship from StepRepr
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity PropertyDefinitionRelationship

uses
    HAsciiString from TCollection,
    PropertyDefinition from StepRepr

is
    Create returns PropertyDefinitionRelationship from StepRepr;
	---Purpose: Empty constructor

    Init (me: mutable; aName: HAsciiString from TCollection;
                       aDescription: HAsciiString from TCollection;
                       aRelatingPropertyDefinition: PropertyDefinition from StepRepr;
                       aRelatedPropertyDefinition: PropertyDefinition from StepRepr);
	---Purpose: Initialize all fields (own and inherited)

    Name (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Name
    SetName (me: mutable; Name: HAsciiString from TCollection);
	---Purpose: Set field Name

    Description (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Description
    SetDescription (me: mutable; Description: HAsciiString from TCollection);
	---Purpose: Set field Description

    RelatingPropertyDefinition (me) returns PropertyDefinition from StepRepr;
	---Purpose: Returns field RelatingPropertyDefinition
    SetRelatingPropertyDefinition (me: mutable; RelatingPropertyDefinition: PropertyDefinition from StepRepr);
	---Purpose: Set field RelatingPropertyDefinition

    RelatedPropertyDefinition (me) returns PropertyDefinition from StepRepr;
	---Purpose: Returns field RelatedPropertyDefinition
    SetRelatedPropertyDefinition (me: mutable; RelatedPropertyDefinition: PropertyDefinition from StepRepr);
	---Purpose: Set field RelatedPropertyDefinition

fields
    theName: HAsciiString from TCollection;
    theDescription: HAsciiString from TCollection;
    theRelatingPropertyDefinition: PropertyDefinition from StepRepr;
    theRelatedPropertyDefinition: PropertyDefinition from StepRepr;

end PropertyDefinitionRelationship;
