-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class CameraModelD2 from StepVisual 

inherits CameraModel from StepVisual 

uses

	PlanarBox from StepVisual, 
	Boolean from Standard, 
	HAsciiString from TCollection
is

	Create returns CameraModelD2;
	---Purpose: Returns a CameraModelD2


	Init (me : mutable;
	      aName : HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      aName : HAsciiString from TCollection;
	      aViewWindow : PlanarBox from StepVisual;
	      aViewWindowClipping : Boolean from Standard) is virtual;

	-- Specific Methods for Field Data Access --

	SetViewWindow(me : mutable; aViewWindow : PlanarBox);
	ViewWindow (me) returns PlanarBox;
	SetViewWindowClipping(me : mutable; aViewWindowClipping : Boolean);
	ViewWindowClipping (me) returns Boolean;

fields

	viewWindow : PlanarBox from StepVisual;
	viewWindowClipping : Boolean from Standard;

end CameraModelD2;
