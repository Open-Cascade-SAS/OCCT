-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class RightCircularCylinder from StepShape 

inherits GeometricRepresentationItem from StepGeom

uses

	Axis1Placement from StepGeom,
	Real from Standard, 
	HAsciiString from TCollection
is

	Create returns mutable RightCircularCylinder;
	---Purpose: Returns a RightCircularCylinder


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aPosition : mutable Axis1Placement from StepGeom;
	      aHeight : Real from Standard;
	      aRadius : Real from Standard) is virtual;

	-- Specific Methods for Field Data Access --

	SetPosition(me : mutable; aPosition : mutable Axis1Placement);
	Position (me) returns mutable Axis1Placement;
	SetHeight(me : mutable; aHeight : Real);
	Height (me) returns Real;
	SetRadius(me : mutable; aRadius : Real);
	Radius (me) returns Real;

fields

	position : Axis1Placement from StepGeom;
	height : Real from Standard;
	radius : Real from Standard;

end RightCircularCylinder;
