-- Created on: 2002-12-12
-- Created by: data exchange team
-- Copyright (c) 2002-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class CurveElementEndOffset from StepFEA
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity CurveElementEndOffset

uses
    CurveElementEndCoordinateSystem from StepFEA,
    HArray1OfReal from TColStd

is
    Create returns CurveElementEndOffset from StepFEA;
	---Purpose: Empty constructor

    Init (me: mutable; aCoordinateSystem: CurveElementEndCoordinateSystem from StepFEA;
                       aOffsetVector: HArray1OfReal from TColStd);
	---Purpose: Initialize all fields (own and inherited)

    CoordinateSystem (me) returns CurveElementEndCoordinateSystem from StepFEA;
	---Purpose: Returns field CoordinateSystem
    SetCoordinateSystem (me: mutable; CoordinateSystem: CurveElementEndCoordinateSystem from StepFEA);
	---Purpose: Set field CoordinateSystem

    OffsetVector (me) returns HArray1OfReal from TColStd;
	---Purpose: Returns field OffsetVector
    SetOffsetVector (me: mutable; OffsetVector: HArray1OfReal from TColStd);
	---Purpose: Set field OffsetVector

fields
    theCoordinateSystem: CurveElementEndCoordinateSystem from StepFEA;
    theOffsetVector: HArray1OfReal from TColStd;

end CurveElementEndOffset;
