-- File:	StepVisual_ExternallyDefinedCurveFont.cdl
-- Created:	Wed May 10 15:09:07 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class ExternallyDefinedCurveFont from StepVisual
inherits ExternallyDefinedItem from StepBasic

    ---Purpose: Representation of STEP entity ExternallyDefinedCurveFont

uses
    SourceItem from StepBasic,
    ExternalSource from StepBasic

is
    Create returns ExternallyDefinedCurveFont from StepVisual;
	---Purpose: Empty constructor

end ExternallyDefinedCurveFont;
