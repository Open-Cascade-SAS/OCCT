-- Created on: 2005-10-05
-- Created by: Mikhail KLOKOV
-- Copyright (c) 2005-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class SurfaceRangeSample from IntTools
uses
    Range from IntTools,
    CurveRangeSample from IntTools

is
    Create
    	returns SurfaceRangeSample from IntTools;

    Create(theIndexU, theDepthU,theIndexV, theDepthV: Integer from Standard)
    	returns SurfaceRangeSample from IntTools;
	
    Create(theRangeU, theRangeV: CurveRangeSample from IntTools)
    	returns SurfaceRangeSample from IntTools;

    Create(Other: SurfaceRangeSample from IntTools)
    	returns SurfaceRangeSample from IntTools;
    
    Assign(me: in out; Other: SurfaceRangeSample from IntTools)
    	returns SurfaceRangeSample from IntTools;
    	---C++:  alias  operator = 
    	---C++:  return  & 

    SetRanges(me: in out; theRangeU, theRangeV: CurveRangeSample from IntTools);
    	---C++: inline

    GetRanges(me; theRangeU, theRangeV: out CurveRangeSample from IntTools);
	---C++: inline

    SetIndexes(me: in out; theIndexU, theIndexV: Integer from Standard);
	---C++: inline
	
    GetIndexes(me; theIndexU: out Integer from Standard;
    	    	   theIndexV: out Integer from Standard);
	---C++: inline

    GetDepths(me; theDepthU: out Integer from Standard;
    	    	  theDepthV: out Integer from Standard);
	---C++: inline
	
    SetSampleRangeU(me: in out; theRangeSampleU: CurveRangeSample from IntTools);
    	---C++: inline
    
    GetSampleRangeU(me)
    	returns CurveRangeSample from IntTools;
	---C++: return const &
	---C++: inline

    SetSampleRangeV(me: in out; theRangeSampleV: CurveRangeSample from IntTools);
    	---C++: inline
    
    GetSampleRangeV(me)
    	returns CurveRangeSample from IntTools;
	---C++: return const &
	---C++: inline

    SetIndexU(me: in out; theIndexU: Integer from Standard);
    	---C++: inline

    GetIndexU(me)
	returns Integer from Standard;
	---C++: inline

    SetIndexV(me: in out; theIndexV: Integer from Standard);
	---C++: inline
	
    GetIndexV(me)
    	returns Integer from Standard;
	---C++: inline

--
    SetDepthU(me: in out; theDepthU: Integer from Standard);
    	---C++: inline

    GetDepthU(me)
	returns Integer from Standard;
	---C++: inline

    SetDepthV(me: in out; theDepthV: Integer from Standard);
	---C++: inline
	
    GetDepthV(me)
    	returns Integer from Standard;
	---C++: inline


    GetRangeU(me; theFirstU, theLastU: Real from Standard; 
    	    	 theNbSampleU: Integer from Standard)
    	returns Range from IntTools;

    GetRangeV(me; theFirstV, theLastV: Real from Standard; 
    	    	 theNbSampleV: Integer from Standard)
    	returns Range from IntTools;

    IsEqual(me; Other: SurfaceRangeSample from IntTools)
    	returns Boolean from Standard;
	---C++: inline

    GetRangeIndexUDeeper(me; theNbSampleU: Integer from Standard)
    	returns Integer from Standard;
	---C++: inline


    GetRangeIndexVDeeper(me; theNbSampleV: Integer from Standard)
    	returns Integer from Standard;
	---C++: inline

fields
    myRangeU: CurveRangeSample from IntTools;
    myRangeV: CurveRangeSample from IntTools;
    
end SurfaceRangeSample from IntTools;
