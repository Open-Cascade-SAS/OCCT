-- Created on: 2005-01-21
-- Created by: Alexander SOLOVYOV
-- Copyright (c) 2005-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class SensitivePolyhedron from MeshVS inherits SensitiveEntity from Select3D

uses
    EntityOwner                from SelectBasics,
    Projector                  from Select3D,
    Location                   from TopLoc,
    Real                       from Standard,
    Boolean                    from Standard,
    Array1OfPnt2d              from TColgp,
    SequenceOfInteger          from TColStd,
    Box2d                      from Bnd,
    Lin                        from gp,
    ListOfBox2d                from SelectBasics,
    Array1OfPnt                from TColgp,
    HArray1OfPnt               from TColgp,
    HArray1OfPnt2d             from TColgp,
    HArray1OfSequenceOfInteger from MeshVS,
    XY                         from gp

is
    Create( Owner : EntityOwner from SelectBasics;
            Nodes : Array1OfPnt from TColgp;
            Topo  : HArray1OfSequenceOfInteger from MeshVS ) returns mutable SensitivePolyhedron from MeshVS;

    Project( me:mutable; aProjector: Projector from Select3D ) is redefined;

    GetConnected( me:mutable; aLocation: Location from TopLoc ) returns SensitiveEntity from Select3D 
       is redefined;
   
    Matches( me   : mutable; 
             X,Y  : Real from Standard;
             aTol : Real from Standard;
             DMin : out Real from Standard ) returns Boolean is redefined;

    Matches( me                  : mutable; 
             XMin,YMin,XMax,YMax : Real from Standard;
             aTol                : Real from Standard ) returns Boolean from Standard is redefined;

    Matches( me       : mutable; 
             Polyline : Array1OfPnt2d from TColgp;
	     aBox     : Box2d from Bnd;
             aTol     : Real from Standard ) returns Boolean from Standard is redefined;

    GetBox2d( me; aBox : out Box2d from Bnd ) is protected;

    FindIntersection( me; NodesIndices : SequenceOfInteger from TColStd;
                          EyeLine      : Lin from gp ) returns Real is protected;

    ComputeDepth( me; EyeLine: Lin from gp ) returns Real from Standard is redefined;

--  ComputeSize( me ) returns Real from Standard is redefined;

    Areas( me: mutable; aResult : in out ListOfBox2d from SelectBasics ) is redefined;

fields
    myNodes   : HArray1OfPnt from TColgp;
    myNodes2d : HArray1OfPnt2d from TColgp;
    myTopo    : HArray1OfSequenceOfInteger from MeshVS;
    myCenter  : XY from gp;

end SensitiveEntity;

