-- File:	RWStepAP203_RWCcDesignSecurityClassification.cdl
-- Created:	Fri Nov 26 16:26:33 1999 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0
-- Copyright:	Matra Datavision 1999

class RWCcDesignSecurityClassification from RWStepAP203

    ---Purpose: Read & Write tool for CcDesignSecurityClassification

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    CcDesignSecurityClassification from StepAP203

is
    Create returns RWCcDesignSecurityClassification from RWStepAP203;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : CcDesignSecurityClassification from StepAP203);
	---Purpose: Reads CcDesignSecurityClassification

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: CcDesignSecurityClassification from StepAP203);
	---Purpose: Writes CcDesignSecurityClassification

    Share (me; ent : CcDesignSecurityClassification from StepAP203;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWCcDesignSecurityClassification;
