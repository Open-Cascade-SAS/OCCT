-- Created on: 1995-04-25
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



package LocOpe

	---Purpose: Provides  tools to implement local     topological
	--          operations on a shape.

uses MMgt,
     StdFail,
     TCollection,
     TColStd,
     gp, 
     Geom,
     TColGeom,
     TColgp,

     TopAbs,
     TopoDS,
     TopExp,
     TopTools,
     BRepFill,
     BRepAlgo,
     BRepSweep, 
     BOP,
     TopOpeBRepDS
--     TopOpeBRepBuild

is

    class Builder;

    class SplitShape;

    deferred class ProjectedWires;      -- inherits TShared from MMgt
    
    class WiresOnShape;                 -- inherits ProjectedWires from LocOpe


    class Spliter;

    class Generator;

    deferred class GeneratedShape;      -- inherits TShared from MMgt
    
    class GluedShape;                   -- inherits GeneratedShape from LocOpe
    class Prism;
    class Revol;

    class Pipe;

    class DPrism;

    class LinearForm;

    class RevolutionForm;

    class Gluer;

    class FindEdges;

    class FindEdgesInFace;

    class DataMapOfShapePnt instantiates DataMap from TCollection
    	(Shape          from TopoDS,
	 Pnt            from gp,
	 ShapeMapHasher from TopTools);

    class PntFace;
    
    class CurveShapeIntersector;
    
    class CSIntersector;
    

    class BuildShape;

    class SplitDrafts;


    class SequenceOfPntFace instantiates Sequence from TCollection
    	(PntFace from LocOpe);

    class SequenceOfLin instantiates Sequence from TCollection
    	(Lin from gp);

    class SequenceOfCirc instantiates Sequence from TCollection
    	(Circ from gp);

    private class HBuilder;    -- inherits HBuilder from TopOpeBRepBuild

    private class BuildWires;   -- used in LocOpe_Spliter

    enumeration Operation is
    	FUSE,
	CUT,
	INVALID
    end Operation;


    Closed(W: Wire from TopoDS; OnF: Face from TopoDS)
	---Purpose: Returns Standard_True  when the wire <W> is closed
	--          on the face <OnF>.
    	returns Boolean from Standard;
    

    Closed(E: Edge from TopoDS; OnF: Face from TopoDS)
	---Purpose: Returns Standard_True  when the edge <E> is closed
	--          on the face <OnF>.
    	returns Boolean from Standard;

    TgtFaces(E : Edge from TopoDS; 
    	     F1: Face from TopoDS;
    	     F2: Face from TopoDS)
	---Purpose: Returns Standard_True  when the faces are tangent
    	returns Boolean from Standard;


    
--    IsInside(F1: Face from TopoDS; F2: Face from TopoDS)
-- 	---Purpose: Returns Standard_True when  the face F1 is in  the
-- 	--          F2 .
--    	returns Boolean from Standard;
   

    SampleEdges(S : Shape from TopoDS;
    	        Pt: in out SequenceOfPnt from TColgp);


end LocOpe;





