-- Created on: 1994-10-28
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class EdgeVertexInterference from TopOpeBRepDS 
    inherits ShapeShapeInterference from TopOpeBRepDS

    ---Purpose: An interference with a parameter.

uses

    Transition from TopOpeBRepDS,
    Config     from TopOpeBRepDS,
    Kind       from TopOpeBRepDS,    	
    OStream    from Standard    
    
is

    Create(T  : Transition from TopOpeBRepDS;
	   ST : Kind from TopOpeBRepDS;
	   S  : Integer from Standard;
	   G  : Integer from Standard;
      	   GIsBound : Boolean from Standard;
    	   C  : Config from TopOpeBRepDS;
	   P  : Real from Standard)
	   
    returns mutable EdgeVertexInterference from TopOpeBRepDS; 

    	---Purpose: Create an interference of VERTEX <G> on a crossed EDGE E.
    	--  
    	--  if support type <ST> == EDGE : <S> is edge E
    	--                          FACE : <S> is the face with bound E. 
    	--  <T> is the transition along the edge, crossing the crossed edge.
    	--   E  is the crossed edge.
    	--  <GIsBound> indicates if <G> is a bound of the edge.
    	--  <P> is the parameter of <G> on the edge.
    	--  
    	--  interference is stored in the list of interfs of the edge.
    	--  


    Create(T : Transition from TopOpeBRepDS;
	   S : Integer from Standard;
	   G : Integer from Standard;
      	   GIsBound : Boolean from Standard;
    	   C : Config from TopOpeBRepDS;
	   P : Real from Standard) 
	   
    	---Purpose: Create an interference of VERTEX <G> on crossed EDGE <S>.
    	--          
    	--  <T> is the transition along the edge, crossing the crossed edge.
    	--  <S> is the crossed edge.
    	--  <GIsBound> indicates if <G> is a bound of the edge.
    	--  <C> indicates the geometric configuration between
    	--        the edge and the crossed edge.
    	--  <P> is the parameter of <G> on the edge.
    	--  
    	--  interference is stored in the list of interfs of the edge.
    	--  

    returns mutable EdgeVertexInterference from TopOpeBRepDS; 
	    
    Parameter(me) returns Real from Standard
    is static;
    
    Parameter(me : mutable; P : Real from Standard)
    is static;

    Dump(me; OS : in out OStream from Standard) returns OStream
    is redefined;
    ---C++: return &
    
fields

    myParam : Real from Standard;

end EdgeVertexInterference from TopOpeBRepDS;
