-- Created on: 2001-07-09
-- Created by: Julia DOROVSKIKH
-- Copyright (c) 2001-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class ADriver from XmlMDF inherits TShared from MMgt

        ---Purpose: Attribute Storage/Retrieval Driver.

uses
    AsciiString         from TCollection,
    ExtendedString      from TCollection,
    Attribute           from TDF,
    MessageDriver       from CDM,
    RRelocationTable    from XmlObjMgt,
    SRelocationTable    from XmlObjMgt,
    Persistent          from XmlObjMgt,
    Element             from XmlObjMgt

is
    Initialize (theMessageDriver : MessageDriver from CDM;
                theNamespace     : CString from Standard;
                theName          : CString from Standard = NULL);

    VersionNumber(me) returns Integer from Standard
        is virtual;
        ---Purpose: Returns the version number from which the driver
        --          is available.

    NewEmpty    (me)
        returns Attribute from TDF
        is deferred;
        ---Purpose: Creates a new attribute from TDF.

    SourceType  (me) returns Type from Standard;
        ---Purpose: Returns the type of source object,
        --          inheriting from Attribute from TDF.

    TypeName    (me)
        returns AsciiString from TCollection
        is static;
        ---C++: return const &
        ---Purpose: Returns the full XML tag name (including NS prefix)

    Paste       (me; aSource     : Persistent from XmlObjMgt;
                     aTarget     : Attribute from TDF;
                     aRelocTable : out RRelocationTable from XmlObjMgt)
        returns Boolean from Standard
        is deferred;
        ---Purpose: Translate the contents of <aSource> and put it
        --          into <aTarget>, using the relocation table
        --          <aRelocTable> to keep the sharings.

    Paste       (me; aSource     : Attribute from TDF;
                     aTarget     : in out Persistent from XmlObjMgt;
                     aRelocTable : out SRelocationTable from XmlObjMgt)
        is deferred;
        ---Purpose: Translate the contents of <aSource> and put it
        --          into <aTarget>, using the relocation table
        --          <aRelocTable> to keep the sharings.

    WriteMessage (me; theMessage : ExtendedString from TCollection);
        ---Purpose: Send message to Application (usually when error occurres)

fields

    myMessageDriver : MessageDriver from CDM;
    myTypeName      : AsciiString from TCollection is protected;

end ADriver;
