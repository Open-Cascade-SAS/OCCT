-- Created on: 1998-02-04
-- Created by: Christian CAILLET
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class SignType  from Interface    inherits SignText from MoniTool

    	---Purpose : Provides the basic service to get a type name, according
    	--           to a norm
    	--           It can be used for other classes (general signatures ...)

uses CString, Transient, AsciiString, InterfaceModel

is

--    Name (me) returns CString  is deferred;  already in SignText
    ---Purpose : Returns an identification of the Signature (a word), given at
    --           initialization time

    Text  (me; ent : any Transient; context : any Transient)
    	returns AsciiString from TCollection;
    ---Purpose : Specialised to consider context as an InterfaceModel


    Value (me; ent : any Transient; model : InterfaceModel)
    	returns CString  is deferred;
    ---Purpose : Returns the Signature for a Transient object. It is specific
    --           of each sub-class of Signature. For a Null Handle, it should
    --           provide ""
    --           It can work with the model which contains the entity

    ClassName (myclass; typnam : CString) returns CString;
    ---Purpose : From a CDL Type Name, returns the Class part (package dropped)
    --           WARNING : buffered, to be immediately copied or printed

end SignType;
