-- Created on: 1995-12-07
-- Created by: FMA
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class GeometricRepresentationContextAndParametricRepresentationContext from StepGeom 

inherits RepresentationContext from StepRepr


	--- This classe is an implementation of EXPRESS
	--  ANDOR Subtype Declaration.
	--  
	--  Hand made by FMA - 1995 Feb 9th
uses

	GeometricRepresentationContext from StepGeom, 
	ParametricRepresentationContext from StepRepr, 
	HAsciiString from TCollection, 
	Integer from Standard

is

	Create returns GeometricRepresentationContextAndParametricRepresentationContext;
	---Purpose: empty constructor


	Init (me : mutable;
	      aContextIdentifier : HAsciiString from TCollection;
	      aContextType : HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      aContextIdentifier : HAsciiString from TCollection;
	      aContextType : HAsciiString from TCollection;
	      aGeometricRepresentationContext : GeometricRepresentationContext from StepGeom;
	      aParametricRepresentationContext : ParametricRepresentationContext from StepRepr) is virtual;

	Init (me : mutable;
	      aContextIdentifier : HAsciiString from TCollection;
	      aContextType : HAsciiString from TCollection;
	      aCoordinateSpaceDimension : Integer from Standard) is virtual;

	-- Specific Methods for Field Data Access --

	SetGeometricRepresentationContext(me : mutable; aGeometricRepresentationContext : GeometricRepresentationContext);
	GeometricRepresentationContext (me) returns GeometricRepresentationContext;
	SetParametricRepresentationContext(me : mutable; aParametricRepresentationContext : ParametricRepresentationContext);
	ParametricRepresentationContext (me) returns ParametricRepresentationContext;

	-- Specific Methods for ANDOR Field Data Access --

	SetCoordinateSpaceDimension(me : mutable; aCoordinateSpaceDimension : Integer);
	CoordinateSpaceDimension (me) returns Integer;


fields

	geometricRepresentationContext : GeometricRepresentationContext from StepGeom;
	parametricRepresentationContext : ParametricRepresentationContext from StepRepr;

end GeometricRepresentationContextAndParametricRepresentationContext;
