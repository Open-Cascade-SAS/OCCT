-- File:	STEPSelections_AssemblyExplorer.cdl
-- Created:	Wed Mar 24 15:12:12 1999
-- Author:	data exchange team
--		<det@friendox.nnov.matra-dtv.fr>
---Copyright:	 Matra Datavision 1999


class AssemblyExplorer from STEPSelections 

	---Purpose: 

uses
    
    Graph from Interface,
    SequenceOfAssemblyComponent        from STEPSelections,
    IndexedDataMapOfTransientTransient from TColStd,
    ProductDefinition                  from StepBasic,
    ShapeDefinitionRepresentation      from StepShape,
    AssemblyComponent                  from STEPSelections,
    NextAssemblyUsageOccurrence        from StepRepr
    
is
    
    Create (G: Graph) returns AssemblyExplorer from STEPSelections;
    
    Init(me: in out; G: Graph);
    
    Dump(me; os: in out OStream from Standard);
    
    FindSDRWithProduct(me; product: ProductDefinition from StepBasic)
    returns ShapeDefinitionRepresentation from StepShape;
    
    FillListWithGraph(me: in out; cmp: AssemblyComponent from STEPSelections);
    
    FindItemWithNAUO(me; nauo: NextAssemblyUsageOccurrence from StepRepr)
    returns Transient from Standard;
    
    --Methods for fetching the results
    
    NbAssemblies(me) returns Integer;
    	---Purpose: Returns the number of root assemblies;
	---C++: inline
    
    Root(me; rank: Integer = 1) returns AssemblyComponent from STEPSelections;
    	---Purpose: Returns root of assenbly by its rank;
	---C++: inline
    

fields

    myRoots: SequenceOfAssemblyComponent from STEPSelections;
    myGraph: Graph from Interface;
    myMap  : IndexedDataMapOfTransientTransient from TColStd;    

end AssemblyExplorer;
