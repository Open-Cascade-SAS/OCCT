-- Created on: 1995-10-24
-- Created by: Mister rmi
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PolygonOnClosedTriangulation from PBRep 
    
    inherits PolygonOnTriangulation  from  PBRep


    	---Purpose: A representation by two arrays of nodes on a 
    	--          triangulation.


uses PolygonOnTriangulation from PPoly,
     Location               from PTopLoc,
     Triangulation          from PPoly


is

    Create(P1, P2   : PolygonOnTriangulation from PPoly;
    	   S        : Triangulation    from PPoly;
	   L        : Location         from PTopLoc)
    returns PolygonOnClosedTriangulation from PBRep;


    IsPolygonOnClosedTriangulation(me)    returns Boolean
    	---Purpose: Returns True.
    is redefined;

    PolygonOnTriangulation2(me) 
    returns any PolygonOnTriangulation from PPoly;

fields

    myPolygon2:  PolygonOnTriangulation from PPoly;

end PolygonOnClosedTriangulation;
