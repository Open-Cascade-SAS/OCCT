-- Created on: 1995-02-23
-- Created by: Mister rmi
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class ViewerSelector2d from StdSelect inherits ViewerSelector from SelectMgr

	---Purpose: A viewer selection framework.
    	-- The objects defined in this framework can be passed to a selection manager.
        
uses

    View          from V2d,
    Projector     from Select2D,
    Selection     from SelectMgr,
    GraphicObject from Graphic2d

is

    Create returns mutable ViewerSelector2d from StdSelect;

    	--- Purpose: Constructs an empty viewer selection framework.
    
    Create (aProjector: Projector from Select2D) 
    returns mutable ViewerSelector2d from StdSelect;
    	---Purpose: Constructs the viewer selection framework defined by
    	-- the projector aProjector.
    
    Set(me:mutable; aSensitivity : Integer) is static;
    	---Level: Public 
    	---Purpose: Sets a pixel tolerance for the selection.
    	--         will be converted for picking in a view.


    Set(me:mutable; aProjector: Projector from Select2D) is static;
    	---Purpose: Sets the new projector aProjector.   

    Convert(me:mutable;aSelection:mutable Selection from SelectMgr) 
    is redefined static;

    Pick (me           : mutable;XPix,YPix:Integer;
    	  aView        : View from V2d) is static;
    	---Purpose: Returns the pixel coordinates of the mouse Xpix, Ypix
    	-- in the view aView. 

    Pick (me:mutable;XPMin,YPMin,XPMax,YPMax:Integer;aView:View from V2d) is static;
    	---Purpose: Returns the minimum and maximum pixel coordinates
    	-- XPMin, YPMin and XPMax, YPMax defining a 2D area in the view aView.



    Projector (me) returns any Projector from Select2D;
    	---Purpose: Returns the projector which defines this framework.
    	---C++: inline

    	
    DisplayAreas (me:mutable;aView:View from V2d) is static;
    	---Purpose: Displays the active areas in the given view;



    ClearAreas(me:mutable) is static;    
    	---Purpose: Clear the displayed sensitive areas from this framework..
	


fields

    myprj    : Projector from Select2D;
    mypixtol : Integer;
    
    mygo     : GraphicObject from Graphic2d;
    
end ViewerSelector2d;


