-- Created on: 1993-06-17
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package TopOpeBRep 

	---Purpose: This package provides  the topological  operations
	--          on the BRep data structure.

uses

    Standard,
    MMgt,
    TColStd,
    TopAbs,
    TopoDS,
    TopTools,
    TopExp,
    gp,
    Geom,
    Geom2d,
    GeomAbs,
    Geom2dAdaptor,
    Bnd,
    BRep,
    BRepClass,
    BRepAdaptor,
    BRepTopAdaptor,
    ProjLib,
    IntRes2d,
    Geom2dInt,    
    
    IntSurf,
    IntPatch,

    GeomAdaptor,
    IntCurveSurface,
    BRepIntCurveSurface,

    TopOpeBRepDS,
    TopOpeBRepTool,
    TCollection
    
is

    enumeration TypeLineCurve is
    	ANALYTIC,RESTRICTION,WALKING,
        LINE,CIRCLE,ELLIPSE,PARABOLA,HYPERBOLA,
	OTHERTYPE
    end TypeLineCurve;

    class VPointInter;

    imported Array1OfVPointInter;

    imported transient class HArray1OfVPointInter;

    pointer PThePointOfIntersection to Point from IntPatch;
    class VPointInterIterator;

    pointer PPntOn2S to PntOn2S from IntSurf;
    class WPointInter;
    
    class WPointInterIterator;
	 
    class LineInter;
    pointer PLineInter to LineInter from TopOpeBRep;
	
    imported Array1OfLineInter;

    imported transient class HArray1OfLineInter;

    imported DataMapOfTopolTool;

    imported DataMapIteratorOfDataMapOfTopolTool;

    pointer PIntRes2d_IntersectionPoint to IntersectionPoint from IntRes2d;
    class Hctxff2d;
    class Hctxee2d;

    enumeration P2Dstatus is
    	P2DUNK,P2DINT,P2DSGF,P2DSGL,P2DNEW 
    end P2Dstatus;
    
    class Point2d;
    imported SequenceOfPoint2d;
    
    class PointClassifier;

    class VPointInterClassifier;

    class GeomTool;
     
    class FacesIntersector;

    pointer PFacesIntersector to FacesIntersector from TopOpeBRep;
	
    class EdgesIntersector;

    pointer PEdgesIntersector to EdgesIntersector from TopOpeBRep;

    class FaceEdgeIntersector;

    class ShapeScanner;

    class ShapeIntersector;

    class ShapeIntersector2d;

    class PointGeomTool;
    
    class FFTransitionTool;

    class Bipoint;
    imported ListOfBipoint;
    imported ListIteratorOfListOfBipoint;
    
    class FacesFiller;
    pointer PFacesFiller to FacesFiller from TopOpeBRep;
    class FFDumper;

    class EdgesFiller;

    class FaceEdgeFiller;

    class DSFiller;

    Print(TLC  : TypeLineCurve from TopOpeBRep; OS  : in out OStream) 
    ---C++: return &
    returns OStream;
    ---Purpose: Prints the name  of  <TLC>  as  a String  on the
    --          Stream <S> and returns <S>.

end TopOpeBRep;
