-- Created on: 1991-06-27
-- Created by: Remi LEQUETTE
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



package BRep 

	---Purpose: This package describes  a Boundary  Representation
	--          Data   Structure   inherited  from   the  abstract
	--          Topology   defined  in the   TopoDS  package.  The
	--          geometric data are provided by the Geom and Geom2d
	--          packages.
	--          
	--          The TVertex,  TEdge,  and TFace  are  redefined in
	--          this package to add geometric information.

        ---Level : Public  
        --  All methods of all  classes will be public.

uses
    MMgt,        -- Memory management
    TCollection, -- Basic data structures
    TColStd,     -- HArray1OfInteger
    gp,          -- Elementary geometry
    Bnd,         -- Bounding boxes
    TopLoc,      -- Local coordinate systems
    TopAbs,      -- Enumerations : Orientation, ShapeType
    TopoDS,      -- Abstract topological data structure
    GeomAbs,     -- Enumerations : Shape
    Geom,        -- 3D geometry : curves and surfaces
    Geom2d,      -- 2D geometry : curves in parametric space
    Poly         -- Triangulations and Polygons

is

    --
    --  Face
    --  

    class TFace;
	---Purpose: The TFace  class is inherited  from the TFace from
	--          TopoDS. It contains a  surface, a tolerance  and a
	--          natural restriction flag.
	
    --
    --  Edge
    --
    --  An Edge is  defined by a list  of curve representations  which
    --  are either :
    --  
    --  Geometric representations :
    --  
    --  * A 3d curve (at most one)
    --  
    --  * A curve on surface, curve in parametric space.
    --  
    --  * A curve on closed surface, two curves in parametric space.
    --  
    --  Polygonal representations :
    --  
    --  * A 3d polygon (at most one).
    --  
    --  * A Polygon on triangulation (array of node indices)
    --  
    --  * A Polygon on closed triangulation (2 arrays of node indices)
    --  
    --  * A polygon on surface (array of 2d points in parametric space)
    --  
    --  Curve on 2 surfaces :
    --  
    --  * This is used for storing shape continuity.
    --  

    deferred class CurveRepresentation;
	---Purpose: Root      for curve representations.    Contains a
	--          location.

    class ListOfCurveRepresentation instantiates
    List from TCollection (CurveRepresentation from BRep);
    
    deferred class GCurve;
	---Purpose: Root class  for geometric curves  representations.
	--          Contains a first an a last parameter.

    class Curve3D;
	---Purpose: Representation by a 3d curve.

    class CurveOnSurface;
	---Purpose: Representation by a curve in the  parametric space
	--          of a surface.

    class CurveOnClosedSurface;
	---Purpose: Representation  by two   curves in the  parametric
	--          space of a closed surface.

    class Polygon3D;
	---Purpose: Representation by a 3D polygon.

    class PolygonOnTriangulation;
	---Purpose: Representation by    an array  of  indices  on   a
	--          triangulation.
	
    class PolygonOnClosedTriangulation;
	---Purpose: Representation   by two  arrays  of indices   on a
	--          triangulation.
	
    class PolygonOnSurface;
	---Purpose: Representation by 2d polygon in the parametric space
	--          of a surface.

    class PolygonOnClosedSurface;
	---Purpose: Representation by two 2d polygons in the parametric
	--          space of the  surface.
	
    class CurveOn2Surfaces;
	---Purpose: Geometric continuity bewtween two surfaces.

    class TEdge;
	---Purpose: The TEdge class is  inherited  from the TEdge from
	--          TopoDS.   It contains a  3d   curve and  a list of
	--          representations.

	
    --
    --  Vertex
    --

    deferred class PointRepresentation;
	---Purpose: Root  for   point   representations.  Contains   a
	--          location. 
	
    class ListOfPointRepresentation instantiates
    List from TCollection (PointRepresentation from BRep);
    
    class PointOnCurve;
	---Purpose: Representation by a parameter on a 3D curve.
	
    deferred class PointsOnSurface;
	---Purpose: Root for points on surface.
    
    class PointOnCurveOnSurface;
	---Purpose: Representation by   a parameter on  a curve   on a
	--          surface. 

    class PointOnSurface;
	---Purpose: Representation by two parameters on a surface.

    class TVertex;
	---Purpose: The TVertex class  is  inherited from the  TVertex
	--          from    TopoDS.  It contains  a  3d  point   and a
	--          location.

    class Builder;
	---Purpose: The  Builder  from BRep is   inherited    from the
	--          Builder3D   from  TopoDS.    It  is  used to build
	--          Shapes.

    class Tool;
	---Purpose: The Tool from BRep is used to access the geometric
	--          data.


end BRep;
