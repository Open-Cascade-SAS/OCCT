-- Created on: 1993-11-08
-- Created by: Laurent BUCHARD
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



generic class WLine from ApproxInt ( 
    TheCurve        as any;
    TheCurveTool    as any;
    TheCurve2d      as any;
    TheCurveTool2d  as any)
    
    inherits TShared from MMgt
    
   
uses PntOn2S           from IntSurf,
     LineOn2S          from IntSurf
     
is 
     
     Create(CurveXYZ: TheCurve;
            CurveUV1: TheCurve2d;
	    CurveUV2: TheCurve2d)
	
	 returns mutable WLine from ApproxInt;

     Create(lin: LineOn2S from IntSurf;  Tang: Boolean from Standard)
     
	 returns mutable WLine from ApproxInt;
	 
     NbPnts(me) 
     
         returns Integer from Standard
	 is static;
	 
     Point(me: mutable; Index: Integer from Standard)
     
         returns PntOn2S from IntSurf
	 is static;
	 
fields 

    curvxyz  : TheCurve;
    curvuv1  : TheCurve2d;
    curvuv2  : TheCurve2d;
    pnton2s  : PntOn2S    from IntSurf;
    linon2s  : LineOn2S   from IntSurf;
end WLine;

