-- Created on: 2009-04-06
-- Created by: Sergey ZARITCHNY
-- Copyright (c) 2009-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Point from TDataXtd inherits Attribute from TDF

	---Purpose: 
    	-- The basis to define a point attribute.
    	-- The topological attribute must contain a vertex.
    	-- You use this class to create reference points in a design.
	--          
	--  Warning:  Use TDataXtd_Geometry  attribute  to retrieve the
	--          gp_Pnt of the Point attribute

uses Attribute       from TDF,
     Label           from TDF,
     GUID            from Standard,
     Pnt             from gp,
     DataSet         from TDF,
     RelocationTable from TDF

is    


    ---Purpose: class methods
    --          =============
      
    GetID(myclass)    
    	---C++: return const & 
    returns GUID from Standard;   
    	---Purpose:
    	-- Returns the GUID for point attributes.

    Set (myclass ; label : Label from TDF) 
    	---Purpose: 
    	-- Sets the label Label as a point attribute.
    	-- If no object is found, a point attribute is created.
    returns Point from TDataXtd;      

    Set (myclass ; label : Label from TDF; P : Pnt from gp)
    	---Purpose: 
    	-- Sets the label Label as a point attribute containing the point P.
    	-- If no object is found, a point attribute is created.
    returns Point from TDataXtd;    

    ---Purpose: Point methods
    --          =============    

    Create
    returns mutable Point from TDataXtd;  

    ---Category: TDF_Attribute methods
    --           =====================

    
    ID (me)  
    	---C++: return const & 
    returns GUID from Standard;

    Restore (me: mutable; With : Attribute from TDF);

    NewEmpty (me)
    returns mutable Attribute from TDF;

    Paste (me; Into : mutable Attribute from TDF;
	       RT   : mutable RelocationTable from TDF);  

    Dump (me; anOS : in out OStream from Standard) 
    	returns OStream from Standard
    	is redefined;
	---C++: return &

end Point;

