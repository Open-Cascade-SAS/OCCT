-- Created on: 1993-01-29
-- Created by: Isabelle GRIGNON
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PolyLine from IntPatch

inherits Polygo from IntPatch

uses Pnt2d from gp,
     Box2d from Bnd,
     IType from IntPatch,
     WLine from IntPatch,
     RLine from IntPatch

is

    Create
    returns PolyLine from IntPatch;

    Create (InitDefle: Real from Standard)
   	returns PolyLine from IntPatch;

    SetWLine(me: in out; OnFirst: Boolean from Standard; Line: WLine from IntPatch)
    	is static;

    SetRLine(me: in out; OnFirst: Boolean from Standard; Line: RLine from IntPatch)
      	is static;

    Prepare(me: in out)
      	is static private;

    ResetError(me: in out);

    NbPoints(me) returns Integer;
  
    Point(me; Index : Integer) 
    	returns Pnt2d from gp;
                                      	    	 

fields

    pnt      : Pnt2d   from gp;
    typ      : IType   from IntPatch;
    onfirst  : Boolean from Standard;
    wpoly    : WLine from IntPatch;
    rpoly    : RLine from IntPatch;

end PolyLine;
