-- Created on: 1993-01-28
-- Created by: Gilles DEBARBOUILLE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class Parameter from Dynamic 
inherits

    TShared from MMgt


	---Purpose: A  parameter is defined  as  the association of  a
	--          name and a value.  For easy use, inherited classes
	--          have been  created  to manipulate  values by their
	--          C++ type.  This class is the root class of all the
	--          derived parameter classes.  Only the identifier of
	--          the parameter is  stored  in it.   The  associated
	--          value is stored in the  inherited classes where it
	--          is more  easy to overload the methods manipulating
	--          the  value.   No  instance of  this class  must be
	--          created. It is for this  reason that this class is
	--          deferred.

uses

    OStream from Standard,
    CString from Standard,
    HAsciiString from TCollection,
    AsciiString  from TCollection


is

    Initialize(aname : CString from Standard) ;
    
    ---Level: Internal 
    
    ---Purpose: Initializer of this class  taking in argument the name
    --          of the parameter <aname>.
    
    Name(me) returns AsciiString from TCollection
    
    ---Level: Public 

    ---Purpose: Returns in an AsciiString the name of the parameter.

    is static;
        
    Dump(me ; astream : in out OStream from Standard)
    
    ---Level: Internal 
    
    ---Purpose: Useful for debugging.
    
    is virtual;
    
fields

    theparametername : HAsciiString from TCollection;
    
end Parameter;
