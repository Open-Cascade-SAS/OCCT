-- Created on: 1993-03-10
-- Created by: JCV
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class CylindricalSurface from Geom inherits ElementarySurface from Geom

       
        ---Purpose : This class defines the infinite cylindrical surface.
        --  
        --  The local coordinate system of the CylindricalSurface is defined
        --  with an axis placement (see class ElementarySurface).
        --  
        --  The "ZAxis" is the symmetry axis of the CylindricalSurface, 
        --  it gives the direction of increasing parametric value V.
        --  
        --  The parametrization range is :
        --       U [0, 2*PI],  V ]- infinite, + infinite[
        --       
        --  The "XAxis" and the "YAxis" define the placement plane of the 
        --  surface (Z = 0, and parametric value V = 0)  perpendicular to 
        --  the symmetry axis. The "XAxis" defines the origin of the 
        --  parameter U = 0.  The trigonometric sense gives the positive 
        --  orientation for the parameter U.
        -- 
        --  When you create a CylindricalSurface the U and V directions of
        --  parametrization are such that at each point of the surface the
        --  normal is oriented towards the "outside region".
        -- 
        --  The methods UReverse VReverse change the orientation of the 
        --  surface.

uses Ax3      from gp, 
     Cylinder from gp,
     Pnt      from gp, 
     Trsf     from gp,
     GTrsf2d  from gp,
     Vec      from gp,
     Curve    from Geom, 
     Geometry from Geom

raises ConstructionError from Standard,
       RangeError        from Standard


is

  Create (A3 : Ax3; Radius : Real)    returns mutable CylindricalSurface
        ---Purpose :
        --  A3 defines the local coordinate system of the cylindrical surface.
        --  The "ZDirection" of A3 defines the direction of the surface's
        --  axis of symmetry.
        --  At the creation the parametrization of the surface is defined
        --  such that the normal Vector (N = D1U ^ D1V) is oriented towards
        --  the "outside region" of the surface.
        --- Warnings :
        --  It is not forbidden to create a cylindrical surface with 
        --  Radius = 0.0
     raises ConstructionError;
        ---Purpose : Raised if Radius < 0.0



  Create (C : Cylinder)  returns mutable CylindricalSurface;
        ---Purpose :
        --  Creates a CylindricalSurface from a non transient Cylinder
        --  from package gp.



  SetCylinder (me : mutable; C : Cylinder);
        ---Purpose :
        --  Set <me> so that <me> has the same geometric properties as C.


  SetRadius (me : mutable; R : Real)
        ---Purpose : Changes the radius of the cylinder.
     raises ConstructionError;
        ---Purpose : Raised if R < 0.0


  Cylinder (me)   returns Cylinder;
        ---Purpose :
        --  returns a non transient cylinder with the same geometric 
        --  properties as <me>.


  UReversedParameter (me; U : Real) returns Real;
	---Purpose: Return the  parameter on the  Ureversed surface for
	--          the point of parameter U on <me>.
	--          Return 2.PI - U.


  VReversedParameter (me; V : Real) returns Real;
	---Purpose: Return the  parameter on the  Vreversed surface for
	--          the point of parameter V on <me>.
	--          Return -V

  TransformParameters(me; U,V : in out Real; T : Trsf from gp)
	---Purpose: Computes the  parameters on the  transformed  surface for
	-- the transform of the point of parameters U,V on <me>.
	--          me->Transformed(T)->Value(U',V')
	--          is the same point as
	--          me->Value(U,V).Transformed(T)
	--   Where U',V' are the new values of U,V after calling
	--          me->TranformParameters(U,V,T)
	--          This methods multiplies V by T.ScaleFactor()
     is redefined;  

  ParametricTransformation(me; T : Trsf from gp) returns GTrsf2d from gp
    	---Purpose: Returns a 2d transformation  used to find the  new
    	--          parameters of a point on the transformed surface.
	--          me->Transformed(T)->Value(U',V')
	--          is the same point as
	--          me->Value(U,V).Transformed(T)
	--  Where U',V' are  obtained by transforming U,V with
	--          th 2d transformation returned by
	--          me->ParametricTransformation(T)
	--    This  methods  returns  a scale  centered  on  the
	--          U axis with T.ScaleFactor
     is redefined;  



  Bounds (me; U1, U2, V1, V2 : out Real);
        ---Purpose :
        --  The CylindricalSurface is infinite in the V direction so
        --  V1 = Realfirst, V2 = RealLast from package Standard.
        --  U1 = 0 and U2 = 2*PI.


  Coefficients (me; A1, A2, A3, B1, B2, B3, C1, C2, C3, D : out Real);
       	---Purpose :
       	--  Returns the coefficients of the implicit equation of the quadric
       	--  in the absolute cartesian coordinate system :
       	--  These coefficients are normalized.
       	--  A1.X**2 + A2.Y**2 + A3.Z**2 + 2.(B1.X.Y + B2.X.Z + B3.Y.Z) +
       	--  2.(C1.X + C2.Y + C3.Z) + D = 0.0


  Radius (me)   returns Real;
    	---Purpose: Returns the radius of this cylinder.

  IsUClosed (me)  returns Boolean;
        ---Purpose : Returns True.


  IsVClosed (me)  returns Boolean;
        ---Purpose : Returns False.


  IsUPeriodic (me)  returns Boolean;
        ---Purpose : Returns True.


  IsVPeriodic (me)  returns Boolean;
        ---Purpose : Returns False.


  UIso (me; U : Real)  returns mutable Curve;
        ---Purpose :
        --  The UIso curve is a Line. The location point of this line is
        --  on the placement plane (XAxis, YAxis) of the surface.
        --  This line is parallel to the axis of symmetry of the surface.


  VIso (me; V : Real)   returns mutable Curve;
        ---Purpose :
        --  The VIso curve is a circle. The start point of this circle 
        --  (U = 0) is defined with the "XAxis" of the surface.
        --  The center of the circle is on the symmetry axis.


  D0 (me; U, V : Real; P : out Pnt);
        ---Purpose :
        --  Computes the  point P (U, V) on the surface.
        --  P (U, V) = Loc + Radius * (cos (U) * XDir + sin (U) * YDir) + 
        --             V * ZDir
        --  where Loc is the origin of the placement plane (XAxis, YAxis)
        --  XDir is the direction of the XAxis and YDir the direction of
        --  the YAxis.


  D1 (me; U, V : Real; P : out Pnt; D1U, D1V : out Vec);
        ---Purpose :
        --  Computes the current point and the first derivatives in the
        --  directions U and V.


  D2 (me; U, V : Real; P : out Pnt; D1U, D1V, D2U, D2V, D2UV : out Vec);
        ---Purpose :
        --  Computes the current point, the first and the second derivatives
        --  in the directions U and V.


  D3 (me; U, V : Real; P : out Pnt; 
      D1U, D1V, D2U, D2V, D2UV, D3U, D3V, D3UUV, D3UVV : out Vec);
        ---Purpose :
        --  Computes the current point, the first, the second and the 
        --  third   derivatives in the directions U and V.


  DN (me; U, V : Real; Nu, Nv : Integer)   returns Vec
        ---Purpose :
        --  Computes the derivative of order Nu in the direction u and Nv
        --  in the direction v.
     raises RangeError;
        ---Purpose : Raised if Nu + Nv < 1 or Nu < 0 or Nv < 0.



  Transform (me : mutable; T : Trsf);
    	---Purpose:  Applies the transformation T to this cylinder.
  Copy (me)  returns mutable like me;
    	---Purpose:  Creates a new object which is a copy of this cylinder.
fields

  radius : Real;
        
end;
