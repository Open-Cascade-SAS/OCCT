-- Created on: 1996-07-26
-- Created by: Maria PUMBORIOS
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package FilletSurf 

	---Purpose:  This package contains the API giving 
	--           only geometric informations about fillets
	--           for Toyota Project UV4. 
        
uses
    TopoDS,
    TopTools,
    ChFi3d,
    ChFiDS,
    BRepAdaptor,
    Adaptor3d,
    math,
    Geom,
    Geom2d,
    gp,
    StdFail,
    TopAbs
is

---------------------------------------------------------- 
--  enumeration used to describe the status of start and end section
--  of the fillet 
--   TwoExtremityOnEdge
--   OneExtremityOnEdge
--   NoExtremityOnEdge
----------------------------------------------------------
--                                                               
--    
enumeration StatusType  is  TwoExtremityOnEdge, OneExtremityOnEdge, 
                            NoExtremityOnEdge  
end  StatusType;
    
---------------------------------------------------------- 
--  enumeration used to describe the status of the computation of the fillet
-- IsOk  
-- IsNotOk 
-- IsPartial    
--   
----------------------------------------------------------

enumeration StatusDone  is  IsOk, IsNotOk,IsPartial 
                      
end  StatusDone;

---------------------------------------------------------- 
--  enumeration used to describe the  status error  
--   EmptyList 
--   EdgeNotG1 
--   FacesNotG1
--    EdgeNotOnShape    
--    NotSharpEdge
--    PbFilletCompute
----------------------------------------------------------

enumeration ErrorTypeStatus  is  EmptyList, EdgeNotG1,FacesNotG1,EdgeNotOnShape,
                                 NotSharpEdge, PbFilletCompute                    
end  ErrorTypeStatus ;



--  this class is the API giving geometric informations about fillets:
 
    class Builder; 


-- this class is private and is only used by the class Builder:


    private class InternalBuilder;
    

end FilletSurf;
















