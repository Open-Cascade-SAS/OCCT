-- File:	RWStepFEA_RWNodeGroup.cdl
-- Created:	Thu Dec 12 17:51:06 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWNodeGroup from RWStepFEA

    ---Purpose: Read & Write tool for NodeGroup

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    NodeGroup from StepFEA

is
    Create returns RWNodeGroup from RWStepFEA;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : NodeGroup from StepFEA);
	---Purpose: Reads NodeGroup

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: NodeGroup from StepFEA);
	---Purpose: Writes NodeGroup

    Share (me; ent : NodeGroup from StepFEA;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWNodeGroup;
