-- Created on: 1993-08-06
-- Created by: Denis PASCAL
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package GraphDS 

    ---Purpose: This  package  <GraphDS> provides  generic  classes to
    --          describe transient graph data structure.

uses Standard,
     MMgt,
     TCollection,
     TColStd

is
    enumeration EntityRole is 
    	OnlyInput, 
    	OnlyOutput, 
    	InputAndOutput
    end EntityRole;
    
    enumeration RelationRole is 
        OnlyFront, 
    	OnlyBack, 
    	FrontAndBack
    end RelationRole;

    class EntityRoleMap instantiates DataMap from TCollection
                                    (Transient  from Standard,
				     EntityRole from GraphDS,
				     MapTransientHasher from TColStd);

    generic class DirectedGraph,
                  Vertex,
		  Edge,
		  VerticesIterator,
		  EdgesIterator;
		 
    
    generic class RelationGraph,
                  Entity,
		  Relation,
    	    	  EntitiesIterator,
                  IncidentEntitiesIterator,
                  RelationsIterator,
                  IncidentRelationsIterator;		  

end GraphDS;










