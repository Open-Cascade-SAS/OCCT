-- Created on: 1998-02-11
-- Created by: Philippe MANGIN
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

private  class SectionPlacement from BRepFill 

	---Purpose: Place a shape in a local axis coordinate         

uses 
    LocationLaw  from  BRepFill,
    Shape        from  TopoDS, 
    Trsf   from  gp

is 
   Create(Law             :  LocationLaw  from  BRepFill; 
          Section         :  Shape        from  TopoDS;  
          WithContact     :  Boolean  =  Standard_False; 
          WithCorrection  :  Boolean  =  Standard_False)  
	   ---Purpose: Automatic placement         
   returns   SectionPlacement from  BRepFill;   
    
   Create(Law             :  LocationLaw  from  BRepFill; 
          Section         :  Shape        from  TopoDS; 
	  Vertex          :  Shape        from  TopoDS;   
          WithContact     :  Boolean  =  Standard_False; 
          WithCorrection  :  Boolean  =  Standard_False)  
	   ---Purpose: Placement on vertex       
   returns   SectionPlacement from  BRepFill;     
   
   Perform(me:in  out; 
           WithContact :  Boolean;  
           WithCorrection :  Boolean;
    	   Vertex         :  Shape        from  TopoDS)   
    is  private; 
    
   Transformation(me) 
   ---C++: return const &    
   returns  Trsf  from  gp;   
    
   AbscissaOnPath(me:in  out)   
   returns  Real;

fields
    myLaw :  LocationLaw  from  BRepFill; 
    mySection  :  Shape from  TopoDS; 
    myTrsf     :  Trsf  from  gp; 
    myParam    :  Real; 
    myIndex    :  Integer;
end SectionPlacement;
