-- Created on: 2014-03-15
-- Created by: Laurent PAINNOT
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class NewtonFunctionRoot from math 
     ---Purpose:
     -- This class implements the calculation of a root of a function of
     -- a single variable starting from an initial near guess using the
     -- Newton algorithm. Knowledge of the derivative is required.


uses Vector from math, Matrix from math,
     FunctionWithDerivative from math,
     OStream from Standard
     
raises NotDone from StdFail

is 

    Create(F: in out FunctionWithDerivative;
    	   Guess, EpsX, EpsF: Real;
	   NbIterations: Integer = 100)
    ---Purpose:
    -- The Newton method is done to find the root of the function F 
    -- from the initial guess Guess.
    -- The tolerance required on the root is given by Tolerance.
    -- The solution is found when :
    --  abs(Xi - Xi-1) <= EpsX and abs(F(Xi))<= EpsF
    -- The maximum number of iterations allowed is given by NbIterations.
    returns NewtonFunctionRoot;


    Create(F: in out FunctionWithDerivative;
    	   Guess, EpsX, EpsF, A, B: Real;
	   NbIterations: Integer = 100)
    ---Purpose:
    -- The Newton method is done to find the root of the function F 
    -- from the initial guess Guess.
    -- The solution must be inside the interval [A, B].
    -- The tolerance required on the root is given by Tolerance.
    -- The solution is found when :
    --  abs(Xi - Xi-1) <= EpsX and abs(F(Xi))<= EpsF
    -- The maximum number of iterations allowed is given by NbIterations.
    returns NewtonFunctionRoot;


    Create(A, B, EpsX, EpsF: Real; 
           NbIterations: Integer = 100)
        ---Purpose: is used in a sub-class to initialize correctly all the fields
        --          of this class.

    returns NewtonFunctionRoot;
    

    Perform(me: in out; F: in out FunctionWithDerivative;
    	    Guess: Real)
        ---Purpose: is used internally by the constructors.

    is static;


    IsDone(me)
    	---Purpose: Returns true if the computations are successful, otherwise returns false.
      	---C++: inline
  returns Boolean
    is static;
    
    
    Root(me)
    	---Purpose: Returns the value of the root of function <F>.
        -- Exception NotDone is raised if the root was not found.
    	---C++: inline

    returns Real
    raises NotDone
    is static;
    

    Derivative(me)
    	---Purpose: returns the value of the derivative at the root.
        -- Exception NotDone is raised if the root was not found.
    	---C++: inline
    returns Real
    raises NotDone
    is static;
    

    Value(me)
    	---Purpose: returns the value of the function at the root.
        -- Exception NotDone is raised if the root was not found.
    	---C++: inline
    returns Real
    raises NotDone
    is static;
    

    NbIterations(me)
        ---Purpose: Returns the number of iterations really done on the 
        -- computation of the Root.
        -- Exception NotDone is raised if the root was not found.
    	---C++: inline
    returns Integer
    raises NotDone
    is static;


    Dump(me; o:in out OStream)
    	---Purpose: Prints information on the current state of the object.

    is static;


fields

Done: Boolean;
X   : Real;
Fx  : Real;
DFx : Real;
It  : Integer;
EpsilonX: Real;
EpsilonF: Real;
Itermax: Integer;
Binf: Real;
Bsup: Real;

end NewtonFunctionRoot;

