-- Created on: 1992-11-10
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class PathPoint from IntSurf 

	---Purpose: 

uses Pnt           from gp,
     Vec           from gp,
     Dir2d         from gp,
     HSequenceOfXY from TColgp

raises UndefinedDerivative from StdFail,
       OutOfRange          from Standard

is

    Create
    
    	returns PathPoint from IntSurf;


    Create (P: Pnt from gp; U,V: Real from Standard)
    
    	returns PathPoint from IntSurf;


    SetValue (me: in out; P: Pnt from gp; U,V: Real from Standard)
    
    	is static;


    AddUV(me: in out; U,V : Real from Standard)
    
	---C++: inline

    	is static;
	

    SetDirections(me: in out; V: Vec from gp; D: Dir2d from gp)
    
	---C++: inline

    	is static;
	

    SetTangency(me: in out; Tang: Boolean from Standard)
    
	---C++: inline

    	is static;



    SetPassing(me: in out; Pass: Boolean from Standard)
    
	---C++: inline

    	is static;


    Value(me)
    
    	returns Pnt from gp
	---C++: return const &
	---C++: inline

	is static;


    Value2d(me; U,V: out Real from Standard)
    
	---C++: inline
    	is static;


    IsPassingPnt(me)
    
    	returns Boolean from Standard
	---C++: inline

	is static;


    IsTangent(me)
    
    	returns Boolean from Standard
	---C++: inline

	is static;


    Direction3d(me)
    
    	returns Vec from gp
	---C++: return const &
	---C++: inline

	raises UndefinedDerivative from StdFail
	is static;


    Direction2d(me)
    
    	returns Dir2d from gp
	---C++: return const &
	---C++: inline

	raises UndefinedDerivative from StdFail
	is static;


    Multiplicity(me)
    
    	returns Integer from Standard
	---C++: inline

	is static;


    Parameters(me; Index: Integer from Standard;
                   U,V: out Real from Standard)

	---C++: inline

    	raises OutOfRange from Standard
    	is static;


fields

    pt     : Pnt           from gp;
    ispass : Boolean       from Standard;
    istgt  : Boolean       from Standard;
    vectg  : Vec           from gp;
    dirtg  : Dir2d         from gp;
    sequv  : HSequenceOfXY from TColgp;

end PathPoint;
