-- Created on: 1995-02-23
-- Created by: Mister rmi
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SensitivePoint from Select3D 
inherits SensitiveEntity from Select3D

	---Purpose: A framework to define sensitive 3D points.

uses
    Pnt             from gp,
    Pnt2d           from gp,
    Projector       from Select3D,
    Lin             from gp,
    EntityOwner     from SelectBasics,
    ListOfBox2d     from SelectBasics,
    PickArgs        from SelectBasics,
    Location        from TopLoc,
    Box2d             from Bnd,
    Array1OfPnt2d     from TColgp, 
    Pnt               from Select3D,
    Pnt2d             from Select3D

is

    Create (OwnerId : EntityOwner from SelectBasics;
    	    Point   : Pnt from gp)
    returns mutable SensitivePoint;
    	---Purpose: Constructs a sensitive point object defined by the
    	-- owner OwnerId and the point Point. 


    Project (me:mutable;aProjector : Projector from Select3D) 
    is redefined static;
    ---Level: Public 
    ---Purpose:Converts the stored 3D point into a 2D point according 
    --         to <aProjector> ; this method is called by the selection Manager.

    
    Areas(me:mutable; aresult : in out ListOfBox2d from SelectBasics) 
    is redefined static;
    ---Level: Public 
    ---Purpose: stores in <aresult> the 2D sensitive box which represents 
    --          the point area in the selection process. 

    GetConnected(me:mutable;aLocation: Location from TopLoc)
    returns SensitiveEntity from Select3D is redefined static;

    Matches (me : mutable;
             thePickArgs : PickArgs from SelectBasics;
             theMatchDMin, theMatchDepth : out Real from Standard)
    returns Boolean is redefined static;
    ---Level: Public
    ---Purpose: Checks whether the sensitive entity matches the picking
    -- detection area (close to the picking line).
    -- For details please refer to base class declaration.

    Matches (me  :mutable; 
             XMin,YMin,XMax,YMax : Real from Standard;
             aTol: Real from Standard) 
    returns Boolean
    is static;

     
    Matches (me  :mutable; 
             Polyline:Array1OfPnt2d from TColgp;
	     aBox:Box2d from Bnd;
             aTol: Real from Standard) 
    returns Boolean
    is redefined virtual;
    ---Level: Public 
    

    ComputeDepth(me;EyeLine: Lin from gp) 
    returns Real from Standard;

      
    Point(me) returns Pnt from gp;
    ---Purpose: Returns the point used at the time of construction.


    Dump(me; S: in out OStream;FullDump : Boolean from Standard = Standard_True) is redefined virtual;

fields

    mypoint   : Pnt from Select3D;
    myprojpt  : Pnt2d from Select3D;
    
    
end SensitivePoint;


