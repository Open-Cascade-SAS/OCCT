-- Created on: 1993-01-09
-- Created by: CKY / Contract Toubro-Larsen ( Deepak PRABHU )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package IGESDimen

        ---Purpose : This package represents Entities applied to Dimensions
        --           ie. Annotation Entities and attached Properties and
        --           Associativities.

uses

        Standard, 
        TCollection, 
        gp,
	TColStd,
	TColgp,
	Message,
        Interface, 
        IGESData, 
        IGESBasic,
        IGESGraph,
        IGESGeom

is

        class CenterLine;                  

        class Section;                     

        class WitnessLine;                 

        class AngularDimension;            

        class CurveDimension;              

        class DiameterDimension;           

        class FlagNote;                    

        class GeneralLabel;                

        class GeneralNote;                 

        class NewGeneralNote;              

        class LeaderArrow;                 

        class LinearDimension;            

        class OrdinateDimension;           

        class PointDimension;              

        class RadiusDimension;             

        class GeneralSymbol;               

        class SectionedArea;               

        class DimensionedGeometry;         

        class NewDimensionedGeometry;      

        class DimensionUnits;              

        class DimensionTolerance;          

        class DimensionDisplayData;        

        class BasicDimension;              

    	--    Tools for Entities    --

        class ToolCenterLine;
        class ToolSection;
        class ToolWitnessLine;                 
        class ToolAngularDimension;            
        class ToolCurveDimension;              
        class ToolDiameterDimension;           
        class ToolFlagNote;                    
        class ToolGeneralLabel;                
        class ToolGeneralNote;                 
        class ToolNewGeneralNote;              
        class ToolLeaderArrow;                 
        class ToolLinearDimension;            
        class ToolOrdinateDimension;           
        class ToolPointDimension;              
        class ToolRadiusDimension;             
        class ToolGeneralSymbol;               
        class ToolSectionedArea;               
        class ToolDimensionedGeometry;         
        class ToolNewDimensionedGeometry;      
        class ToolDimensionUnits;              
        class ToolDimensionTolerance;          
        class ToolDimensionDisplayData;        
        class ToolBasicDimension;              

    -- Definition and Exploitation of Entities defined in this Package

    class Protocol;
    class ReadWriteModule;
    class GeneralModule;
    class SpecificModule;

    -- Instantiations :

    class  Array1OfLeaderArrow instantiates
    	 Array1 from TCollection (LeaderArrow);
    class  Array1OfGeneralNote instantiates
    	 Array1 from TCollection (GeneralNote);

    class HArray1OfLeaderArrow instantiates
    	HArray1 from TCollection (LeaderArrow,Array1OfLeaderArrow);
    class HArray1OfGeneralNote instantiates
    	HArray1 from TCollection (GeneralNote,Array1OfGeneralNote);

    -- Package Methods

    Init;
    ---Purpose : Prepares dynamic data (Protocol, Modules) for this package

    Protocol  returns Protocol from IGESDimen;
    ---Purpose : Returns the Protocol for this Package

end IGESDimen;
