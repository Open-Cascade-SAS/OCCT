-- File:	MakeEllipse.cdl
-- Created:	Mon Sep 28 11:49:44 1992
-- Author:	Remi GILET
--		<reg@sdsun2>
---Copyright:	 Matra Datavision 1992

class MakeEllipse from GC inherits Root from GC

    	---Purpose :This class implements construction algorithms for an ellipse in
    	-- 3D space. The result is a Geom_Ellipse ellipse.
    	-- A MakeEllipse object provides a framework for:
    	-- -   defining the construction of the ellipse,
    	-- -   implementing the construction algorithm, and
    	-- -   consulting the results. In particular, the Value
    	--   function returns the constructed ellipse.

uses Pnt     from gp,
     Ax2     from gp,
     Hypr    from gp,
     Ellipse from Geom,
     Elips   from gp

raises NotDone from StdFail

is

Create (E : Elips from gp)  returns MakeEllipse;
    	--- Purpose :
    	--  Creates an ellipse from a non persistent ellipse E from package gp by its conversion. 

Create (A2                       : Ax2  from gp      ; 
    	MajorRadius, MinorRadius : Real from Standard) returns MakeEllipse;
    	--- Purpose : Constructs an ellipse with major and minor radii MajorRadius and
    	--   MinorRadius, and located in the plane defined by
    	--   the "X Axis" and "Y Axis" of the coordinate system A2, where:
    	--   -   its center is the origin of A2, and
    	--   -   its major axis is the "X Axis" of A2;
	--  Warnings :
	--  The MakeEllipse class does not prevent the
    	-- construction of an ellipse where MajorRadius is equal to MinorRadius.
    	-- If an error occurs (that is, when IsDone returns
    	-- false), the Status function returns:
    	-- -   gce_InvertRadius if MajorRadius is less than MinorRadius;
    	-- -   gce_NegativeRadius if MinorRadius is less than 0.0;
    	-- -   gce_NullAxis if the points S1 and Center are coincident; or
    	-- -   gce_InvertAxis if:
    	--   -   the major radius computed with Center and S1
    	--    is less than the minor radius computed with Center, S1 and S2, or
    	--   -   Center, S1 and S2 are collinear.

Create(S1,S2  : Pnt from gp;
       Center : Pnt from gp) returns MakeEllipse;
	---Purpose: Constructs an ellipse centered on the point Center, where
    	--   -   the plane of the ellipse is defined by Center, S1 and S2,
    	--   -   its major axis is defined by Center and S1,
    	--   -   its major radius is the distance between Center and S1, and
    	--   -   its minor radius is the distance between S2 and the major axis.
		
Value(me) returns Ellipse from Geom
    raises NotDone
    is static;
    	---Purpose: Returns the constructed ellipse.
    	-- Exceptions StdFail_NotDone if no ellipse is constructed.
        ---C++: return const&

Operator(me) returns Ellipse from Geom
    is static;
    	---C++: return const&
    	---C++: alias "Standard_EXPORT operator Handle_Geom_Ellipse() const;"

fields

    TheEllipse : Ellipse from Geom;
    --The solution from Geom.
    
end MakeEllipse;
