-- Created on: 1995-03-15
-- Created by: Christian CAILLET
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package  XSDRAWIGES

    ---Purpose : XSDRAW for IGES : commands IGESSelect, Controller, transfer

uses Standard, Interface, Transfer, IFSelect, IGESControl  , Draw

is

--    class Controller;  see IGESControl

    InitSelect;
    ---Purpose : Inits IGESSelect commands, for DRAW

    InitToBRep   (theCommands : in out Interpretor from Draw);
    ---Purpose : Inits IGESToBRep for DRAW

    InitFromBRep (theCommands : in out Interpretor from Draw);
    ---Purpose : Inits BRepToIGES for DRAW

end XSDRAWIGES;
