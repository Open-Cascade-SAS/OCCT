-- Created on: 1997-04-17
-- Created by: Christophe MARION
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Hider from HLRBRep

uses
    Integer         from Standard,
    Boolean         from Standard,
    Real            from Standard,
    ShortReal       from Standard,
    ListOfInteger   from TColStd,
    MapOfShapeTool  from BRepTopAdaptor,
    Data            from HLRBRep

is
    Create(DS : Data from HLRBRep)
    returns Hider from HLRBRep;
	---Purpose: Creates a Hider processing  the set  of  Edges and
	--          hiding faces described by <DS>.  Stores the hidden
	--          parts in <DS>.

    OwnHiding(me : in out; FI : Integer from Standard)
	---Purpose: own hiding the side face number <FI>.
    is static;

    Hide(me : in out; FI :        Integer from Standard;
                      MST: in out MapOfShapeTool from BRepTopAdaptor)
	---Purpose: Removes from the edges,   the parts hidden by  the
	--          hiding face number <FI>.
    is static;

fields
    myDS : Data from HLRBRep;

end Hider;
