-- Created on: 2001-07-17
-- Created by: Julia DOROVSKIKH <jfa@hotdox.nnov.matra-dtv.fr>
-- Copyright (c) 2001-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Persistent from XmlObjMgt

uses
    Element from XmlObjMgt,
    DOMString from XmlObjMgt

is
    Create      returns Persistent from XmlObjMgt;
      ---Purpose: empty constructor

    Create (theElement : Element from XmlObjMgt)
                returns Persistent from XmlObjMgt;
      ---Purpose: constructor

    Create (theElement : Element from XmlObjMgt;
            theRef     : DOMString from XmlObjMgt)
                returns Persistent from XmlObjMgt;
      ---Purpose: constructor from sub-element of Element referenced by theRef

    CreateElement (me:in out; theParent: out Element   from XmlObjMgt;
                              theType:       DOMString from XmlObjMgt;
                              theID:         Integer   from Standard);
      ---Purpose: myElement := <theType id="theID"/>

    SetId (me:in out; theId: Integer from Standard)
    is static;
      ---Level: Internal

    Element (me) returns Element from XmlObjMgt;
      ---C++: inline
      ---C++: return const &
      ---C++: alias "inline operator const XmlObjMgt_Element&() const;"
      ---Purpose: return myElement

    Element (me:in out) returns Element from XmlObjMgt;
      ---C++: inline
      ---C++: return &
      ---C++: alias "inline operator XmlObjMgt_Element&();"
      ---Purpose: return myElement

    Id(me) returns Integer from Standard
    is static;
      ---C++: inline
      ---Level: Internal

fields
    myElement: Element from XmlObjMgt;
    myID     : Integer from Standard;

end Persistent;
