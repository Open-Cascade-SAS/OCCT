-- Created on: 1993-06-23
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SurfaceCurveInterference from TopOpeBRepDS 
    inherits Interference from TopOpeBRepDS

    ---Purpose: an interference with a 2d curve

uses

    Transition  from TopOpeBRepDS,
    Kind        from TopOpeBRepDS,
    Curve       from Geom2d,
    OStream     from Standard
    
is

    Create returns mutable SurfaceCurveInterference from TopOpeBRepDS;

    Create(Transition   : Transition from TopOpeBRepDS;
	   SupportType  : Kind from TopOpeBRepDS;
	   Support      : Integer;
	   GeometryType : Kind from TopOpeBRepDS;
	   Geometry     : Integer;
    	   PC : Curve from Geom2d) 
    returns mutable SurfaceCurveInterference from TopOpeBRepDS; 

    Create(I : Interference from TopOpeBRepDS)
    returns mutable SurfaceCurveInterference from TopOpeBRepDS; 
	    
    PCurve(me) returns any Curve from Geom2d is static;
	---C++: return const &

    PCurve(me : mutable; PC : Curve from Geom2d) is static;

    DumpPCurve(me; OS : in out OStream from Standard; 
                   compact : Boolean = Standard_True)
    ---C++: return &
    returns OStream from Standard
    is static;

    Dump(me; OS : in out OStream from Standard)
    ---C++: return &
    returns OStream from Standard
    is redefined;
    
fields

    myPCurve : Curve from Geom2d;

end SurfaceCurveInterference from TopOpeBRepDS;
