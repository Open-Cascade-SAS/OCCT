-- Created on: 1993-09-28
-- Created by: Bruno DUMORTIER
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Filling from GeomFill
	---Purpose: Root class for Filling;

uses
    Array1OfPnt    from TColgp,
    Array2OfPnt    from TColgp,
    HArray2OfPnt   from TColgp,
    Array1OfReal   from TColStd,
    Array2OfReal   from TColStd,
    HArray2OfReal  from TColStd
    
raises
    NoSuchObject from Standard

is
    Create;
    
    NbUPoles(me) returns Integer from Standard
    is static;
    
    NbVPoles(me) returns Integer from Standard
    is static;

    Poles(me; Poles : in out Array2OfPnt from TColgp)
    is static;
    
    isRational(me) returns Boolean from Standard
    is static;
    
    Weights(me; Weights : in out Array2OfReal from TColStd)
    raises
    	NoSuchObject from Standard
    is static;    
    
    
fields
    
    IsRational : Boolean        from Standard is protected;
    myPoles    : HArray2OfPnt   from TColgp   is protected;
    myWeights  : HArray2OfReal  from TColStd  is protected;

end Filling;
