-- Created on: 1998-12-09
-- Created by: Xuan PHAM PHU
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class connexity from TopOpeBRepTool

uses 
    Shape from TopoDS,
    ListOfShape from TopTools,
    Array1OfListOfShape from TopTools
is
    Create returns connexity from TopOpeBRepTool;
    Create (Key : Shape from TopoDS) returns connexity from TopOpeBRepTool;
    SetKey (me : in out; Key : Shape from TopoDS);	        	
    Key (me) returns Shape from TopoDS;
    ---C++: return const &
    
    Item(me; OriKey : Integer; Item : out ListOfShape from TopTools) 
    returns Integer;
    -- if <theKey> is oriented <OriKey> in all shapes of <Item>, returns
    -- the <Item>'s length.
    
    AllItems(me; Item : out ListOfShape from TopTools)
    returns Integer;
    -- returns all items attached to <theKey>
    
    AddItem(me : in out; OriKey : Integer; Item : ListOfShape from TopTools);
    AddItem(me : in out; OriKey : Integer; Item : Shape from TopoDS);
    RemoveItem(me : in out; OriKey : Integer; Item : Shape from TopoDS)
    returns Boolean;
    -- returns true if <Item> is stored in the list.
    RemoveItem(me : in out; Item : Shape from TopoDS)
    returns Boolean;
    
    ChangeItem(me : in out; OriKey : Integer)
    returns ListOfShape from TopTools;
    ---C++: return & 
   
    IsMultiple(me)
    returns Boolean;
    -- returns true if <theKey> is multiple.   

    IsFaulty(me)
    returns Boolean;

    IsInternal(me; Item : out ListOfShape from TopTools)
    returns Integer;
    -- <theKey> is INTERNAL in shapes of <Item> oriented FORWARD.
    
fields
    theKey : Shape from TopoDS;
    theItems : Array1OfListOfShape from TopTools; 
	-- <theKey> is FORWARD in shapes of theItems(1)  
	-- <theKey> is REVERSED in shapes of theItems(2)  
	-- <theKey> is INTERNAL in shapes of theItems(3)  
	-- <theKey> is EXTERNAL in shapes of theItems(4) 
	-- <theKey> appears FORWARD and REVERSED in shapes of theItems(5)  
end connexity;
