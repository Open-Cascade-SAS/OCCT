-- Created on: 2000-04-09
-- Created by: Sergey MOZOKHIN
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package STEPCAFControl

    ---Purpose : This package provides external access and control for STEP,
    --           on the level of CAF (shapes with attributes, external 
    --           references etc.)

uses 
    Dico,
    TCollection,
    TColStd,
    TopTools,
    TopoDS,
    IFSelect,
    Transfer,
    XSControl,
    STEPControl,
    STEPConstruct,
    StepShape,
    StepRepr,
    StepBasic,
    ShapeBuild,
    TDF,
    TDocStd,
    XCAFDoc,
    MoniTool

is

    class Reader;
    	---Purpose: Reader for DECAF documents
    
    class Writer;
    	---Purpose: Writer for DECAF documents

    class ExternFile;
        ---Purpose: Auxiliary class to store results of translation of external file

    class ActorWrite;
    class Controller;
    	---Purpose: Extensions of standard STEP tools for DECAF specifics
    
    class DictionaryOfExternFile instantiates 
    	  Dictionary from Dico (ExternFile from STEPCAFControl);

    class DataMapOfShapeSDR instantiates 
    	  DataMap from TCollection (Shape from TopoDS,
	    	    	    	    ShapeDefinitionRepresentation from StepShape,
				    ShapeMapHasher from TopTools);

    --- skl
    class DataMapOfShapePD instantiates 
    	  DataMap from TCollection (Shape from TopoDS,
	    	    	    	    ProductDefinition from StepBasic,
				    ShapeMapHasher from TopTools);

    class DataMapOfSDRExternFile instantiates 
    	  DataMap from TCollection (ShapeDefinitionRepresentation from StepShape,
				    ExternFile from STEPCAFControl,
				    MapTransientHasher from TColStd);

    --- skl
    class DataMapOfPDExternFile instantiates 
    	  DataMap from TCollection (ProductDefinition from StepBasic,
				    ExternFile from STEPCAFControl,
				    MapTransientHasher from TColStd);

    class DataMapOfLabelShape instantiates
    	  DataMap from TCollection (Label from TDF,
				    Shape from TopoDS,
	    	    	    	    LabelMapHasher from TDF);

    class DataMapOfLabelExternFile instantiates
    	  DataMap from TCollection (Label from TDF,
				    ExternFile from STEPCAFControl,
	    	    	    	    LabelMapHasher from TDF);

end STEPCAFControl;
