-- Created on: 2007-05-29
-- Created by: Vlad Romashko
-- Copyright (c) 2007-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ReferenceListDriver from XmlMDataStd inherits ADriver from XmlMDF

uses

    SRelocationTable from XmlObjMgt,
    RRelocationTable from XmlObjMgt,
    Persistent       from XmlObjMgt,
    MessageDriver    from CDM,
    Attribute        from TDF

is

    Create (theMessageDriver:MessageDriver from CDM)
    returns mutable ReferenceListDriver from XmlMDataStd;

    NewEmpty (me)
    returns mutable Attribute from TDF;

    Paste(me; Source     : Persistent from XmlObjMgt;
              Target     : mutable Attribute from TDF;
              RelocTable : out RRelocationTable from XmlObjMgt)
    returns Boolean from Standard;

    Paste(me; Source     : Attribute from TDF;
              Target     : in out Persistent from XmlObjMgt;
              RelocTable : out SRelocationTable from XmlObjMgt);

end ReferenceListDriver;
