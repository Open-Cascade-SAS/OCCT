-- Created on: 1994-10-28
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class FaceEdgeInterference from TopOpeBRepDS 
    inherits ShapeShapeInterference from TopOpeBRepDS

uses

    Transition from TopOpeBRepDS,
    Config     from TopOpeBRepDS,
    OStream    from Standard    
    
is

    Create(T : Transition from TopOpeBRepDS;
	   S : Integer from Standard;
	   G : Integer from Standard;
      	   GIsBound : Boolean from Standard;
    	   C : Config from TopOpeBRepDS)
	   
    	---Purpose: Create an interference of EDGE <G> on FACE <S>.

    returns mutable FaceEdgeInterference from TopOpeBRepDS; 
	    
    Dump(me; OS : in out OStream from Standard) returns OStream
    is redefined;
    ---C++: return &
    
end FaceEdgeInterference from TopOpeBRepDS;
