-- Created on: 1997-05-21
-- Created by: Christian CAILLET
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class DescrGeneral  from StepData    inherits GeneralModule  from StepData

    ---Purpose : Works with a Protocol by considering its entity descriptions


uses Transient,
     EntityIterator from Interface,
     ShareTool      from Interface,
     Check          from Interface,
     CopyTool       from Interface,
     Protocol  from StepData

is

    Create (proto : Protocol from StepData) returns DescrGeneral;

    FillSharedCase (me; CN : Integer; ent : Transient;
        iter : in out EntityIterator);

    CheckCase (me; CN : Integer; ent : Transient; shares : ShareTool;
    	ach : in out Check);

    CopyCase (me; CN : Integer; entfrom : Transient; entto : mutable Transient;
    	TC : in out CopyTool);

    NewVoid (me; CN : Integer; ent : out mutable Transient) returns Boolean;

fields

    theproto : Protocol from StepData;

end DescrGeneral;
