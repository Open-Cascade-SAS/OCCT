-- Created on: 1994-11-14
-- Created by: Bruno DUMORTIER
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

private class MultiLine from BRepFill 

	---Purpose: Private class used to compute the 3d curve and the
	--          two 2d curves resulting from the intersection of a
	--          surface of linear extrusion( Bissec, Dz) and the 2
	--          faces.    
	--          This 3 curves will  have  the same parametrization 
	--          as the Bissectrice.
	--          This  class  is  to  be  send  to an approximation 
	--          routine. 

uses
    Face  from TopoDS,
    Edge  from TopoDS,
    Curve from Geom,
    Curve from Geom2d,
    Curve from Geom2dAdaptor,
    Pnt   from gp,
    Pnt2d from gp,
    Shape from GeomAbs
    
raises
    DomainError from Standard
    
is
    Create;
    
    Create( Face1, Face2 : Face    from TopoDS;
    	    Edge1, Edge2 : Edge    from TopoDS;
	    Inv1 , Inv2  : Boolean from Standard;
    	    Bissec       : Curve   from Geom2d );

    IsParticularCase(me)
    returns Boolean from Standard
	---Purpose: Search if the Projection of the Bissectrice on the
	--          faces needs an approximation or not.
	--          Returns true if the approximation is not needed.
    is static;

    Continuity (me) returns Shape from GeomAbs
	---Purpose: Returns   the continuity  betwwen  the two  faces
	--          seShape         from GeomAbsparated by myBis.
    is static;
	    
    Curves(me; Curve   : in out Curve from Geom;
    	       PCurve1 : in out Curve from Geom2d;
	       PCurve2 : in out Curve from Geom2d)
    raises 
    	DomainError from Standard
	---Purpose: raises if IsParticularCase is <False>.
    is static;

    FirstParameter(me) 
	---Purpose: returns the first parameter of the Bissectrice.
    returns Real from Standard is static;		    

    LastParameter(me) 
	---Purpose: returns the last parameter of the Bissectrice.
    returns Real from Standard is static;		    

    Value ( me; U : Real from Standard)
	---Purpose: Returns the current point on the 3d curve
    returns Pnt from gp is static;

    ValueOnF1(me; U : Real from Standard)
	---Purpose: returns the current point on the PCurve of the
	--          first face
    returns Pnt2d from gp is static;
	
    ValueOnF2(me; U : Real from Standard)
	---Purpose: returns the current point on the PCurve of the
	--          first face
    returns Pnt2d from gp is static;
    
    Value3dOnF1OnF2(me; 
    	    	    U   : Real         from Standard;
		    P3d : in out Pnt   from gp;
		    PF1 : in out Pnt2d from gp;
		    PF2 : in out Pnt2d from gp)
    is static;		    
		    	
	
fields
    myFace1 : Face    from TopoDS;
    myFace2 : Face    from TopoDS;
    myU1    : Curve   from Geom2dAdaptor;
    myV1    : Curve   from Geom2dAdaptor;
    myU2    : Curve   from Geom2dAdaptor;
    myV2    : Curve   from Geom2dAdaptor;
    myIsoU1 : Boolean from Standard;
    myIsoU2 : Boolean from Standard;
    myBis   : Curve   from Geom2dAdaptor;
    myKPart : Integer from Standard;
    myCont  : Shape   from GeomAbs;	
    
end MultiLine;
