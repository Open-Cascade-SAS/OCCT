-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class LoopAndPath from StepShape 

inherits TopologicalRepresentationItem from StepShape 


	--- This classe is an implementation of EXPRESS
	--  ANDOR Subtype Declaration.
uses

	Loop from StepShape, 
	Path from StepShape, 
	HAsciiString from TCollection, 
	HArray1OfOrientedEdge from StepShape, 
	OrientedEdge from StepShape
is

	Create returns mutable LoopAndPath;
	---Purpose: Returns a LoopAndPath


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aLoop : mutable Loop from StepShape;
	      aPath : mutable Path from StepShape) is virtual;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aEdgeList : mutable HArray1OfOrientedEdge from StepShape) is virtual;

	-- Specific Methods for Field Data Access --

	SetLoop(me : mutable; aLoop : mutable Loop);
	Loop (me) returns mutable Loop;
	SetPath(me : mutable; aPath : mutable Path);
	Path (me) returns mutable Path;

	-- Specific Methods for ANDOR Field Data Access --


	-- Specific Methods for ANDOR Field Data Access --

	SetEdgeList(me : mutable; aEdgeList : mutable HArray1OfOrientedEdge);
	EdgeList (me) returns mutable HArray1OfOrientedEdge;
	EdgeListValue (me; num : Integer) returns mutable OrientedEdge;
	NbEdgeList (me) returns Integer;

fields

	loop : Loop from StepShape;
	path : Path from StepShape;

end LoopAndPath;
