-- Created on: 1999-07-29
-- Created by: Roman LYGIN
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



package Message 

    	---Purpose: Defines
   	--          - tools to work with messages
    	--          - basic tools intended for progress indication

uses

    MMgt,
    TColStd,
    TCollection,
    Standard

is

    enumeration Gravity is
    	---Purpose: Defines gravity level of messages
	-- - Trace: low-level details on algorithm execution (usually for debug purposes)
	-- - Info: informative message
	-- - Warning: warning message
	-- - Alarm: non-critical error
	-- - Fail: fatal error 
	Trace,
        Info,
        Warning,
        Alarm,
	Fail
    end Gravity;

    imported Status;
    imported StatusType;
    imported ExecStatus;

    class Msg;
    	---Purpose: Defines message.
    class MsgFile;
    	---Purpose: Defines file storing messages.
	
    class Messenger;
    	---Purpose: Messenger is API class providing general-purpose interface for 
	--          libraries that may issue text messages without knowledge
	--          of how these messages will be further processed.
	
    class Algorithm;
	---Purpose: Class Message_Algorithm is the root class for all algorithms.
	--          It provides generic mechanism for management execution status,
	--          collection and output of corresponding error/warning messages

    deferred class Printer;
    	---Purpose: Defines basic message printer.
	
	class PrinterOStream;
	    ---Purpose: Defines printer associated with an ostream
    
    class ListOfMsg instantiates List from TCollection (Msg from Message);
    
    class SequenceOfPrinters instantiates 
    Sequence from TCollection (Printer from Message);

    -- Progress indication
    deferred class ProgressIndicator;
    class ProgressScale;
    class ProgressSentry;
    class SequenceOfProgressScale instantiates
         Sequence from TCollection (ProgressScale from Message);
    
    DefaultMessenger returns Messenger from Message;
        ---Purpose: Defines default messenger for OCCT applications.
        --          This is global static instance of the messenger.
	--          By default, it contains single printer directed to cout.
	--          It can be customized according to the application needs.
	---C++: return const &

    FillTime (Hour, Minute: Integer; Second: Real) returns AsciiString from TCollection;
    	---Purpose: Returns the string filled with values of hours, minutes and seconds.
	-- Example:
    	--          1. (5, 12, 26.3345) returns "05h:12m:26.33s",
	--          2. (0,  6, 34.496 ) returns "06m:34.50s",
	--          3. (0,  0,  4.5   ) returns "4.50s"

end Message;
