-- Created on: 1995-07-17
-- Created by: Stagiaire Alain JOURDAIN
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package IntPoly

    	  ---Purpose:


uses    Standard,
    	TCollection,
    	gp,
        TColStd,
	TColgp,
    	TopoDS,
    	TopAbs,
    	TopExp,
        TopLoc,
	Poly
	
is   class SequenceOfSequenceOfPnt2d
    	instantiates Sequence from TCollection (SequenceOfPnt2d from TColgp);

     class Pnt2dHasher;

     class IndexedMapOfPnt2d
     	instantiates IndexedMap from TCollection (Pnt2d       from gp,
                                                  Pnt2dHasher from IntPoly);
        
     class PlaneSection;
     
     class SequenceOfSequenceOfPnt
    	instantiates Sequence from TCollection (SequenceOfPnt from TColgp);

     class PntHasher;

     class IndexedMapOfPnt
     	instantiates IndexedMap from TCollection (Pnt       from gp,
                                                  PntHasher from IntPoly);
        
     class ShapeSection;


end IntPoly;












