-- Created on: 1994-12-16
-- Created by: Frederic MAUPAS
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class TranslateEdge from StepToTopoDS
    inherits Root from StepToTopoDS
    
    ---Purpose:
    --         

uses

    Edge               from StepShape,
    Tool               from StepToTopoDS,
    TranslateEdgeError from StepToTopoDS,
    Shape              from TopoDS,
    Edge               from TopoDS,
    Vertex             from TopoDS,
    Curve              from Geom2d,
    Surface            from Geom,
    EdgeCurve          from StepShape,
    Curve              from StepGeom,
    Vertex             from StepShape,
    Pcurve             from StepGeom,
    NMTool             from StepToTopoDS

raises NotDone from StdFail

is

    Create returns TranslateEdge;
    
    Create (E      : Edge from StepShape;
            T      : in out Tool from StepToTopoDS;
            NMTool : in out NMTool from StepToTopoDS)
    	returns TranslateEdge;
	    
    Init (me     : in out;
          E      : Edge from StepShape;
          T      : in out Tool from StepToTopoDS;
          NMTool : in out NMTool from StepToTopoDS);

    MakeFromCurve3D (me : in out; C3D : Curve from StepGeom;
    	    	     EC     : EdgeCurve from StepShape;        -- for messages
		     Vend   : Vertex from StepShape;      -- case of null edge
		     preci  : Real; E : in out Edge from TopoDS;
		     V1, V2 : in out Vertex from TopoDS;
		     T      : in out Tool from StepToTopoDS);
    ---Purpose:  Warning! C3D is assumed to be a Curve 3D ...
    --    other cases to checked before calling this

    MakePCurve (me; PCU : Pcurve from StepGeom; ConvSurf : Surface from Geom)
    	returns Curve from Geom2d;
    --  Null if failed

    Value (me) returns Shape from TopoDS
    	raises NotDone
	is static;
	---C++: return const &

    Error (me) returns TranslateEdgeError from StepToTopoDS;
    
fields

    myError  : TranslateEdgeError from StepToTopoDS;
    
    myResult : Shape              from TopoDS;
    
end TranslateEdge;
