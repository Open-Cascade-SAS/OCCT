-- Created on: 2000-05-18
-- Created by: Peter KURNEV
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Range from IntTools 

	---Purpose: The class describes the  1-d range 
        --          [myFirst, myLast].  	 

--uses
is 
    Create   
    	returns  Range from IntTools ;
	---Purpose:
	--- Empty constructor
	---
     
    Create  (aFirst:Real  from  Standard;  aLast:Real  from  Standard) 
    	returns  Range from IntTools ; 
	---Purpose:
	--- Initialize me by range boundaries
	---
	 
    SetFirst(me:out; aFirst:Real  from  Standard); 
    	---Purpose:
	--- Modifier
	---
     
    SetLast (me:out; aLast:Real  from  Standard);  
    	---Purpose:
	--- Modifier
	---
     
    First   (me) 
    	returns  Real  from  Standard; 
	---Purpose:
	--- Selector
	---
     
    Last   (me) 
    	returns  Real  from  Standard;  
	---Purpose:
	--- Selector
	---
	 
    Range  (me; aFirst:out Real  from  Standard;   
    	    	aLast :out Real  from  Standard);
    	---Purpose:
	--- Selector
	---
	    	
fields
    myFirst:  Real  from  Standard;
    myLast :  Real  from  Standard;
end Range;
