-- File:	RWStepElement_RWSurfaceElementProperty.cdl
-- Created:	Thu Dec 12 17:29:04 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWSurfaceElementProperty from RWStepElement

    ---Purpose: Read & Write tool for SurfaceElementProperty

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    SurfaceElementProperty from StepElement

is
    Create returns RWSurfaceElementProperty from RWStepElement;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : SurfaceElementProperty from StepElement);
	---Purpose: Reads SurfaceElementProperty

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: SurfaceElementProperty from StepElement);
	---Purpose: Writes SurfaceElementProperty

    Share (me; ent : SurfaceElementProperty from StepElement;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWSurfaceElementProperty;
