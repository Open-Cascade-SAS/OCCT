-- Created on: 1996-01-26
-- Created by: Philippe MANGIN
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

private class BattenLaw from FairCurve inherits Function from math

	---Purpose: This class compute the Heigth of an batten 

is
     Create(Heigth, Slope, Sliding : Real)
    ---Purpose: Constructor of linear batten with
    --          Heigth : the Heigth at the middle point
    --          Slope  : the geometric slope of the batten
    --          Sliding : Active Length of the batten without extension
     returns BattenLaw;
     
     SetSliding(me : in out; Sliding : Real);
     ---Purpose: Change the value of sliding
     ---C++: inline
     
     SetHeigth(me : in out; Heigth : Real);
     ---Purpose: Change the value of Heigth at the middle point.
     ---C++: inline
     
     SetSlope(me : in out; Slope : Real);
     ---Purpose: Change the value of the geometric slope.
     ---C++: inline
     
    
     Value(me: in out; T: Real; THeigth: out Real) returns Boolean
     ---Purpose: computes the value of  the heigth for the parameter T
     --          on  the neutral fibber
     ---C++: inline
     is redefined;




fields
MiddleHeigth   : Real; -- the Heigth at the middle point
GeometricSlope : Real; -- the geometric slope of the batten
LengthSliding  : Real; -- the length of sliding of the batten
end BattenLaw;
