-- Created on: 1997-02-05
-- Created by: Alexander BRIVIN
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Instancing from Vrml 

	---Purpose: defines  "instancing" - using  the  same  instance  of  a  node   
	--          multiple  times.
	--  It  is  accomplished  by  using  the  "DEF"  and  "USE"  keywords.      
    	--  The  DEF  keyword  both  defines  a  named  node,  and  creates  a  single 
	--  instance  of  it.   
    	--  The  USE  keyword  indicates  that  the  most  recently  defined  instance 
    	--  should  be  used  again.   
    	--  If  several  nades  were  given  the  same  name,  then  the  last  DEF 
	--  encountered  during  parsing  "wins". 
	--  DEF/USE  is  limited  to  a  single  file.
uses

     AsciiString from TCollection

is
 
    Create ( aString        : AsciiString from TCollection ) 
        returns Instancing from Vrml;
 
        ---Purpose: Adds "DEF  <myName>" in  anOStream  (VRML  file).
    DEF ( me;  anOStream: in out OStream from Standard) returns OStream from Standard;
    ---C++:  return  & 

        ---Purpose: Adds "USE  <myName>" in  anOStream (VRML  file).
    USE ( me;  anOStream: in out OStream from Standard) returns OStream from Standard;
    ---C++:  return  & 

fields
 
    myName  : AsciiString from TCollection;  --  Name  using  DEF/USE  for a  node

end Instancing;

