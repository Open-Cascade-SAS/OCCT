-- Created on: 2001-12-20
-- Created by: Pavel TELKOV
-- Copyright (c) 2001-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Curve2d from ShapeCustom 

	---Purpose: Converts curve2d to analytical form with given 
    	--          precision or simpify curve2d.
    	
uses
    Curve         from Geom2d,
    Line          from Geom2d,
    Array1OfPnt2d from TColgp,
    BSplineCurve  from Geom2d
is
    
    -- static methods
    IsLinear (myclass; thePoles : Array1OfPnt2d from TColgp;
    	    	       theTolerance : Real from Standard;
		       theDeviation : in out Real from Standard)
    returns Boolean from Standard;
    	---Purpose: Check if poleses is in the plane with given precision
    	--          Returns false if no.
	
    ConvertToLine2d (myclass; theCurve : Curve from Geom2d;
    	    	    	      theFirstIn, theLastIn : Real from Standard;
			      theTolerance : Real from Standard;
			      theNewFirst, theNewLast : in out Real from Standard;
			      theDeviation: in out Real from Standard)
    returns Line from Geom2d;
    	---Purpose: Try to convert BSpline2d or Bezier2d to line 2d
    	--          only if it is linear. Recalculate first and last parameters.
    	--          Returns line2d or null curve2d.

    SimplifyBSpline2d (myclass; theBSpline2d : in out BSplineCurve from Geom2d;
    	    	    	    	theTolerance : Real from Standard )
    returns Boolean from Standard;
    	---Purpose: Try to remove knots from bspline where local derivatives are the same.
    	--          Remove knots with given precision.
    	--          Returns false if Bsplien was not modified

--fields


end Curve2d;
