-- Created on: 1997-02-11
-- Created by: Alexander BRIVIN
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Texture2Transform from Vrml 

	---Purpose: defines a Texture2Transform node of VRML specifying properties of geometry
	---          and its appearance.
    	--  This  node  defines  a 2D  transformation  applied  to  texture  coordinates.   
	--  This  affect  the  way  textures  are  applied  to  the  surfaces  of  subsequent 
    	--  shapes. 
    	--  Transformation  consisits  of(in  order)  a  non-uniform  scale  about  an   
    	--  arbitrary  center  point,  a  rotation  about  that  same  point,  and 
	--  a  translation.  This  allows  a  user  to  change  the  size  and  position  of 
	--  the  textures  on  the  shape.
    	--  By  default  : 
	--    myTranslation (0 0)
	--    myRotation (0)
	--    myScaleFactor (1 1)
	--    myCenter (0 0) 
 
uses
 
   Vec2d from gp 

is
 
    Create  returns  Texture2Transform from Vrml;
 
    Create  ( aTranslation  :  Vec2d   from  gp;
    	      aRotation     :  Real    from  Standard; 
    	      aScaleFactor  :  Vec2d   from  gp;
    	      aCenter       :  Vec2d   from  gp ) 
        returns  Texture2Transform from Vrml;

    SetTranslation ( me : in out; aTranslation : Vec2d  from  gp );
    Translation ( me  )  returns  Vec2d  from  gp;

    SetRotation ( me : in out; aRotation : Real from Standard );
    Rotation ( me )  returns  Real from Standard;

    SetScaleFactor( me : in out; aScaleFactor : Vec2d  from  gp );
    ScaleFactor( me )  returns  Vec2d  from  gp;

    SetCenter ( me : in out; aCenter : Vec2d  from  gp );
    Center ( me )  returns  Vec2d  from  gp;

    Print  ( me;  anOStream: in out OStream from Standard) returns OStream from Standard;
    ---C++:  return  & 

fields
 
    myTranslation  :  Vec2d  from  gp;       -- Translation vector
    myRotation     :  Real   from  Standard; -- Rotation
    myScaleFactor  :  Vec2d  from  gp;       -- Scale factors
    myCenter       :  Vec2d  from  gp;       -- Center point for scale and rotate
    
end Texture2Transform;

