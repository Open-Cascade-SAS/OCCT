-- File:        SweptSurface.cdl
-- Created:     Fri Dec  1 11:11:29 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class SweptSurface from StepGeom 

inherits Surface from StepGeom 

uses

	Curve from StepGeom, 
	HAsciiString from TCollection
is

	Create returns mutable SweptSurface;
	---Purpose: Returns a SweptSurface


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aSweptCurve : mutable Curve from StepGeom) is virtual;

	-- Specific Methods for Field Data Access --

	SetSweptCurve(me : mutable; aSweptCurve : mutable Curve);
	SweptCurve (me) returns mutable Curve;

fields

	sweptCurve : Curve from StepGeom;

end SweptSurface;
