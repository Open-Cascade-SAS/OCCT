-- Created on: 2002-12-12
-- Created by: data exchange team
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class RepresentedDefinition from StepRepr
inherits SelectType from StepData

    ---Purpose: Representation of STEP SELECT type RepresentedDefinition

uses
    GeneralProperty from StepBasic,
    PropertyDefinition from StepRepr,
    PropertyDefinitionRelationship from StepRepr,
    ShapeAspect from StepRepr,
    ShapeAspectRelationship from StepRepr

is
    Create returns RepresentedDefinition from StepRepr;
	---Purpose: Empty constructor

    CaseNum (me; ent: Transient) returns Integer;
	---Purpose: Recognizes a kind of RepresentedDefinition select type
	--          1 -> GeneralProperty from StepBasic
	--          2 -> PropertyDefinition from StepRepr
	--          3 -> PropertyDefinitionRelationship from StepRepr
	--          4 -> ShapeAspect from StepRepr
	--          5 -> ShapeAspectRelationship from StepRepr
	--          0 else

    GeneralProperty (me) returns GeneralProperty from StepBasic;
	---Purpose: Returns Value as GeneralProperty (or Null if another type)

    PropertyDefinition (me) returns PropertyDefinition from StepRepr;
	---Purpose: Returns Value as PropertyDefinition (or Null if another type)

    PropertyDefinitionRelationship (me) returns PropertyDefinitionRelationship from StepRepr;
	---Purpose: Returns Value as PropertyDefinitionRelationship (or Null if another type)

    ShapeAspect (me) returns ShapeAspect from StepRepr;
	---Purpose: Returns Value as ShapeAspect (or Null if another type)

    ShapeAspectRelationship (me) returns ShapeAspectRelationship from StepRepr;
	---Purpose: Returns Value as ShapeAspectRelationship (or Null if another type)

end RepresentedDefinition;
