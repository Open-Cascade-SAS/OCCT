-- Created on: 1994-09-02
-- Created by: Christian CAILLET
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SelectIncorrectEntities  from IFSelect  inherits SelectFlag

    ---Purpose : A SelectIncorrectEntities sorts the Entities which have been
    --           noted as Incorrect in the Graph of the Session
    --             (flag "Incorrect")
    --           It can find a result only if ComputeCheck has formerly been
    --           called on the WorkSession. Else, its result will be empty.

uses AsciiString from TCollection, InterfaceModel, Graph, EntityIterator

is

    Create returns mutable SelectIncorrectEntities;
    ---Purpose : Creates a SelectIncorrectEntities
    --           i.e. a SelectFlag("Incorrect")

end SelectIncorrectEntities;
