-- File:	RWStepAP203_RWCcDesignPersonAndOrganizationAssignment.cdl
-- Created:	Fri Nov 26 16:26:32 1999 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0
-- Copyright:	Matra Datavision 1999

class RWCcDesignPersonAndOrganizationAssignment from RWStepAP203

    ---Purpose: Read & Write tool for CcDesignPersonAndOrganizationAssignment

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    CcDesignPersonAndOrganizationAssignment from StepAP203

is
    Create returns RWCcDesignPersonAndOrganizationAssignment from RWStepAP203;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : CcDesignPersonAndOrganizationAssignment from StepAP203);
	---Purpose: Reads CcDesignPersonAndOrganizationAssignment

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: CcDesignPersonAndOrganizationAssignment from StepAP203);
	---Purpose: Writes CcDesignPersonAndOrganizationAssignment

    Share (me; ent : CcDesignPersonAndOrganizationAssignment from StepAP203;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWCcDesignPersonAndOrganizationAssignment;
