-- Created on: 1991-04-22
-- Created by: jean pierre TIRAULT
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

generic class Hash from PCollection (key as Storable) inherits Storable
    is
    
    
    
    Create returns Hash;
    ---Purpose : Empty constructor.



    HashCode (me; MyKey : key ; Upper : Integer) 
             returns Integer is virtual;
    ---Level: Public
    ---Purpose: Returns a hashcod value of key bounded by Upper.



    Compare (me; One , Two : key) returns Boolean is virtual;    
    ---Level: Public
    ---Purpose : Compare two keys and returns a boolean value

end;

