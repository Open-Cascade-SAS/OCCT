-- Created on: 1993-09-28
-- Created by: Denis PASCAL
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class TSNode from GraphTools 

uses SequenceOfInteger from TColStd

is

    Create returns TSNode from GraphTools;
    
    Reset (me : in out);

    IncreaseRef  (me : in out);

    DecreaseRef  (me : in out);

    NbRef        (me) returns Integer from Standard;

    AddSuccessor (me : in out; s : Integer from Standard);

    NbSuccessors (me) returns Integer from Standard;

    GetSuccessor (me; index : Integer from Standard)
    returns Integer from Standard;

fields

    referenceCount : Integer from Standard;
    mySuccessors   : SequenceOfInteger from TColStd;

end TSNode;




