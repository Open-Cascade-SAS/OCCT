-- Created on: 1997-04-29
-- Created by: Alexander BRIVIN
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DeflectionCurve from VrmlConverter 

    	---Purpose: DeflectionCurve    -  computes the presentation of
    	--          objects to be seen as  curves,   converts this  one into
    	--          VRML    objects    and    writes (adds)  into
    	--          anOStream.     All  requested properties  of   the
    	--          representation  are specify in  aDrawer.   
	--          This  kind of the presentation
    	--          is converted into IndexedLineSet ( VRML ).
        --          The computation will be made according to a maximal
        --          chordial deviation. 

uses
 
    Length       from Quantity,
    Curve        from Adaptor3d,
    Drawer       from VrmlConverter

is

    Add(myclass; anOStream: in out OStream from Standard; 
    	    	 aCurve       : in out Curve        from Adaptor3d;
    	    	 aDrawer      : Drawer       from VrmlConverter);

    ---Purpose: adds to the OStream the drawing of the curve aCurve with  
    --          respect to the maximal chordial deviation defined
    --          by the drawer aDrawer.
    --          The aspect is defined by LineAspect in aDrawer.
    --          

 
    Add(myclass; anOStream: in out OStream from Standard; 
    	    	 aCurve       : in out Curve        from Adaptor3d;
                 U1, U2       : Real         from Standard;
    	    	 aDrawer      : Drawer       from VrmlConverter);
		    
    ---Purpose: adds to the OStream the drawing of the curve aCurve with  
    --          respect to the maximal chordial deviation defined
    --          by the drawer aDrawer.
    --          The aspect is defined by LineAspect in aDrawer.
    --          The drawing will be limited between the points of parameter
    --          U1 and U2.


    Add(myclass; anOStream: in out OStream from Standard; 
    	    	 aCurve       : in out Curve        from Adaptor3d;
    	    	 aDeflection  : Real         from Standard;
    	    	 aLimit       : Real         from Standard);

    ---Purpose: adds to the OStream the drawing of the curve aCurve with  
    --          respect to the maximal chordial deviation aDeflection.
    --          The aspect is the current aspect


    Add(myclass; anOStream:  in out OStream from Standard;
    	    	 aCurve       : in out Curve        from Adaptor3d;
    	    	 aDeflection  : Real         from Standard;
    	    	 aDrawer      : Drawer       from VrmlConverter);

    ---Purpose: adds to the OStream the drawing of the curve aCurve with  
    --          respect to the maximal chordial deviation aDeflection.
    --          The aspect is the current aspect


    Add(myclass; anOStream: in out OStream from Standard; 
    	    	 aCurve       : in out Curve        from Adaptor3d;
                 U1, U2       : Real         from Standard;
    	    	 aDeflection  : Real         from Standard);
		 
    ---Purpose: adds to the OStream the drawing of the curve aCurve with  
    --          respect to the maximal chordial deviation aDeflection.
    --          The aspect is the current aspect
    --          The drawing will be limited between the points of parameter
    --          U1 and U2.


end DeflectionCurve;
