-- Created on: 1995-03-24
-- Created by: Robert COUBLANC
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SensitiveFace from Select3D 
inherits SensitivePoly from Select3D

    ---Purpose: Sensitive Entity to make a face selectable.
    -- In some cases this class can raise Standard_ConstructionError and 
    -- Standard_OutOfRange exceptions. For more details see Select3D_SensitivePoly.

uses
    EntityOwner       from SelectBasics,
    Projector         from Select3D,
    Lin               from gp,
    ListOfBox2d       from SelectBasics,
    PickArgs          from SelectBasics,
    Array1OfPnt       from TColgp,
    HArray1OfPnt      from TColgp,
    Array1OfPnt2d     from TColgp,
    Box2d             from Bnd,
    TypeOfSensitivity from Select3D,
    Location          from TopLoc, 
    SensitiveEntity   from Select3D

raises
    ConstructionError from Standard,
    OutOfRange from Standard

is

    Create (OwnerId      : EntityOwner from SelectBasics;
            ThePoints    : Array1OfPnt from TColgp;
            Sensitivity  : TypeOfSensitivity = Select3D_TOS_INTERIOR)
     returns mutable SensitiveFace;
        ---Level: Public 
        ---Purpose: Constructs a sensitive face object defined by the
        -- owner OwnerId, the array of points ThePoints, and
        -- the sensitivity type Sensitivity.
        -- The array of points is the outer polygon of the geometric face.

    Create (OwnerId      : EntityOwner from SelectBasics;
            ThePoints    : HArray1OfPnt from TColgp;
            Sensitivity  : TypeOfSensitivity = Select3D_TOS_INTERIOR)
     returns mutable SensitiveFace;
        ---Level: Public 
        ---Purpose: Constructs a sensitive face object defined by the
        -- owner OwnerId, the array of points ThePoints, and
        -- the sensitivity type Sensitivity.
        -- The array of points is the outer polygon of the geometric face.
   
    Matches (me : mutable;
             thePickArgs : PickArgs from SelectBasics;
             theMatchDMin, theMatchDepth : out Real from Standard)
    returns Boolean is redefined virtual;
    ---Level: Public
    ---Purpose: Checks whether the sensitive entity matches the picking
    -- detection area (close to the picking line).
    -- For details please refer to base class declaration.

    Matches (me  :mutable; 
             XMin,YMin,XMax,YMax : Real from Standard;
             aTol: Real from Standard) 
    returns Boolean
    is redefined virtual;
    ---Level: Public 
     
    Matches (me  :mutable; 
             Polyline:Array1OfPnt2d from TColgp;
             aBox:Box2d from Bnd;
             aTol: Real from Standard) 
    returns Boolean
    is redefined virtual;
    ---Level: Public 
    

    ComputeDepth (me;
                  thePickLine : Lin from gp;
                  theDepthMin, theDepthMax : Real from Standard)
    returns Real from Standard
    is virtual;
    ---Level: Public
    ---Purpose: Computes the depth values for all 3D points defining this face and returns
    -- the minimal value among them.
    -- If the "minimal depth" approach is not suitable and gives wrong detection results
    -- in some particular case, a custom sensitive face class can redefine this method.

    ComputeDepth(me;EyeLine: Lin from gp)
    is private;
    ---Level: Public
    ---Purpose: Warning: Obsolete.
    -- Use newer version of the method with min, max limits passed as arguments.

    Dump(me; S: in out OStream;FullDump : Boolean from Standard = Standard_True) is redefined virtual; 

    GetConnected(me: mutable; theLocation : Location from TopLoc) 
    returns SensitiveEntity from Select3D 
    is redefined virtual; 
        ---Level: Public 
        ---Purpose: Returns the copy of this


fields

    mytype          : TypeOfSensitivity;
end SensitiveFace;
