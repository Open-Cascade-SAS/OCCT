-- File:        CurveStyle.cdl
-- Created:     Mon Dec  4 12:02:25 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWCurveStyle from RWStepVisual

	---Purpose : Read & Write Module for CurveStyle

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     CurveStyle from StepVisual,
     EntityIterator from Interface

is

	Create returns RWCurveStyle;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable CurveStyle from StepVisual);

	WriteStep (me; SW : in out StepWriter; ent : CurveStyle from StepVisual);

	Share(me; ent : CurveStyle from StepVisual; iter : in out EntityIterator);

end RWCurveStyle;
