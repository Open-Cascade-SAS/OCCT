-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class RepresentationContext from StepRepr 

inherits TShared from MMgt

uses

	HAsciiString from TCollection
is

	Create returns RepresentationContext;
	---Purpose: Returns a RepresentationContext

	Init (me : mutable;
	      aContextIdentifier : HAsciiString from TCollection;
	      aContextType : HAsciiString from TCollection) is virtual;

	-- Specific Methods for Field Data Access --

	SetContextIdentifier(me : mutable; aContextIdentifier : HAsciiString);
	ContextIdentifier (me) returns HAsciiString;
	SetContextType(me : mutable; aContextType : HAsciiString);
	ContextType (me) returns HAsciiString;

fields

	contextIdentifier : HAsciiString from TCollection;
	contextType : HAsciiString from TCollection;

end RepresentationContext;
