-- Created on: 2002-10-29
-- Created by: Michael SAZONOV
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ADriverTable from BinMDF inherits TShared from MMgt

        ---Purpose: A driver table is an object building links between
        --          object types and object drivers. In the
        --          translation process, a driver table is asked to
        --          give a translation driver for each current object
        --          to be translated.

uses
    Type               from Standard,
    ADriver            from BinMDF,    
    TypeADriverMap     from BinMDF,
    IndexedMapOfTransient from TColStd,
    SequenceOfAsciiString from TColStd,
    TypeIdMap from BinMDF

is
    Create returns mutable ADriverTable from BinMDF;
        ---Purpose: Constructor

    AddDriver(me : mutable; theDriver : ADriver from BinMDF);
        ---Purpose: Adds a translation driver <theDriver>.

    AssignId(me : mutable; theType	: Type from Standard;
			   theId	: Integer from Standard)
    	is private;
	---C++: inline
        ---Purpose: Assigns the ID to the driver of the Type

    AssignIds(me : mutable; theTypes	: IndexedMapOfTransient from TColStd);
        ---Purpose: Assigns the IDs to the drivers of the given Types.
        --          It uses indices in the map as IDs.
        --          Useful in storage procedure.

    AssignIds(me : mutable; theTypeNames : SequenceOfAsciiString from TColStd);
        ---Purpose: Assigns the IDs to the drivers of the given Type Names;
        --          It uses indices in the sequence as IDs.
        --          Useful in retrieval procedure.

    GetDriver(me; theType     : Type from Standard;
                  theDriver   : in out ADriver from BinMDF)
        returns Integer from Standard;
	---C++: inline
        ---Purpose: Gets a driver <theDriver> according to <theType>.
        --          Returns Type ID if the driver was assigned an ID; 0 otherwise.

    GetDriver(me; theTypeId   : Integer from Standard)
    	returns ADriver from BinMDF;
	---C++: inline
        ---Purpose: Returns a driver according to <theTypeId>.
        --          Returns null handle if a driver is not found

fields
    myMap	: TypeADriverMap from BinMDF;
    myMapId	: TypeIdMap from BinMDF;

end ADriverTable;
