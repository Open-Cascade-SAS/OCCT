-- Created on: 1997-06-10
-- Created by: Yves FRICAUD
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



private class Localizer from TNaming 

	---Purpose: 

uses
    Shape                                  from TopoDS,
    ShapeEnum                              from TopAbs,
    Label                                  from TDF,
    LabelList                              from TDF,
    LabelMap                               from TDF,
    UsedShapes                             from TNaming,
    NamedShape                             from TNaming,
    MapOfNamedShape                        from TNaming,
    ListOfNamedShape                       from TNaming,
    Evolution                              from TNaming,
    ShapesSet                              from TNaming,	
    ListOfShape                            from TopTools,
    MapOfShape                             from TopTools,
    IndexedDataMapOfShapeListOfShape       from TopTools,
    ListOfMapOfShape                       from TNaming,
    ListOfIndexedDataMapOfShapeListOfShape from TNaming
	    
is


    Create returns Localizer from TNaming;
    
    Init (me       : in out;
    	  US       : UsedShapes from TNaming;
	  CurTrans : Integer    from Standard );

    SubShapes (me : in out; S : Shape from TopoDS; Type : ShapeEnum from TopAbs) 
    returns MapOfShape from TopTools;
    ---C++: return const&
  
    Ancestors    (me : in out; S : Shape from TopoDS; Type : ShapeEnum from TopAbs)
    returns IndexedDataMapOfShapeListOfShape from TopTools;
    ---C++: return const&
    
    FindFeaturesInAncestors (me            : in out;
    	    	    	     S             :        Shape      from TopoDS;
			     In            :        Shape      from TopoDS;
			     AncInFeatures : in out MapOfShape from TopTools);
			     
			     
    GoBack (me     : in out;
    	    S      : Shape                   from TopoDS;
	    Lab    : Label                   from TDF;
	    Evol   : Evolution               from TNaming;
	    OldS   : in out ListOfShape      from TopTools;
	    OldLab : in out ListOfNamedShape from TNaming);
	    

    Backward (me          : in out;
    	      NS          :        NamedShape      from TNaming;
    	      S           :        Shape           from TopoDS;
	      Primitives  : in out MapOfNamedShape from TNaming;
	      ValidShapes : in out MapOfShape      from TopTools);
	      
    FindNeighbourg (me         : in out;
    	            Cont       :       Shape from TopoDS;
		    S          :       Shape from TopoDS;
		    Neighbourg : in out MapOfShape from TopTools);
		    	
    IsNew (myclass ;S  : Shape      from TopoDS;
    	            NS : NamedShape from TNaming)
    returns Boolean from Standard;
    
    FindGenerator (myclass ; NS :        NamedShape from TNaming;
	    		     S  :        Shape      from TopoDS;
    	    theListOfGenerators : in out ListOfShape from TopTools );

    
    FindShapeContext (myclass ; NS    :        NamedShape from TNaming;
    	    	    	    	theS  :        Shape      from TopoDS; 
				theSC : in out Shape      from TopoDS); 
    ---Purpose: Finds context of the shape <S>.		    				

fields

    myCurTrans           : Integer                                from Standard;	
    myUS                 : UsedShapes                             from TNaming;

    myShapeWithSubShapes : ListOfShape                            from TopTools;
    mySubShapes          : ListOfMapOfShape                       from TNaming;
    
    myShapeWithAncestors : ListOfShape                            from TopTools;
    myAncestors          : ListOfIndexedDataMapOfShapeListOfShape from TNaming;
    
end Localizer;









