-- Created on: 1993-04-26
-- Created by: Jean-Louis Frenkel
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

--   GG  : GER61351 17/11/1999 Change SetColor() with a compatible Quantity_Color instead
--				       the restricted NameOfColor.


class IsoAspect from Prs3d inherits LineAspect from Prs3d
    	---Purpose: A framework to define the display attributes of isoparameters.
    	-- This framework can be used to modify the default
    	-- setting for isoparameters in AIS_Drawer.
        
uses 

    NameOfColor from Quantity,
    Color from Quantity,
    TypeOfLine from Aspect

is
    Create (aColor: NameOfColor from Quantity;
	    aType: TypeOfLine from Aspect;
    	    aWidth: Real from Standard;
          aNumber: Integer from Standard)    
	    returns mutable IsoAspect from Prs3d;
    	---Purpose: Constructs a framework to define display attributes of isoparameters.
    	-- These include:
    	-- -   the color attribute aColor
    	-- -   the type of line aType
    	-- -   the width value aWidth
    	-- -   aNumber, the number of isoparameters to be   displayed.
        
    Create (aColor: Color from Quantity;
	    aType: TypeOfLine from Aspect;
    	    aWidth: Real from Standard;
          aNumber: Integer from Standard)	    
	    returns mutable IsoAspect from Prs3d;
	    

    SetNumber (me: mutable; aNumber: Integer from Standard) 
    	---Purpose: defines the number of U or V isoparametric curves 
    	--         to be drawn for a single face.
    	--          Default value: 10
    is static;

    Number (me) returns Integer from Standard 
    	---Purpose: returns the number of U or V isoparametric curves drawn for a single face.
    is static;
    
fields

    myNumber: Integer from Standard;
    
end IsoAspect from Prs3d;
