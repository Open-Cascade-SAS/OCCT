-- Created on: 1999-03-24
-- Created by: data exchange team
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class AssemblyExplorer from STEPSelections 

	---Purpose: 

uses
    
    Graph from Interface,
    SequenceOfAssemblyComponent        from STEPSelections,
    IndexedDataMapOfTransientTransient from TColStd,
    ProductDefinition                  from StepBasic,
    ShapeDefinitionRepresentation      from StepShape,
    AssemblyComponent                  from STEPSelections,
    NextAssemblyUsageOccurrence        from StepRepr
    
is
    
    Create (G: Graph) returns AssemblyExplorer from STEPSelections;
    
    Init(me: in out; G: Graph);
    
    Dump(me; os: in out OStream from Standard);
    
    FindSDRWithProduct(me; product: ProductDefinition from StepBasic)
    returns ShapeDefinitionRepresentation from StepShape;
    
    FillListWithGraph(me: in out; cmp: AssemblyComponent from STEPSelections);
    
    FindItemWithNAUO(me; nauo: NextAssemblyUsageOccurrence from StepRepr)
    returns Transient from Standard;
    
    --Methods for fetching the results
    
    NbAssemblies(me) returns Integer;
    	---Purpose: Returns the number of root assemblies;
	---C++: inline
    
    Root(me; rank: Integer = 1) returns AssemblyComponent from STEPSelections;
    	---Purpose: Returns root of assenbly by its rank;
	---C++: inline
    

fields

    myRoots: SequenceOfAssemblyComponent from STEPSelections;
    myGraph: Graph from Interface;
    myMap  : IndexedDataMapOfTransientTransient from TColStd;    

end AssemblyExplorer;
