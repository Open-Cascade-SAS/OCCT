-- Created on: 1997-06-26
-- Created by: Laurent PAINNOT
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

private class Classifier from BRepMesh



uses  
    Pnt2d                         from gp,
    SequenceOfPnt2d               from TColgp,
    Face                          from TopoDS,
    State                         from TopAbs,
    SequenceOfInteger             from TColStd,
    SeqOfPtr                      from BRepTopAdaptor, 
    DataMapOfShapePairOfPolygon   from BRepMesh,
    IndexedMapOfInteger           from TColStd,
    IndexedMapOfVertex            from BRepMesh,
    Status                        from BRepMesh,
    DataStructureOfDelaun         from BRepMesh

is 
    
    Create   (theFace      : Face                          from TopoDS; 
              theTolUV     : Real                          from Standard;
              theEdges     : DataMapOfShapePairOfPolygon   from BRepMesh;
              theMap       : IndexedMapOfInteger           from TColStd;
              theStructure : DataStructureOfDelaun         from BRepMesh;
              theUmin, theUmax, theVmin, theVmax : Real    from Standard)
    returns Classifier from BRepMesh;


    Perform(me; thePoint: Pnt2d from gp)
    returns State from TopAbs;


    State (me)
    returns Status from BRepMesh;
        ---C++: inline


    Destroy(me: in out);
        ---C++: alias ~


    AnalizeWire (me          : in out;
                 theSeqPnt2d : in SequenceOfPnt2d from TColgp;
                 theUmin, theUmax, theVmin, theVmax: in Real from Standard)
    is private;
    -- Private method called from constructor after some (piece of) wire 
    -- has been explored and put into <theSeqPnt2d>. 
    -- Here it is triangulated if it is a hole and anyway added to the bulk.
    
fields 

    myTabClass  : SeqOfPtr          from BRepTopAdaptor;
    myTabOrient : SequenceOfInteger from TColStd;
    myTolUV     : Real              from Standard;
    myFace      : Face              from TopoDS;
    myState     : Status            from BRepMesh;

end Classifier from BRepMesh;
