-- Created on: 1991-11-18
-- Created by: Remi GILET
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

generic class ParGenCurve from GccGeo (TheCurve as any)

    ---Purpose: Definition of a virtual curve.

uses Pnt2d  from gp,
     Vec2d  from gp
     
is

Create returns ParGenCurve;

Create(C : TheCurve) returns ParGenCurve;

Create(C : TheCurve               ;
       D : Real     from Standard ) returns ParGenCurve;

Value(me; U : Real)returns Pnt2d;
    --- Purpose : Computes the point of parameter U on the curve 

D1 (me; U : Real; P : out Pnt2d from gp ; V : out Vec2d from gp);
    --- Purpose : Computes the point of parameter U on the curve with its
    --  first derivative.

D2 (me; U : Real; P : out Pnt2d from gp ; V1,V2 : out Vec2d from gp);
    --- Purpose : Computes the point of parameter U on the curve with its
    --  first derivative and second derivative.


FirstParameter(me)  returns Real;
    	
LastParameter(me) returns Real;

GetResolution(me) returns Real;

GetIntervals(me) returns Integer;

fields

Cu  : TheCurve              ;
Dep : Real     from Standard;

end ParGenCurve;
