-- Created on: 1995-04-06
-- Created by: Jean-Louis Frenkel
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


deferred class Viewer from Viewer inherits TShared from MMgt

uses
    AsciiString,ExtendedString from TCollection,
    GraphicDriver from Graphic3d
    
is
    Initialize( aDriver: GraphicDriver from Graphic3d;
                aName: ExtString from Standard;
                aDomain: CString from Standard;
                aNextCount: Integer from Standard);
    
    Update(me: mutable) is deferred;


    Driver(me) returns mutable GraphicDriver from Graphic3d
    is static;
    ---C++: return const &
    
    NextName(me) returns ExtString from Standard
    is static;

    Domain(me) returns CString from  Standard
    is static;

    IncrCount(me:mutable) is static protected;
    
fields
    	myNextCount: Integer from Standard;
        myDomain: AsciiString from TCollection;    
        myName: ExtendedString from TCollection;
        myDriver: GraphicDriver from Graphic3d;
end Viewer  from Viewer;
