-- Created on: 1998-09-01
-- Created by: Stephanie HUMEAU
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ACRLaw from BRepFill inherits LocationLaw  from  BRepFill 

	---Purpose: Build Location Law,  with a Wire.   In the case 
	--          of guided contour and trihedron by reduced
	--          curvilinear abscissa
	       
       

uses
  Wire  from  TopoDS,
  LocationLaw from GeomFill, 
  LocationGuide from GeomFill, 
  HArray1OfReal from TColStd

is 
    Create (Path   :  Wire  from  TopoDS;  
            Law    : LocationGuide from GeomFill)  
    returns ACRLaw from BRepFill; 
    
fields 
     OrigParam  : HArray1OfReal  from TColStd; 
 
end ACRLaw;
