-- File:        Placement.cdl
-- Created:     Mon Dec  4 12:02:28 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWPlacement from RWStepGeom

	---Purpose : Read & Write Module for Placement

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     Placement from StepGeom,
     EntityIterator from Interface

is

	Create returns RWPlacement;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable Placement from StepGeom);

	WriteStep (me; SW : in out StepWriter; ent : Placement from StepGeom);

	Share(me; ent : Placement from StepGeom; iter : in out EntityIterator);

end RWPlacement;
