-- Created by: CAL
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

--              11/97 ; CAL : retrait des DataStructure

deferred class DataStructureManager from Graphic3d inherits TShared

	---Version:

	---Purpose:	This class allows the definition of a manager to
	--		which the graphic objects are associated.
	--		It allows them to be globally manipulated.
	--		It defines the global attributes.

	---Keywords:

	---Warning:
	---References:

is
	-------------------------
	-- Category: Constructors
	-------------------------

	Initialize;
	---Level: Public
	---Purpose: Initializes the manager <me>.
	---Category: Constructors

	------------------------
	-- Category: Destructors
	------------------------

	Destroy (me: mutable)
		is virtual;
	---Level: Public
	---Purpose: Deletes the manager <me>.
	---C++: alias ~
	---Category: Destructors

end DataStructureManager from Graphic3d;
