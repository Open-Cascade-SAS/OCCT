-- Created on: 1995-07-02
-- Created by: Laurent BUCHARD
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

generic class HContToolGen from Contap  (
     TheHVertex      as any;
     TheHCurve2d     as any;
     TheHSurface     as any;
     TheHCurve2dTool as any;
     TheHSurfaceTool as any)

	---Purpose: Tool for the intersection between 2 surfaces.
	--          Regroupe pour l instant les methodes hors Adaptor3d...



uses 
     Pnt2d    from gp,
     Pnt      from gp

is


    NbSamplesU(myclass; S: TheHSurface; u1,u2: Real from Standard)
        returns Integer from Standard;

    NbSamplesV(myclass; S: TheHSurface; v1,v2: Real from Standard)
        returns Integer from Standard;

-- Methodes pour recherche des points interieurs

    NbSamplePoints(myclass; S: TheHSurface)

    	returns Integer from Standard;


    SamplePoint(myclass; S    : TheHSurface;
    	    	         Index: Integer from Standard;
                         U,V: out Real from Standard);


-- Methodes sur un arc de restriction

    HasBeenSeen(myclass; C: TheHCurve2d)

	---Purpose: Returns True if all the intersection point and edges
	--          are known on the Arc.
	--          The intersection point are given as vertices.
	--          The intersection edges are given as intervals between
	--          two vertices.

    	returns Boolean from Standard;

    NbSamplesOnArc(myclass; A: TheHCurve2d)
    
    	---Purpose: returns the number of points which is used to make 
    	--          a sample on the arc. this number is a function of
    	--          the Surface and the CurveOnSurface complexity.
    
        returns Integer from Standard;


    Bounds(myclass; C: TheHCurve2d; 
                    Ufirst,Ulast: out Real from Standard);

	---Purpose: Returns the parametric limits on the arc C.
	--          These limits must be finite : they are either
	--          the real limits of the arc, for a finite arc,
	--          or a bounding box for an infinite arc.


    Project(myclass; C: TheHCurve2d;
                     P: Pnt2d from gp;
                     Paramproj: out Real from Standard;
                     Ptproj   : out Pnt2d from gp)

	---Purpose: Projects the point P on the arc C.
	--          If the methods returns Standard_True, the projection is
	--          successful, and Paramproj is the parameter on the arc
	--          of the projected point, Ptproj is the projected Point.
	--          If the method returns Standard_False, Param proj and Ptproj
	--          are not significant.
	--          

	returns Boolean from Standard;


-- Methods on a vertex


    Tolerance(myclass; V: TheHVertex; C: TheHCurve2d)

	---Purpose: Returns the parametric tolerance used to consider
	--          that the vertex and another point meet, i-e
	--          if Abs(parameter(Vertex) - parameter(OtherPnt))<=
	--          Tolerance, the points are "merged".

    	returns Real from Standard;


    Parameter(myclass; V: TheHVertex; C: TheHCurve2d)
    
	---Purpose: Returns the parameter of the vertex V on the arc A.

	returns Real from Standard;


-- The following methods are used when HasBeenSeen returns Standard_True

    NbPoints(myclass; C: TheHCurve2d)
    
	---Purpose: Returns the number of intersection points on the arc A.
    
    	returns Integer from Standard;


    Value(myclass; C: TheHCurve2d; Index: Integer from Standard;
                   Pt: out Pnt from gp; Tol: out Real from Standard;
                   U: out Real from Standard);

	---Purpose: Returns the value (Pt), the tolerance (Tol), and
	--          the parameter (U) on the arc A , of the intersection
	--          point of range Index.


    IsVertex(myclass; C: TheHCurve2d;
                      Index: Integer from Standard)
    
	---Purpose: Returns True if the intersection point of range Index
	--          corresponds with a vertex on the arc A.

    	returns Boolean from Standard;


    Vertex(myclass; C: TheHCurve2d; Index: Integer from Standard;
                    V: out TheHVertex);

	---Purpose: When IsVertex returns True, this method returns the
	--          vertex on the arc A.


    NbSegments(myclass; C: TheHCurve2d)
    
	---Purpose: returns the number of part of A solution of the
	--          of intersection problem.
    
    	returns Integer from Standard;


    HasFirstPoint(myclass; C: TheHCurve2d; 
                           Index: Integer from Standard;
                           IndFirst: out Integer from Standard)
    
	---Purpose: Returns True when the segment of range Index is not
	--          open at the left side. In that case, IndFirst is the
	--          range in the list intersection points (see NbPoints)
	--          of the one which defines the left bound of the segment.
	--          Otherwise, the method has to return False, and IndFirst
	--          has no meaning.

    	returns Boolean from Standard;


    HasLastPoint(myclass; C: TheHCurve2d;
                          Index: Integer from Standard;
                          IndLast: out Integer from Standard)
    
	---Purpose: Returns True when the segment of range Index is not
	--          open at the right side. In that case, IndLast is the
	--          range in the list intersection points (see NbPoints)
	--          of the one which defines the right bound of the segment.
	--          Otherwise, the method has to return False, and IndLast
	--          has no meaning.

    	returns Boolean from Standard;


    IsAllSolution(myclass; C: TheHCurve2d)
    
	---Purpose: Returns True when the whole restriction is solution
	--          of the intersection problem.
    
    	returns Boolean from Standard;


end HContToolGen;
