-- File:        BRepMesh.cdl
-- Created:     Wed Sep 22 17:34:57 1993
-- Author:      Didier PIFFAULT
--              <dpf@zerox>
---Copyright:    Matra Datavision 1993, 1994
 

package BRepMesh

        ---Purpose: Instantiated   package for the   class of packages

        ---Level : Advanced.  
        --  All methods of all  classes will be advanced.


uses    Standard,
        gp,
        Bnd,
        TColStd,
        TColgp,
        GCPnts,
        BRepAdaptor,
        BRepTopAdaptor,
        TCollection,
        MMgt,
        TopoDS,
        TopAbs,
        TopExp,
        TopTools,
        Poly,
        Geom2d,
        GeomAbs,
        GeomAdaptor,
        TopLoc,
        SortTools


is    enumeration DegreeOfFreedom is 
        Free,
        InVolume,
        OnSurface,
        OnCurve,
        Fixed,
        Frontier,
        Deleted;

      enumeration Status  is 
      ---Purpose: Discribes the wires discretisation.
        NoError,
        OpenWire,
        SelfIntersectingWire,
        Failure,
        ReMesh
      end Status;
       
      enumeration FactoryError is 
        FE_NOERROR,  
        FE_LIBRARYNOTFOUND,
        FE_FUNCTIONNOTFOUND,
        FE_CANNOTCREATEALGO
      end FactoryError;   
      
      class Vertex;

      class Edge;

      class Triangle;

      class ShapeTool;

      class Circ;

      deferred class DiscretRoot; 
      class DiscretFactory;
      --
      pointer PDiscretRoot to DiscretRoot from BRepMesh;
      --
      imported MapOfIntegerInteger from BRepMesh;
      imported MapOfInteger from BRepMesh;
      imported ListOfInteger from BRepMesh;
      imported BaseAllocator from BRepMesh;
      imported PairOfIndex from BRepMesh;
      imported CircleInspector from BRepMesh;
      imported CellFilter from BRepMesh;

      class ComparatorOfVertexOfDelaun;
      class ComparatorOfIndexedVertexOfDelaun;
      class SelectorOfDataStructureOfDelaun;
      class Delaun;
      class DataStructureOfDelaun;
      class CircleTool;

      class Array1OfVertexOfDelaun instantiates Array1 from TCollection
        (Vertex from BRepMesh);

      class HArray1OfVertexOfDelaun instantiates HArray1 from TCollection
        (Vertex from BRepMesh, Array1OfVertexOfDelaun);

      class HeapSortVertexOfDelaun instantiates  HeapSort from SortTools
        (Vertex from BRepMesh, Array1OfVertexOfDelaun,
        ComparatorOfVertexOfDelaun from BRepMesh);

      class HeapSortIndexedVertexOfDelaun instantiates  HeapSort from SortTools
        (Integer, Array1OfInteger from TColStd,
        ComparatorOfIndexedVertexOfDelaun from BRepMesh);

      class NodeHasherOfDataStructureOfDelaun instantiates MapHasher from TCollection
        (Vertex from BRepMesh);
      class LinkHasherOfDataStructureOfDelaun instantiates MapHasher from TCollection
        (Edge from BRepMesh);
      class ElemHasherOfDataStructureOfDelaun instantiates MapHasher from TCollection
        (Triangle from BRepMesh);

      class IDMapOfNodeOfDataStructureOfDelaun  instantiates IndexedDataMap from TCollection
        (Vertex from BRepMesh,
        ListOfInteger from BRepMesh,
        NodeHasherOfDataStructureOfDelaun);

      class IDMapOfLinkOfDataStructureOfDelaun  instantiates IndexedDataMap from TCollection
        (Edge from BRepMesh,
        PairOfIndex from BRepMesh,
        LinkHasherOfDataStructureOfDelaun);

      class IMapOfElementOfDataStructureOfDelaun instantiates IndexedMap from TCollection
        (Triangle from BRepMesh,
        ElemHasherOfDataStructureOfDelaun);

      class DataMapOfVertexInteger instantiates DataMap from TCollection
          (Vertex from TopoDS, Integer from Standard, ShapeMapHasher from TopTools);

      class ListOfVertex instantiates List from TCollection 
          (Vertex from  BRepMesh);

        class ListOfXY instantiates List from TCollection (XY from gp);

      class DataMapOfIntegerListOfXY  instantiates DataMap from TCollection
          (Integer from Standard, ListOfXY from BRepMesh, MapIntegerHasher from TColStd);


      class  VertexHasher  instantiates   MapHasher  from  TCollection(Vertex  from  BRepMesh);

      class IndexedMapOfVertex instantiates IndexedMap from TCollection 
          (Vertex from  BRepMesh,  VertexHasher from  BRepMesh);


      class DataMapOfShapeReal instantiates DataMap from TCollection
                                            (Shape          from TopoDS,
                                             Real           from Standard,
                                             ShapeMapHasher from TopTools);

      class BiPoint;
  
      class Array1OfBiPoint    instantiates Array1  from TCollection(BiPoint from BRepMesh);

      private class FastDiscretFace;
      
      class FastDiscret;
      
      class FaceAttribute;
  
      class DataMapOfFaceAttribute instantiates DataMap from TCollection
                                            (Face           from TopoDS,
                                             FaceAttribute  from BRepMesh,
                                             ShapeMapHasher from TopTools);
              
      private class Classifier;
      imported ClassifierPtr; -- smart pointer on Classifier

      class IncrementalMesh from BRepMesh;
      ---Purpose: meshes faces from a Shape only if necessary.

         ---- classes moved from MeshShape
      class GeomTool;

      class DataMapOfIntegerPnt instantiates
          DataMap from TCollection   (Integer          from Standard,
                                      Pnt              from gp,
                                      MapIntegerHasher from TColStd);

      class PairOfPolygon;

      class DataMapOfShapePairOfPolygon instantiates 
      DataMap from TCollection(Shape          from TopoDS,
                               PairOfPolygon  from BRepMesh,
                               ShapeMapHasher from TopTools);

      Mesh(S: Shape from TopoDS; d: Real from Standard);
      ---Purpose: call to incremental mesh.

  
end BRepMesh;
