-- Created on: 1993-09-07
-- Created by: GG
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class FontMap from Aspect inherits TShared from MMgt

	---Version: 0.0

	---Purpose: This class defines a FontMap object.
	---Keywords:
	---Warning:
	---References:
uses
	FontStyle		from Aspect,
	FontMapEntry 		from Aspect,
	SequenceOfFontMapEntry 	from Aspect

raises
	BadAccess 	from Aspect

is

	Create returns mutable FontMap from Aspect;

        AddEntry (me : mutable; AnEntry : FontMapEntry from Aspect)
	---Level: Public
        ---Purpose: Adds an entry in the font map <me>.
        --  Warning: Raises BadAccess if FontMap size is exceeded.
        raises BadAccess from Aspect;

        AddEntry (me : mutable; aStyle : FontStyle from Aspect)
                                        returns Integer from Standard;
        ---Level: Public
        ---Purpose: Search an identical font style entry in the font map <me>
        -- and returns the FontMapEntry Index if exist.
        -- Or add a new entry and returns the computed FontMapEntry index used.

        Size( me ) returns Integer from Standard is static;
        ---Level: Public
        ---Purpose: Returns the Allocated fontmap Size
 
        Index( me ; aFontmapIndex : Integer ) returns Integer from Standard
        ---Level: Public
        ---Purpose: Returns the FontMapEntry.Index of the FontMap
        --          at rank <aFontmapIndex> .
        raises BadAccess from Aspect is static;
        ---Trigger: Raises BadAccess if the index less than 1 or
        --          greater than Size.

	Dump( me ) ;

	Entry ( me ;
		AnIndex : Integer from Standard )
	returns FontMapEntry from Aspect
	---Level: Public
	---Purpose: Returns the Font map entry with the index <AnIndex>.
	--  Warning: Raises BadAccess if the index less than 1
	--	    or greater than Size.
	raises BadAccess from Aspect is static;

fields

	mydata	    :	SequenceOfFontMapEntry from Aspect is protected;

end FontMap ;
