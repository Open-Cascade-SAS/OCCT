-- Created on: 1995-07-18
-- Created by: Modelistation
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class   GenExtPS from Extrema 

    	---Purpose: It calculates all the extremum distances
    	--          between a point and a surface.
    	--          These distances can be minimum or maximum.

uses  	POnSurf       from Extrema,
    	Pnt           from gp,
	FuncExtPS     from Extrema,
	Surface       from Adaptor3d,
	SurfacePtr    from Adaptor3d,
        HUBTreeOfSphere from Extrema,
        ExtFlag from Extrema,
	ExtAlgo from Extrema,
	HArray1OfSphere from Bnd,
	Vector        from math,
	HArray1OfReal from TColStd,
	POnSurfParams from Extrema,
	HArray2OfPOnSurfParams from Extrema

raises  NotDone      from StdFail,
    	OutOfRange   from Standard,
	TypeMismatch from Standard
	

is

    Create returns GenExtPS;
    
    Create (P: Pnt; S: Surface from Adaptor3d; NbU,NbV: Integer; TolU,TolV: Real; F : ExtFlag from Extrema = Extrema_ExtFlag_MINMAX; A : ExtAlgo from Extrema = Extrema_ExtAlgo_Grad)
    	returns GenExtPS;
      	---Purpose: It calculates all the distances.
        --          The function F(u,v)=distance(P,S(u,v)) has an 
        --          extremum when gradient(F)=0. The algorithm searchs
        --          all the zeros inside the definition ranges of the 
        --          surface.
      	--          NbU and NbV are used to locate the close points
      	--          to find the zeros. They must be great enough
      	--          such that if there is N extrema, there will
      	--          be N extrema between P and the grid.
      	--          TolU et TolV are used to determine the conditions 
      	--          to stop the iterations; at the iteration number n:
      	--           (Un - Un-1) < TolU and (Vn - Vn-1) < TolV .


    Create (P: Pnt; S: Surface from Adaptor3d; NbU,NbV: Integer; 
    	    Umin, Usup, Vmin, Vsup: Real; TolU,TolV: Real; F : ExtFlag from Extrema = Extrema_ExtFlag_MINMAX; A : ExtAlgo from Extrema = Extrema_ExtAlgo_Grad)
    	returns GenExtPS;
      	---Purpose: It calculates all the distances.
        --          The function F(u,v)=distance(P,S(u,v)) has an 
        --          extremum when gradient(F)=0. The algorithm searchs
        --          all the zeros inside the definition ranges of the 
        --          surface.
      	--          NbU and NbV are used to locate the close points
      	--          to find the zeros. They must be great enough
      	--          such that if there is N extrema, there will
      	--          be N extrema between P and the grid.
      	--          TolU et TolV are used to determine the conditions 
      	--          to stop the iterations; at the iteration number n:
      	--           (Un - Un-1) < TolU and (Vn - Vn-1) < TolV .

    
    Initialize(me: in out; S: Surface from Adaptor3d; NbU, NbV: Integer; TolU, TolV: Real)
    	---Pupose: sets the fields of the algorithm.
    is static;


    Initialize(me: in out; S: Surface from Adaptor3d; NbU, NbV: Integer; 
    	       Umin, Usup, Vmin, Vsup: Real; TolU, TolV: Real)
    	---Pupose: sets the fields of the algorithm.
    is static;
    

    Perform(me: in out; P: Pnt from gp)
        ---Purpose: the algorithm is done with the point P.
        --          An exception is raised if the fields have not
        --          been initialized.  
    raises TypeMismatch from Standard
    is static;
    
    SetFlag(me : in out; F : ExtFlag from Extrema)
    	is static;
	
    SetAlgo(me : in out; A : ExtAlgo from Extrema)
    	is static;


    IsDone (me) returns Boolean
    	---Purpose: Returns True if the distances are found.
    	is static;
    
    NbExt (me) returns Integer
    	---Purpose: Returns the number of extremum distances.
    	raises  NotDone from StdFail
	    	-- if IsDone(me)=False.
    	is static;

    SquareDistance (me; N: Integer) returns Real
    	---Purpose: Returns the value of the Nth resulting square distance.
    	raises  NotDone from StdFail,
    	    	-- if IsDone(me)=False.
    	        OutOfRange
		-- if N < 1 or N > NbPoints(me).
    	is static;

    Point (me; N: Integer) returns POnSurf
        ---C++: return const &
    	---Purpose: Returns the point of the Nth resulting distance.
    	raises  NotDone from StdFail,
    	    	-- if IsDone(me)=False.
    	        OutOfRange
		-- if N < 1 or N > NbPoints(me).
    	is static;

    Bidon(me) returns SurfacePtr from Adaptor3d
    is static private;
    
    BuildTree(me : in out)
    is static private;
    
    FindSolution(me: in out; P : Pnt from gp;
         theParams: POnSurfParams from Extrema)
    is static private;
    
    GetGridPoints(me: in out;  theSurf: Surface from Adaptor3d) is private;
    	---Purpose: Selection of points to build grid, depending on the type of surface
    
    BuildGrid(me: in out; thePoint: Pnt from gp) is private;
    	---Purpose: Creation of grid of parametric points

    ComputeEdgeParameters(me: in out;
                          IsUEdge    : Boolean;
                          theParam0  : POnSurfParams from Extrema;
                          theParam1  : POnSurfParams from Extrema;
                          thePoints  : Pnt from gp;
                          theDiffTol : Real) returns POnSurfParams from Extrema
    is private;
      ---Purpose: Compute new edge parameters.
      ---C++: return const &


fields
    myDone    : Boolean;
    myInit    : Boolean;
    myumin    : Real;
    myusup    : Real;
    myvmin    : Real;
    myvsup    : Real;
    myusample : Integer;
    myvsample : Integer;
    mytolu    : Real;
    mytolv    : Real;
    myPoints  : HArray2OfPOnSurfParams from Extrema;
    mySphereUBTree : HUBTreeOfSphere from Extrema;
    mySphereArray : HArray1OfSphere from Bnd;
    myF	      : FuncExtPS from Extrema;
    myS       : SurfacePtr from Adaptor3d;
    myFlag    : ExtFlag from Extrema;
    myAlgo    : ExtAlgo from Extrema;
    myUParams : HArray1OfReal from TColStd;
    myVParams : HArray1OfReal from TColStd;
    myFacePntParams  : HArray2OfPOnSurfParams from Extrema;
    myUEdgePntParams : HArray2OfPOnSurfParams from Extrema;
    myVEdgePntParams : HArray2OfPOnSurfParams from Extrema;
    myGridParam      : POnSurfParams from Extrema;

end GenExtPS;
