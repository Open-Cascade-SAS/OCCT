-- Created on: 1992-10-13
-- Created by: Ramin BARRETO
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


deferred class PManaged from PMMgt

inherits Persistent from Standard

  ---Purpose: 
  --   The class <PManaged> is a persistent abstract class that
  --   provides a strategy for managing  the necessary storage 
  --   for an instance of <PManaged>. The storage is taken from
  --   Persistent cache.
  --
  --   The storage of an instance is returned to persistent cache
  --   when the instance is deleted explicitly.
  --
  --   The persistent classes like the persistent nodes benefit from
  --   the "PManaged" allocator if they inherit from <PManaged>.
  --   
  --  Warning: 
  --    The only way to delete explicitly an instance of <PManaged> is 
  --    to apply the method "Delete()" to a "Handle(PManaged)".
  --    Exemple:
  --       Handle(PManaged) aHand ;
  --       ...
  --       aHand.Delete(); 
  --       

uses  
   Integer from Standard

raises  
    OutOfMemory from Standard
  
is
    --New(myclass; aSize: Integer) returns PManaged
    ---Purpose:
    --   Returns an instance. The storage of the given "size" is 
    --   allocated by <StorageManager>.
    --
    --raises  
    --	OutOfMemory;  
    --	-- If the allocation fails.
    -- -C++: alias "void* operator new (size_t);"
    ---Level: Advanced

    --Delete(myclass; aInstance: PManaged; aSize: Integer);
    ---Purpose: 
    --   Returns the storage of the given size to the <StorageManager>.
    --   The application using "Delete" must guarantee that the
    --   instance is not shared.
    --
    -- -C++: alias "void operator delete (void*, size_t);"
    ---Level: Advanced

    --Destructor(me);
    ---Purpose: 
    --   The virtual Destructor for the class "PManaged". This
    --   declaration is necessary for the C++ compiler to
    --   generate a call to "operator delete" with the real size
    --   of the object.
    --
    -- -C+..+: alias "virtual ~PMMgt_PManaged();"
    ---Level: Advanced
    
    Initialize ;
    
end PManaged from PMMgt;

