-- Created on: 1997-09-27
-- Created by: PCT
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Modified:	03-02-98 : FMN ; Add Flag Normal

class VertexNT from Graphic3d inherits VertexN from Graphic3d

	---Version:

	---Purpose: This class allows the creation and update of
	--	    a vertex with a 3D normal and texture coordinate.

	---Keywords: Vertex, Normal, Coordinate, Point, Texture

	---Warning:
	---References:

uses

	Vector	from Graphic3d,
	Vertex	from Graphic3d

is

	Create
		returns VertexNT from Graphic3d;
	---Level: Public
	---Purpose: Creates a point with 0.0, 0.0, 0.0 coordinates
	--	    for which the normal is 0.0, 0.0, 1.0.
	--          texture coordinate is 0.0, 0.0.

	Create ( AX, AY, AZ	: Real from Standard;
		 ANX, ANY, ANZ	: Real from Standard;
		 ATX            : Real from Standard;
		 ATY            : Real from Standard = 0.0;
		 FlagNormalise  : Boolean from Standard = Standard_True )
		returns VertexNT from Graphic3d;
	---Level: Public
	---Purpose: Creates a point with coordinates <AX>, <AY>, <AZ> and
	--	    for which the normal is <ANX>, <ANY>, <ANZ>,
	--          texture coordinate is <ATX>, <ATY>.
	--	    If <FlagNormalise> is True the normal is already normalised
	--	    Else the normal is not normalised, the graphic do it.

	Create ( APoint		: Vertex from Graphic3d;
		 AVector	: Vector from Graphic3d;
		 ATX            : Real from Standard;
		 ATY            : Real from Standard = 0.0;
		 FlagNormalise  : Boolean from Standard = Standard_True )
		returns VertexNT from Graphic3d;
	---Level: Public
	---Purpose: Creates a point in <APoint> for which the normal is <AVector>. 
        --          <ATX>, <ATY> are texture coordinate.
	--	    If <FlagNormalise> is True the normal is already normalised
	--	    Else the normal is not normalised, the graphic do it.

	---------------------------------------------------
	-- Category: Methods to modify the class definition
	---------------------------------------------------

	SetTextureCoordinate( me        : in out;
			      ATX       : Real from Standard;
			      ATY       : Real from Standard = 0.0)
		is static;
	---Level: Public
	---Purpose: Modifies the texture coordinate to the point <me>.
	---Category: Methods to modify the class definition


	----------------------------
	-- Category: Inquire methods
	----------------------------
	
	TextureCoordinate( me;
			   ATX, ATY : out Real from Standard)
		is static;
	---Level: Public
	---Purpose: Returns the texture coordinate to the point <me>.
	---Category: Inquire methods

--

fields

--
-- Class	:	Graphic3d_VertexNT
--
-- Purpose	:	Declaration of variables specific to points.
--
-- Reminder	:	A point is defined by its coordinates and its normal.

	-- the texel
	MyTX, MyTY      :       Real from Standard;

end VertexNT;
