-- Created on: 2008-04-10
-- Created by: Peter KURNEV <pkv@irinox>
-- Copyright (c) 2008-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DiscretFactory from BRepMesh

    ---Purpose:
    -- This class intended to setup / retrieve default triangulation algorithm.
    -- Use BRepMesh_DiscretFactory::Get() static method to retrieve global Factory instance.
    -- Use BRepMesh_DiscretFactory::Discret() method to retrieve meshing tool.

uses
    DiscretRoot      from BRepMesh,
    FactoryError     from BRepMesh,
    PluginEntryType  from BRepMesh,
    AsciiString      from TCollection,
    MapOfAsciiString from TColStd,
    Shape            from TopoDS,
    MapOfFunctions   from Plugin

--raises

is
    Create
        returns DiscretFactory from BRepMesh
        is protected;
    ---C++: alias "Standard_EXPORT virtual ~BRepMesh_DiscretFactory();"

    Get (myclass)
        returns DiscretFactory from BRepMesh;
    ---C++: return &
    ---Purpose:
    -- Returns the global factory instance.

    Names (me)
        returns MapOfAsciiString from TColStd;
    ---C++: return const &
    ---Purpose:
    -- Returns the list of registered meshing algorithms.

    SetDefaultName (     me : out;
                    theName : AsciiString from TCollection)
        returns Boolean from Standard;
    ---Purpose:
    -- Setup meshing algorithm by name.
    -- Returns true if requested tool is available.
    -- On fail Factory will continue to use previous algo.

    DefaultName (me)
        returns AsciiString from TCollection;
    ---C++: return const &
    ---Purpose:
    -- Returns name for current meshing algorithm.

    SetFunctionName (         me : out;
                     theFuncName : AsciiString from TCollection)
        returns Boolean from Standard;
    ---Purpose:
    -- Advanced function. Changes function name to retrieve from plugin.
    -- Returns true if requested tool is available.
    -- On fail Factory will continue to use previous algo.

    SetDefault (         me : out;
                    theName : AsciiString from TCollection;
                theFuncName : AsciiString from TCollection = "DISCRETALGO")
        returns Boolean from Standard;
    ---Purpose:
    -- Setup meshing algorithm that should be created by this Factory.
    -- Returns true if requested tool is available.
    -- On fail Factory will continue to use previous algo.
    -- Call ::ErrorStatus() method to retrieve fault reason.

    FunctionName (me)
        returns AsciiString from TCollection;
    ---C++: return const &
    ---Purpose:
    -- Returns function name that should be exported by plugin.

    Discret (me            : out;
             theShape      : Shape from TopoDS;
             theDeflection : Real  from Standard;
             theAngle      : Real  from Standard)
        returns DiscretRoot from BRepMesh;
    ---Purpose:
    -- Returns triangulation algorithm instance.

    ErrorStatus (me)
        returns FactoryError from BRepMesh;
    ---Purpose:
    -- Returns error status for last meshing algorithm switch.

    Clear (me : out)
        is protected;

fields
    myPluginEntry    : PluginEntryType from BRepMesh is protected;
    myErrorStatus    : FactoryError from BRepMesh is protected;
    myNames          : MapOfAsciiString from TColStd is protected;
    myDefaultName    : AsciiString from TCollection is protected;
    myFunctionName   : AsciiString from TCollection is protected;
    myFactoryMethods : MapOfFunctions from Plugin is protected;

end DiscretFactory;
