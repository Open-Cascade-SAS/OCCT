-- Created on: 1995-09-21
-- Created by: Philippe GIRODENGO
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MeshTriangle from StlMesh inherits TShared from MMgt

	---Purpose: A  mesh triangle is defined with
	--          three geometric vertices and an orientation
	--          

raises 

    NegativeValue from Standard

is

    Create  returns mutable MeshTriangle;
    	---Purpose: empty constructor


    Create (V1, V2, V3 : Integer; Xn, Yn, Zn : Real)  returns mutable MeshTriangle
        ---Purpose: create a triangle defined with the indexes of its three vertices 
        --          and its orientation
    raises NegativeValue;
    	---Purpose: Raised if V1, V2 or V3 is lower than zero


    GetVertexAndOrientation (me; V1, V2, V3 : out Integer; Xn, Yn, Zn : out Real);
        ---Purpose: get indexes of the three vertices (V1,V2,V3) and the orientation

    SetVertexAndOrientation (me : mutable; V1, V2, V3 : in Integer; Xn, Yn, Zn : in Real)
        ---Purpose: set indexes of the three vertices (V1,V2,V3) and the orientation
    raises NegativeValue;
    	---Purpose: Raised if V1, V2 or V3 is lower than zero


    GetVertex  (me; V1, V2, V3 : out Integer);
        ---Purpose: get indexes of the three vertices (V1,V2,V3)

    SetVertex  (me : mutable; V1, V2, V3 : in Integer)
        ---Purpose: set indexes of the three vertices (V1,V2,V3)
    raises NegativeValue;
    	---Purpose: Raised if V1, V2 or V3 is lower than zero


fields 

    MyV1     : Integer;
    MyV2     : Integer;
    MyV3     : Integer;
    MyXn     : Real;
    MyYn     : Real;
    MyZn     : Real;

end MeshTriangle;


