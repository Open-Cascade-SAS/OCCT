-- Created on: 1993-03-10
-- Created by: JCV
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class TrimmedCurve from Geom inherits BoundedCurve from Geom


        ---Purpose : Describes a portion of a curve (termed the "basis
    	-- curve") limited by two parameter values inside the
    	-- parametric domain of the basis curve.
    	-- The trimmed curve is defined by:
    	-- - the basis curve, and
    	-- - the two parameter values which limit it.
    	-- The trimmed curve can either have the same
    	-- orientation as the basis curve or the opposite orientation.

uses Ax1      from gp,
     Ax2      from gp,
     Pnt      from gp, 
     Trsf     from gp,
     Vec      from gp,
     Curve    from Geom,
     Geometry from Geom,
     Shape    from GeomAbs


raises ConstructionError   from Standard,
       RangeError          from Standard,
       NoSuchObject        from Standard,
       UndefinedDerivative from Geom,
       UndefinedValue      from Geom


is


  Create (C : Curve; U1, U2 : Real; Sense : Boolean = Standard_True)
     returns mutable TrimmedCurve
        ---Purpose : Constructs a trimmed curve from the basis curve C
    	-- which is limited between parameter values U1 and U2.
    	-- Note: - U1 can be greater or less than U2; in both cases,
    	--   the returned curve is oriented from U1 to U2.
    	-- - If the basis curve C is periodic, there is an
    	--   ambiguity because two parts are available. In this
    	--   case, the trimmed curve has the same orientation
    	--   as the basis curve if Sense is true (default value)
    	--   or the opposite orientation if Sense is false.
    	-- - If the curve is closed but not periodic, it is not
    	--   possible to keep the part of the curve which
    	--   includes the junction point (except if the junction
    	--   point is at the beginning or at the end of the
    	--   trimmed curve). If you tried to do this, you could
    	--   alter the fundamental characteristics of the basis
    	--   curve, which are used, for example, to compute
    	--   the derivatives of the trimmed curve. The rules
    	--   for a closed curve are therefore the same as
    	--   those for an open curve.
    	-- Warning: The trimmed curve is built from a copy of curve C.
    	--   Therefore, when C is modified, the trimmed curve
    	--   is not modified.
    	-- - If the basis curve is periodic, the bounds of the
    	--   trimmed curve may be different from U1 and U2
    	--   if the parametric origin of the basis curve is within
    	--   the arc of the trimmed curve. In this case, the
    	--   modified parameter will be equal to U1 or U2
    	--   plus or minus the period.
    	--   Exceptions
    	-- Standard_ConstructionError if:
    	-- - C is not periodic and U1 or U2 is outside the
    	--   bounds of C, or
    	-- - U1 is equal to U2.
     raises ConstructionError;
    



  Reverse (me : mutable);
    	---Purpose : Changes the orientation of this trimmed curve.
    	-- As a result:
    	-- - the basis curve is reversed,
    	-- - the start point of the initial curve becomes the
    	--   end point of the reversed curve,
    	-- - the end point of the initial curve becomes the
    	--   start point of the reversed curve,
    	-- - the first and last parameters are recomputed.
    	--   If the trimmed curve was defined by:
    	-- - a basis curve whose parameter range is [ 0., 1. ],
    	-- - the two trim values U1 (first parameter) and U2 (last parameter),
    	--   the reversed trimmed curve is defined by:
    	-- - the reversed basis curve, whose parameter range is still [ 0., 1. ],
    	-- - the two trim values 1. - U2 (first parameter) and 1. - U1 (last parameter).
     


  ReversedParameter(me; U : Real) returns Real;
	---Purpose: Computes the parameter on the reversed curve for
    	-- the point of parameter U on this trimmed curve.


  SetTrim (me : mutable; U1, U2 : Real; Sense : Boolean = Standard_True)
        ---Purpose :  Changes this trimmed curve, by redefining the
    	-- parameter values U1 and U2 which limit its basis curve.
    	-- Note: If the basis curve is periodic, the trimmed curve
    	-- has the same orientation as the basis curve if Sense
    	-- is true (default value) or the opposite orientation if Sense is false.
    	-- Warning
    	-- If the basis curve is periodic, the bounds of the
    	-- trimmed curve may be different from U1 and U2 if the
    	-- parametric origin of the basis curve is within the arc of
    	-- the trimmed curve. In this case, the modified
    	-- parameter will be equal to U1 or U2 plus or minus the period.
    	-- Exceptions
    	-- Standard_ConstructionError if:
    	-- - the basis curve is not periodic, and either U1 or U2
    	--   are outside the bounds of the basis curve, or
    	-- - U1 is equal to U2.
     raises ConstructionError;
      


  BasisCurve (me)    returns Curve;
        ---Purpose : Returns the basis curve. 
        --   Warning
    	-- This function does not return a constant reference.
    	-- Consequently, any modification of the returned value
    	-- directly modifies the trimmed curve.


  Continuity (me)  returns Shape from GeomAbs;
        ---Purpose :
        --  Returns the continuity of the curve :
        -- C0 : only geometric continuity,
        -- C1 : continuity of the first derivative all along the Curve,
        -- C2 : continuity of the second derivative all along the Curve,
        -- C3 : continuity of the third derivative all along the Curve,
        -- CN : the order of continuity is infinite.


  IsCN (me; N : Integer)   returns Boolean
        ---Purpose : Returns true if the degree of continuity of the basis
    	-- curve of this trimmed curve is at least N. A trimmed
    	-- curve is at least "C0" continuous.
        --  Warnings :
        --  The continuity of the trimmed curve can be greater than
        --  the continuity of the basis curve because you consider
        --  only a part of the basis curve.
     raises RangeError;
        ---Purpose : Raised if N < 0.


  EndPoint (me)   returns Pnt;
	---Purpose :
	--  Returns the end point of <me>. This point is the
	--  evaluation of the curve for the "LastParameter".


  FirstParameter (me)   returns Real;
        ---Purpose :
	--  Returns the value of the first parameter of <me>. 
        --  The first parameter is the parameter of the "StartPoint"
        --  of the trimmed curve.


  IsClosed (me)  returns Boolean;
        ---Purpose :
        --  Returns True if the distance between the StartPoint and
        --  the EndPoint is lower or equal to Resolution from package gp.


  IsPeriodic (me)   returns Boolean;
        ---Purpose : Returns true if the basis curve of this trimmed curve is periodic.


  Period (me) returns Real from Standard 
	---Purpose: Returns the period of the basis curve of this trimmed curve.
    	-- Exceptions
    	-- Standard_NoSuchObject if the basis curve is not periodic.
  raises
    	NoSuchObject from Standard
  is redefined;


  LastParameter (me)  returns Real;
	---Purpose :
	--  Returns the value of the last parameter of <me>.
        --  The last parameter is the parameter of the "EndPoint" of the
        --  trimmed curve.


  StartPoint (me)  returns Pnt;
	---Purpose :
	--  Returns the start point of <me>.
	--  This point is the evaluation of the curve from the 
	--  "FirstParameter".






        ---Purpose  : value and derivatives
        --- Warnings :
        --  The returned derivatives have the same orientation as the
        --  derivatives of the basis curve even if the trimmed curve 
        --  has not the same orientation as the basis curve.


  D0(me; U : Real; P : out Pnt);
	---Purpose: Returns in P the point of parameter U.
	--          
        --  If the basis curve is an OffsetCurve sometimes it is not 
        --  possible to do the evaluation of the curve at the parameter
        --  U (see class OffsetCurve).


  D1 (me; U : Real; P : out Pnt; V1 : out Vec)
     raises UndefinedDerivative;
        ---Purpose : Raised if the continuity of the curve is not C1.


  D2 (me; U : Real; P : out Pnt; V1, V2 : out Vec)
     raises UndefinedDerivative;
        ---Purpose : Raised if the continuity of the curve is not C2.


  D3 (me; U : Real; P : out Pnt; V1, V2, V3 : out Vec)
     raises UndefinedDerivative;
        ---Purpose : Raised if the continuity of the curve is not C3.
        

  DN (me; U : Real; N : Integer)  returns Vec
        ---Purpose  : N is the order of derivation.
     raises  UndefinedDerivative,
        ---Purpose : Raised if the continuity of the curve is not CN.
             RangeError;
        ---Purpose : Raised if N < 1.            





        ---Purpose : geometric transformations

  Transform (me : mutable; T : Trsf);
        --- Purpose: Applies the transformation T to this trimmed curve.
    	-- Warning The basis curve is also modified.

  TransformedParameter(me; U : Real; T : Trsf from gp) returns Real
	---Purpose: Returns the  parameter on the  transformed  curve for
	--          the transform of the point of parameter U on <me>.
	--          
	--          me->Transformed(T)->Value(me->TransformedParameter(U,T))
	--          
	--          is the same point as
	--          
	--          me->Value(U).Transformed(T)
	--          
	--          This methods calls the basis curve method.
     is redefined;  

  ParametricTransformation(me; T : Trsf from gp) returns Real
	---Purpose: Returns a  coefficient to compute the parameter on
	--          the transformed  curve  for  the transform  of the
	--          point on <me>.
	--          
	--          Transformed(T)->Value(U * ParametricTransformation(T))
	--          
	--          is the same point as
	--          
	--          Value(U).Transformed(T)
	--          
	--          This methods calls the basis curve method.
     is redefined;  

  Copy (me)  returns mutable like me;
    	---Purpose: Creates a new object which is a copy of this trimmed curve.
    
fields

    basisCurve : Curve;
    uTrim1     : Real;
    uTrim2     : Real;

end;





