-- Created on: 2000-05-10
-- Created by: Andrey BETENEV
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1

class EffectivityAssignment from StepBasic
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity EffectivityAssignment

uses
    Effectivity from StepBasic

is
    Create returns EffectivityAssignment from StepBasic;
	---Purpose: Empty constructor

    Init (me: mutable; aAssignedEffectivity: Effectivity from StepBasic);
	---Purpose: Initialize all fields (own and inherited)

    AssignedEffectivity (me) returns Effectivity from StepBasic;
	---Purpose: Returns field AssignedEffectivity
    SetAssignedEffectivity (me: mutable; AssignedEffectivity: Effectivity from StepBasic);
	---Purpose: Set field AssignedEffectivity

fields
    theAssignedEffectivity: Effectivity from StepBasic;

end EffectivityAssignment;
