-- Created on: 1997-04-17
-- Created by: Christophe MARION
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Hider from HLRBRep

uses
    Integer         from Standard,
    Boolean         from Standard,
    Real            from Standard,
    ShortReal       from Standard,
    ListOfInteger   from TColStd,
    MapOfShapeTool  from BRepTopAdaptor,
    Data            from HLRBRep

is
    Create(DS : Data from HLRBRep)
    returns Hider from HLRBRep;
	---Purpose: Creates a Hider processing  the set  of  Edges and
	--          hiding faces described by <DS>.  Stores the hidden
	--          parts in <DS>.

    OwnHiding(me : in out; FI : Integer from Standard)
	---Purpose: own hiding the side face number <FI>.
    is static;

    Hide(me : in out; FI :        Integer from Standard;
                      MST: in out MapOfShapeTool from BRepTopAdaptor)
	---Purpose: Removes from the edges,   the parts hidden by  the
	--          hiding face number <FI>.
    is static;

fields
    myDS : Data from HLRBRep;

end Hider;
