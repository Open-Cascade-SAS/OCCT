-- Created on: 1992-11-17
-- Created by: Christian CAILLET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class SelectModelEntities  from IFSelect  inherits SelectBase

    ---Purpose : A SelectModelEntities gets all the Entities of an
    --           InterfaceModel.

uses AsciiString from TCollection, EntityIterator, Graph

is

    Create  returns mutable SelectModelEntities;
    ---Purpose : Creates a SelectModelRoot

    RootResult (me; G : Graph) returns EntityIterator;
    ---Purpose : Returns the list of selected entities : the Entities of the
    --           Model (note that this result assures naturally uniqueness)

    CompleteResult (me; G : Graph) returns EntityIterator  is redefined;
    ---Purpose : The complete list of Entities (including shared ones) ...
    --           is exactly identical to RootResults in this case

    Label (me) returns AsciiString from TCollection;
    ---Purpose : Returns a text defining the criterium : "Model Entities"

end SelectModelEntities;
