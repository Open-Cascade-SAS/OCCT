-- Created on: 1997-04-02
-- Created by: Administrateur Atelier XSTEP
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class EDescr  from StepData    inherits TShared

    ---Purpose : This class is intended to describe the authorized form for an
    --           entity, either Simple or Plex

uses CString,
     Described from StepData

is

    Matches    (me; steptype : CString) returns Boolean  is deferred;
    ---Purpose : Tells if a ESDescr matches a step type : exact or super type

    IsComplex  (me) returns Boolean  is deferred;
    ---Purpose : Tells if a EDescr is complex (ECDescr) or simple (ESDescr)

    NewEntity  (me) returns mutable Described  is deferred;
    ---Purpose : Creates a described entity (i.e. a simple one)

end EDescr;
