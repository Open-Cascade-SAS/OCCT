-- File:	QASamtech.cdl
-- Created:	Mon Mar 18 18:37:01 2002
-- Author:	QA Admin
--		<qa@umnox.nnov.matra-dtv.fr>
---Copyright:	 Matra Datavision 2002

package QASamtech
     uses Draw
is
    Commands(DI : in out Interpretor from Draw);
end;
    
