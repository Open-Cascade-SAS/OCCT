-- File:	MeshAlgo_PntComparator.cdl
-- Created:	Fri Jun 18 13:46:14 1993
-- Author:	Didier PIFFAULT
--		<dpf@zerox>
---Copyright:	 Matra Datavision 1993


generic class PntComparator from MeshAlgo (Point as any; Direction as any)

	---Purpose: Sort two point in a given direction.


uses  Boolean from Standard


is      Create (theDir : Direction; TheTol: Real from Standard) 
    	    returns PntComparator;


    	IsLower (me; Left, Right: Point)
	---Purpose: returns True if <Left> is lower than <Right>
    	    returns Boolean from Standard;
    
    	IsGreater (me; Left, Right: Point)
	---Purpose: returns True if <Left> is greater than <Right>
    	    returns Boolean from Standard;

    	IsEqual(me; Left, Right: Point)
	---Purpose: returns True when <Right> and <Left> are equal.
	    returns Boolean from Standard;


fields  DirectionOfSort : Direction;
    	Tolerance       : Real from Standard;

end PntComparator;
