-- Created on: 2002-12-12
-- Created by: data exchange team
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class ElementMaterial from StepElement
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity ElementMaterial

uses
    HAsciiString from TCollection,
    HArray1OfMaterialPropertyRepresentation from StepRepr

is
    Create returns ElementMaterial from StepElement;
	---Purpose: Empty constructor

    Init (me: mutable; aMaterialId: HAsciiString from TCollection;
                       aDescription: HAsciiString from TCollection;
                       aProperties: HArray1OfMaterialPropertyRepresentation from StepRepr);
	---Purpose: Initialize all fields (own and inherited)

    MaterialId (me) returns HAsciiString from TCollection;
	---Purpose: Returns field MaterialId
    SetMaterialId (me: mutable; MaterialId: HAsciiString from TCollection);
	---Purpose: Set field MaterialId

    Description (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Description
    SetDescription (me: mutable; Description: HAsciiString from TCollection);
	---Purpose: Set field Description

    Properties (me) returns HArray1OfMaterialPropertyRepresentation from StepRepr;
	---Purpose: Returns field Properties
    SetProperties (me: mutable; Properties: HArray1OfMaterialPropertyRepresentation from StepRepr);
	---Purpose: Set field Properties

fields
    theMaterialId: HAsciiString from TCollection;
    theDescription: HAsciiString from TCollection;
    theProperties: HArray1OfMaterialPropertyRepresentation from StepRepr;

end ElementMaterial;
