-- Created on: 1992-12-24
-- Created by: Denis PASCAL
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

generic class TopologicalSortIterator from GraphTools
             (Graph      as any;
    	      Vertex     as any; 
              GIterator  as any;
	      TSIterator as any)
	      
--generic class TopologicalSorIterator from GraphTools
--    	         (Graph     as any;
--    	          Vertex    as any;
--    	          GIterator as GraphIterator (Graph,Vertex))
--	          TSIterator as TopologicalSortFromIterator

	---Purpose: This  generic class defines  an  iterator to visit
	--          each vertex of the  underlying graph,  in  such an
	--          order that noone vertex is reach before any vertex
	--          that point to it. In general the order produced by
	--          topological sort  is  not unique. Usefull  for DAG
	--          Topological Sort.

raises NoSuchObject from Standard,
       NoMoreObject from Standard

    
is

    Create    	
    	---Purpose: Create an empty algorithm. 
    returns TopologicalSortIterator from GraphTools;
    
    Create (G : Graph)
	---Purpose: Create the   algorithm setting each vertex  of <G>
	--          reached by  GIterator tool, as initial conditions.
	--          Use Perform   method before visting  the result of
	--          the algorithm.
    returns TopologicalSortIterator from GraphTools;
    
    FromGraph (me : in out; G : Graph); 
	---Purpose: Add each vertex of <G>  reached by GIterator  tool
	--          as   initial  conditions.   Use  Perform  method
	--          before   visiting the  result  of   the algorithm.
        ---Level: Public
    
    FromVertex (me : in out; V : Vertex);
	---Purpose: Add  <V>  as  initial  condition.  This method  is
	--          cumulative.  Use Perform method before visting the
	--          result of the algorithm.  
	---Level: Public

    Reset (me : in out);
	---Purpose: Reset the algorithm.   It may  be reused with  new
	--          initial conditions.  
	---Level: Public

    Perform (me : in out; G              : Graph ;
                          ignoreSelfLoop : Boolean from Standard;
                          processCycle   : Boolean from Standard);    	
    	---Purpose: Peform the  algorithm  in  <G> from initial setted
    	--          conditions according to  the two following flags.
	--          * <ignoreSelfLoop>  allows the  user to ignore (or
	--          not) any vertex wich contains a self loop.
	--          * <processCycle> allows the user to visit (or not>
	--          vertex which is in a cycle.
       ---Level: Public
    
    More (me) 
    returns Boolean from Standard;
       ---Level: Public
    
    Next (me : in out) 
    raises NoMoreObject from Standard;
       ---Level: Public
    
    Value (me) returns any Vertex
       ---Level: Public
    	---C++: return const &
    raises NoSuchObject from Standard;

    IsInCycle (me) returns Boolean from Standard
	---Purpose: Returns TRUE if the current vertex is in a cycle.
       ---Level: Public
    raises NoSuchObject from Standard;
    
fields

   myIterator : TSIterator; 

end TopologicalSortIterator;




