-- Created by: Peter KURNEV
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class AlgoTools2D from BOPTools 

      ---Purpose: 
      ---  The class contains handy static functions 
      ---  dealing with the topology  
      ---  This is the copy of the BOPTools_AlgoTools2D.cdl
uses 
    Vec  from gp, 
    Dir  from gp, 
    Vertex from TopoDS,
    Edge   from TopoDS, 
    Face   from TopoDS, 
    Surface from BRepAdaptor, 
    Curve from Geom2d,
    Curve from Geom, 
    ProjectedCurve from ProjLib, 
    Context from IntTools, 
    ListOfShape from BOPCol 
    
is   

    BuildPCurveForEdgeOnFace  (myclass; 
              aE:  Edge from TopoDS; 
              aF:  Face from TopoDS); 
          ---Purpose: 
          --- Compute P-Curve for the edge <aE> on the face <aF> 
          --- Raises exception Standard_ConstructionError if projection algorithm fails

    EdgeTangent     (myclass;  
              anE  : Edge from TopoDS; 
              aT   : Real from Standard; 
              Tau  : out Vec  from gp) 
          returns  Boolean from Standard; 
          ---Purpose: 
          --- Compute tangent for the edge  <aE> [in 3D]  at parameter <aT> 
          ---
 
    PointOnSurface  (myclass; 
              aE:  Edge from TopoDS; 
              aF:  Face from TopoDS;  
              aT:  Real from Standard; 
              U : out Real from Standard; 
              V : out Real from Standard); 
          ---Purpose: 
          --- Compute surface parameters <U,V> of the face <aF> 
          --- for  the point from the edge <aE> at parameter <aT>. 
          --- If <aE> has't pcurve on surface, algorithm tries to get it by
          --- projection and can  
          --- raise exception Standard_ConstructionError if projection algorithm fails

    CurveOnSurface  (myclass; 
              aE:  Edge from TopoDS; 
              aF:  Face from TopoDS; 
              aC    : out Curve from Geom2d; 
              aToler: out Real from Standard); 
          ---Purpose:  
          --- Get P-Curve <aC>  for the edge <aE> on surface <aF> . 
          --- If the P-Curve does not exist, build  it using Make2D(). 
          --- [aToler] - reached tolerance 
          --- Raises exception Standard_ConstructionError if algorithm Make2D() fails

    CurveOnSurface  (myclass; 
              aE:  Edge from TopoDS; 
              aF:  Face from TopoDS; 
              aC    : out Curve from Geom2d; 
              aFirst: out Real from Standard; 
              aLast : out Real from Standard; 
              aToler: out Real from Standard); 
                      
          ---Purpose: 
          --- Get P-Curve <aC>  for the edge <aE> on surface <aF> . 
          --- If the P-Curve does not exist, build  it using Make2D(). 
          --- [aFirst, aLast] - range of the P-Curve    
          --- [aToler] - reached tolerance 
          --- Raises exception Standard_ConstructionError if algorithm Make2D() fails

    HasCurveOnSurface  (myclass;  
              aE:  Edge from TopoDS; 
              aF:  Face from TopoDS; 
              aC    : out Curve from Geom2d;
              aFirst: out Real from Standard; 
              aLast : out Real from Standard; 
              aToler: out Real from Standard) 
          returns  Boolean from Standard; 
          ---Purpose:  
          --- Returns TRUE if the edge <aE>  has  P-Curve <aC>           
          --- on surface <aF> .   
          --- [aFirst, aLast] - range of the P-Curve    
          --- [aToler] - reached tolerance 
          --- If the P-Curve does not exist, aC.IsNull()=TRUE. 
          ---
    HasCurveOnSurface  (myclass;  
              aE:  Edge from TopoDS; 
              aF:  Face from TopoDS) 
          returns  Boolean from Standard;  
          ---Purpose:  
          --- Returns TRUE if the edge <aE>  has  P-Curve <aC>           
          --- on surface <aF> .   
          --- If the P-Curve does not exist, aC.IsNull()=TRUE. 
          ---
 
    AdjustPCurveOnFace  (myclass;    
              aF    :  Face from TopoDS; 
              C3D   :  Curve from Geom; 
              aC2D  :  Curve from Geom2d; 
              aC2DA : out Curve from Geom2d);                  
          ---Purpose:   
          --- Adjust P-Curve <aC2D> (3D-curve <C3D>) on surface <aF> .  
          ---
    AdjustPCurveOnFace  (myclass;    
              aF    :  Face from TopoDS; 
              aT1   :  Real from Standard;   
              aT2   :  Real from Standard;   
              aC2D  :  Curve from Geom2d; 
              aC2DA : out Curve from Geom2d); 
          ---Purpose:   
          --- Adjust P-Curve <aC2D> (3D-curve <C3D>) on surface <aF> .  
          --- [aT1,  aT2] - range to adjust 
          ---
    AdjustPCurveOnFace  (myclass;    
              aF    :  Surface from BRepAdaptor; 
              aT1   :  Real from Standard;   
              aT2   :  Real from Standard;   
              aC2D  :  Curve from Geom2d; 
              aC2DA : out Curve from Geom2d); 
          ---Purpose:   
          --- Adjust P-Curve <aC2D> (3D-curve <C3D>) on surface <aF> .  
          --- [aT1,  aT2] - range to adjust 
          --- 
    IntermediatePoint (myclass; 
              aFirst: Real from Standard; 
              aLast : Real from Standard) 
          returns  Real from Standard; 
          ---Purpose:   
          --- Compute intermediate  value in  between [aFirst, aLast] . 
          ---
    IntermediatePoint        (myclass;  
              anE  : Edge from TopoDS) 
          returns  Real from Standard;
          ---Purpose:   
          --- Compute intermediate value of parameter for the edge <anE>. 
          ---
    BuildPCurveForEdgeOnPlane(myclass; 
              theE : Edge from TopoDS; 
              theF : Face from TopoDS); 
	      
    BuildPCurveForEdgesOnPlane(myclass; 
              theLE : ListOfShape from BOPCol; 
              theF : Face from TopoDS);
 
    Make2D  (myclass;  
              aE:  Edge from TopoDS; 
              aF:  Face from TopoDS; 
              aC    : out Curve from Geom2d;
              aFirst: out Real from Standard; 
              aLast : out Real from Standard; 
              aToler: out Real from Standard);            
          ---Purpose:   
          --- Make P-Curve <aC> for the edge <aE> on surface <aF> . 
          --- [aFirst, aLast] - range of the P-Curve    
          --- [aToler] - reached tolerance 
          --- Raises exception Standard_ConstructionError if algorithm fails
          
    MakePCurveOnFace  (myclass;    
              aF:  Face from TopoDS; 
              C3D   :     Curve from Geom; 
              aC    : out Curve from Geom2d; 
              aToler: out Real from Standard) ;   
          ---Purpose:   
          --- Make P-Curve <aC> for the 3D-curve <C3D> on surface <aF> . 
          --- [aToler] - reached tolerance 
          --- Raises exception Standard_ConstructionError if projection algorithm fails

    MakePCurveOnFace  (myclass;    
              aF:  Face from TopoDS; 
              C3D   :     Curve from Geom;  
              aT1   :  Real from Standard;   
              aT2   :  Real from Standard;      
              aC    : out Curve from Geom2d; 
              aToler: out Real from Standard) ;                  
          ---Purpose:   
          --- Make P-Curve <aC> for the 3D-curve <C3D> on surface <aF> .  
          --- [aT1,  aT2] - range to build    
          --- [aToler] - reached tolerance 
          --- Raises exception Standard_ConstructionError if projection algorithm fails

    MakePCurveOfType  (myclass;    
              PC  : ProjectedCurve from ProjLib; 
              aC  : out Curve from Geom2d);         
          ---Purpose:   
          --- Make empty  P-Curve <aC> of relevant to <PC> type  
          ---
    AttachExistingPCurve (myclass;    
              aEold :  Edge from TopoDS; 
              aEnew :  Edge from TopoDS; 
              aF    :  Face from TopoDS; 
              aCtx  :  Context from IntTools) 
        returns Integer from Standard;   
          ---Purpose:   
          --- Attach P-Curve from the edge <aEold> on surface <aF>   
          --- to the edge <aEnew>  
          --- Returns 0 in case of success  
     
end AlgoTools2D;
