-- Created on: 2000-04-18
-- Created by: Andrey BETENEV
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0

class DimensionalSize from StepShape
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity DimensionalSize

uses
    ShapeAspect from StepRepr,
    HAsciiString from TCollection

is
    Create returns DimensionalSize from StepShape;
	---Purpose: Empty constructor

    Init (me: mutable; aAppliesTo: ShapeAspect from StepRepr;
                       aName: HAsciiString from TCollection);
	---Purpose: Initialize all fields (own and inherited)

    AppliesTo (me) returns ShapeAspect from StepRepr;
	---Purpose: Returns field AppliesTo
    SetAppliesTo (me: mutable; AppliesTo: ShapeAspect from StepRepr);
	---Purpose: Set field AppliesTo

    Name (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Name
    SetName (me: mutable; Name: HAsciiString from TCollection);
	---Purpose: Set field Name

fields
    theAppliesTo: ShapeAspect from StepRepr;
    theName: HAsciiString from TCollection;

end DimensionalSize;
