-- Created on: 1994-03-23
-- Created by: Bruno DUMORTIER
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


package Geom2dAPI

	---Purpose: The  Geom2dAPI  package  provides  an  Application
	--          Programming Interface for the Geometry.
	--          
	--          The API is a set of classes aiming to provide :
	--          
	--          * High level and simple calls  for the most common
	--          operations. 
	--          
	--          *    Keeping   an   access  on    the    low-level
	--          implementation of high-level calls.
	--          
	-- 	    
	-- 	    The API  provides classes to  call the algorithmes
	-- 	    of the Geometry
	-- 	    
	-- 	    * The  constructors  of the classes  provides  the
	-- 	    different constructions methods.
	-- 	    
	-- 	    * The  class keeps as fields the   different tools
	-- 	    used by the algorithmes
	-- 	    
	-- 	    *   The class  provides  a  casting  method to get
	-- 	    automatically the  result  with  a   function-like
	-- 	    call. 
	-- 	    
	-- 	    For example to evaluate the distance <D> between a
	-- 	    point <P> and a curve <C>, one can writes :
	-- 	    
	-- 	        D = Geom2dAPI_ProjectPointOnCurve(P,C);
	-- 	    
	-- 	    or
	-- 	    
	-- 	        Geom2dAPI_ProjectPointOnCurve PonC(P,C);
	-- 	        D = PonC.LowerDistance();
	-- 	    


uses

    Geom2d,
    gp,
    TColgp,
    Extrema,
    Geom2dAdaptor,
    Geom2dInt,
    GeomAbs,
    TColStd,
    Quantity, 
    Approx,
    StdFail
    

is

    ------------------------------------------------------------------
    -- This classes  provides algo  to  evaluate  the distance between
    -- points and curves, curves and curves. 
    ------------------------------------------------------------------

    class ProjectPointOnCurve;

    class ExtremaCurveCurve;
    


    ------------------------------------------------------------------
    -- This classes provides algo to evaluate a curve  passing through
    -- an array of points.
    ------------------------------------------------------------------

    --- Approximation:
    --  
    class PointsToBSpline;
    
    
    --- Interpolation:
    --
    class Interpolate;
    
    
    ------------------------------------------------------------------
    -- This classes provides algo to evaluate an intersection between 
    -- two 2d-Curves.
    ------------------------------------------------------------------

    class InterCurveCurve;


end Geom2dAPI;
