-- File:	IGESGraph_ToolDrawingSize.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolDrawingSize  from IGESGraph

    ---Purpose : Tool to work on a DrawingSize. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses DrawingSize from IGESGraph,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolDrawingSize;
    ---Purpose : Returns a ToolDrawingSize, ready to work


    ReadOwnParams (me; ent : mutable DrawingSize;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : DrawingSize;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : DrawingSize;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a DrawingSize <ent>, from
    --           its specific (own) parameters

    OwnCorrect (me; ent : mutable DrawingSize) returns Boolean  is static;
    ---Purpose : Sets automatic unambiguous Correction on a DrawingSize
    --           (NbPropertyValues forced to 2)

    DirChecker (me; ent : DrawingSize) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : DrawingSize;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : DrawingSize; entto : mutable DrawingSize;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : DrawingSize;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolDrawingSize;
