-- Created on: 1993-08-11
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class PointRepresentation from PBRep inherits Persistent

	---Purpose: Root class for points representations.

uses
    Location from PTopLoc

is
    Initialize(P : Real;
    	       L : Location from PTopLoc);
    	---Level: Internal 
	       
    Location(me) returns Location from PTopLoc
    is static;
    	---Level: Internal 
		
    Parameter(me) returns Real
    is static;
    	---Level: Internal 
		
    Parameter(me : mutable; P : Real)
    is static;
    	---Level: Internal 
		
    Next(me) returns PointRepresentation from PBRep
    is static;
    	---Level: Internal 
		
    Next(me : mutable; N :  PointRepresentation from PBRep)
    is static;
    	---Level: Internal 

    ------------------------------------------------------
    -- What kind of representation : used to speed Mapping
    ------------------------------------------------------

    IsPointOnCurve(me)          returns Boolean
	---Purpose: A point on a 3d curve.
    is virtual;
	
    IsPointOnCurveOnSurface(me) returns Boolean
	---Purpose: A point on a 2d curve on a surface.
    is virtual;

    IsPointOnSurface(me)        returns Boolean
	---Purpose: A point on a surface.
    is virtual;
    
fields
    
    myLocation  : Location from PTopLoc;
    myParameter : Real;
    myNext      : PointRepresentation from PBRep;

end PointRepresentation;
