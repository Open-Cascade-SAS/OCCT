-- Created on: 1996-03-08
-- Created by: Robert COUBLANC
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class FaceFilter from StdSelect inherits Filter from SelectMgr

	---Purpose: A framework to define a filter to select a specific type of face.
    	-- The types available include:
    	-- -   any face
    	-- -   a planar face
    	-- -   a cylindrical face
    	-- -   a spherical face
    	-- -   a toroidal face
    	-- -   a revol face.

uses
    TypeOfFace from StdSelect,
    Shape from TopoDS,
    EntityOwner from SelectMgr,
    ShapeEnum from TopAbs
is

    Create (aTypeOfFace: TypeOfFace from StdSelect)
    returns mutable FaceFilter from StdSelect;
    	---Purpose: Constructs a face filter object defined by the type of face aTypeOfFace.    
    SetType(me:mutable;aNewType : TypeOfFace from StdSelect);  
    	--- Purpose: Sets the type of face aNewType. aNewType is to be highlighted in selection.   
    Type(me) returns TypeOfFace from StdSelect;
    	--- Purpose: Returns the type of face to be highlighted in selection.   
    IsOk (me;anobj : EntityOwner from SelectMgr) 
    returns Boolean from Standard is redefined virtual;
  
    ActsOn(me; aStandardMode : ShapeEnum from TopAbs)
    returns Boolean from Standard is redefined virtual;
   
fields

    mytype : TypeOfFace from StdSelect;

end FaceFilter;
