-- Created on: 1993-01-09
-- Created by: CKY / Contract Toubro-Larsen ( SIVA )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PlaneSurface from IGESSolid  inherits IGESEntity

        ---Purpose: defines PlaneSurface, Type <190> Form Number <0,1>
        --          in package IGESSolid
        --          A plane surface entity is defined by a point on the
        --          surface and a normal to it.

uses

        Point           from IGESGeom,
        Direction       from IGESGeom

is

        Create returns mutable PlaneSurface;

        -- Specific Methods pertaining to the class

        Init (me        : mutable;
              aLocation : Point;
              aNormal   : Direction;
              refdir    : Direction);
        ---Purpose : This method is used to set the fields of the class
        --           PlaneSurface
        --       - aLocation : the point on the surface
        --       - aNormal   : the surface normal direction
        --       - refdir    : the reference direction (default NULL) for
        --                    unparameterised curves

        LocationPoint(me) returns Point;
        ---Purpose : returns the point on the surface

        Normal(me) returns Direction;
        ---Purpose : returns the normal to the surface

        ReferenceDir(me) returns Direction;
        ---Purpose : returns the reference direction (for parameterised curve)
        -- returns NULL for unparameterised curve

        IsParametrised(me) returns Boolean;
        ---Purpose : returns True if parameterised, else False

fields

--
-- Class    : IGESSolid_PlaneSurface
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class PlaneSurface.
--
-- Reminder : A PlaneSurface instance is defined by :
--            A plane surface entity is defined by a point(Location) on the
--            surface and a normal(Normal) to it. In case of parameterised
--            surface a reference direction (RefDir) is also given.
--

        theLocationPoint : Point;
            -- the point on the surface

        theNormal        : Direction;
            -- the normal to the surface

        theRefDir        : Direction;
            -- the reference direction of the surface

end PlaneSurface;
