-- Created on: 1996-01-29
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class WireToFace from TopOpeBRepBuild

---Purpose: 
-- This class builds faces from a set of wires  SW and a face F.
-- The face must have and underlying surface, say S.
-- All of the edges of all of the wires must have a 2d representation 
-- on surface S (except if S is planar)

uses

    Wire from TopoDS,
    Face from TopoDS,
    ListOfShape from TopTools

is

    Create returns WireToFace;
     
    Init(me : in out)
    is static;
    
    AddWire(me : in out; W : Wire from TopoDS)
    is  static;
     	
    MakeFaces(me : in out; 
    	      F : Face from TopoDS;
    	      LF : in out ListOfShape from TopTools)
    is static;

fields 

    myLW : ListOfShape from TopTools;
    
end WireToFace;
