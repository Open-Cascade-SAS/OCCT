-- File:        ApprovalDateTime.cdl
-- Created:     Mon Dec  4 12:02:28 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWApprovalDateTime from RWStepBasic

	---Purpose : Read & Write Module for ApprovalDateTime

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     ApprovalDateTime from StepBasic,
     EntityIterator from Interface

is

	Create returns RWApprovalDateTime;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable ApprovalDateTime from StepBasic);

	WriteStep (me; SW : in out StepWriter; ent : ApprovalDateTime from StepBasic);

	Share(me; ent : ApprovalDateTime from StepBasic; iter : in out EntityIterator);

end RWApprovalDateTime;
