-- Created on: 1994-11-04
-- Created by: Christian CAILLET
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class ElemHasher  from MoniTool

    ---Purpose : ElemHasher defines HashCode for Element, which is : ask a
    --           Element its HashCode !  Because this is the Element itself
    --           which brings the HashCode for its Key
    --           
    --           This class complies to the template given in TCollection by
    --           MapHasher itself

uses Element

is

    HashCode (myclass; K : Element; Upper : Integer) returns Integer;
    ---Purpose : Returns a HashCode in the range <0,Upper> for a Element :
    --           asks the Element its HashCode then transforms it to be in the
    --           required range

    IsEqual (myclass; K1, K2 : Element) returns Boolean;
    ---Purpose : Returns True if two keys are the same.
    --           The test does not work on the Elements themselves but by
    --           calling their methods Equates

end ElemHasher;
