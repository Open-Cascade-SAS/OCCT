-- Created on: 1993-11-10
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class WPointInter from TopOpeBRep 

  -- as WPointTool from TopOpeLine
  -- 	 (PntOn2S from IntSurf)
  -- 	 

	---Purpose: 

uses

  PntOn2S from IntSurf,
  PPntOn2S from TopOpeBRep,
  Pnt2d from gp,
  Pnt from gp
  
is

  Create returns WPointInter from TopOpeBRep;
  
  Set(me : in out; P : PntOn2S from IntSurf) is static;

  ParametersOnS1(me; U,V : out Real from Standard) is static;
		  
  ParametersOnS2(me; U,V : out Real from Standard) is static;
		  
  Parameters(me; U1,V1,U2,V2 : out Real from Standard) is static;
	    
  ValueOnS1(me) returns Pnt2d from gp is static;
	
  ValueOnS2(me) returns Pnt2d from gp is static;
	
  Value(me) returns Pnt from gp is static;
   ---C++: return const &

  PPntOn2SDummy(me) returns PPntOn2S from TopOpeBRep;

fields

    myPP2S : PPntOn2S from TopOpeBRep;

end WPointInter;
