-- Created on: 1994-04-01
-- Created by: Modelistation
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package BRepTopAdaptor 

	---Purpose: 
	--          
	--          
	--          *** Class2d    : Low level algorithm for 2d classification
	--          
	--          *** FClass2d   : 2d classification on a Face from TopoDS
	--                           A face is first loaded and then every 
	--                           classification is computed as a rejection.                        
	--                           (call BRepClass algorithms if necessary,
	--                           ie, when the rejection is not efficient)
	--                           
	--          *** TopolTool :  Several tools used by the intersection
	--                           algorithm and topology.
	--         
	--          

	---Level: Internal

uses Adaptor3d, TopExp, TopoDS, BRepAdaptor, gp, TopAbs,  Adaptor2d  ,
     TColgp,TColStd,TCollection,TopTools, CSLib

is

    --class Class2d;

    alias SeqOfPtr is SequenceOfAddress from TColStd;

    class FClass2d; 

    class HVertex; -- inherits HVertex from Adaptor3d

    class TopolTool; -- inherits TopolTool from Adaptor3d
    


    --- the folowing classes are used to compute and store 
    --  informations on shapes. ( TopolTool , Bnd_Box ... )
    
    class Tool; 
    
    class MapOfShapeTool  instantiates DataMap from TCollection
        (Shape          from TopoDS,
         Tool           from BRepTopAdaptor,
         ShapeMapHasher from TopTools);


end BRepTopAdaptor;
