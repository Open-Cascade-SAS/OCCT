-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Hypr   from gp   inherits Storable

        --- Purpose : Describes a branch of a hyperbola in 3D space.
        -- A hyperbola is defined by its major and minor radii and
        -- positioned in space with a coordinate system (a gp_Ax2
        -- object) of which:
        -- -   the origin is the center of the hyperbola,
        -- -   the "X Direction" defines the major axis of the
        --   hyperbola, and
        -- - the "Y Direction" defines the minor axis of the hyperbola.
        -- The origin, "X Direction" and "Y Direction" of this
        -- coordinate system together define the plane of the
        -- hyperbola. This coordinate system is the "local
        -- coordinate system" of the hyperbola. In this coordinate
        -- system, the equation of the hyperbola is:
        -- X*X/(MajorRadius**2)-Y*Y/(MinorRadius**2) = 1.0
        -- The branch of the hyperbola described is the one located
        -- on the positive side of the major axis.
        -- The "main Direction" of the local coordinate system is a
        -- normal vector to the plane of the hyperbola. This vector
        -- gives an implicit orientation to the hyperbola. We refer to
        -- the "main Axis" of the local coordinate system as the
        -- "Axis" of the hyperbola.
        -- The following schema shows the plane of the hyperbola,
        -- and in it, the respective positions of the three branches of
        -- hyperbolas constructed with the functions OtherBranch,
        -- ConjugateBranch1, and ConjugateBranch2:
        --
        --                         ^YAxis                
        --                         |                   
        --                  FirstConjugateBranch     
        --                         |        
        --        Other            |                Main
        --   --------------------- C ------------------------------>XAxis
        --        Branch           |                Branch
        --                         |
        --                         |         
        --                   SecondConjugateBranch
        --                         |                  ^YAxis
        -- Warning
        -- The major radius can be less than the minor radius.
        -- See Also
        -- gce_MakeHypr which provides functions for more
        -- complex hyperbola constructions
        -- Geom_Hyperbola which provides additional functions for
        -- constructing hyperbolas and works, in particular, with the
        -- parametric equations of hyperbolas

uses Ax1  from gp,
     Ax2  from gp,
     Pln  from gp,
     Pnt  from gp,
     Trsf from gp,
     Vec  from gp

raises ConstructionError from Standard,
       DomainError       from Standard

is



  Create   returns Hypr;
        ---C++: inline
        --- Purpose : Creates of an indefinite hyperbola.


  Create (A2 : Ax2; MajorRadius, MinorRadius : Real)  returns Hypr
        ---C++: inline
	--- Purpose : Creates a hyperbola with radii MajorRadius and
        --   MinorRadius, positioned in the space by the
        --   coordinate system A2 such that:
        --   -   the origin of A2 is the center of the hyperbola,
        --   -   the "X Direction" of A2 defines the major axis of
        --    the hyperbola, that is, the major radius
        --    MajorRadius is measured along this axis, and
        --   -   the "Y Direction" of A2 defines the minor axis of
        --    the hyperbola, that is, the minor radius
        --    MinorRadius is measured along this axis.
        -- Note: This class does not prevent the creation of a
        -- hyperbola where:
        -- -   MajorAxis is equal to MinorAxis, or
        -- -   MajorAxis is less than MinorAxis.
        -- Exceptions
        -- Standard_ConstructionError if MajorAxis or MinorAxis is negative.   
        --     Raises ConstructionError if MajorRadius < 0.0 or MinorRadius < 0.0
      
     raises ConstructionError;
	--- Purpose : Raised if MajorRadius < 0.0 or MinorRadius < 0.0


  SetAxis (me : in out; A1 : Ax1)
        ---C++: inline
        --- Purpose : Modifies this hyperbola, by redefining its local coordinate
        -- system so that:
        -- -   its origin and "main Direction" become those of the
        --   axis A1 (the "X Direction" and "Y Direction" are then
        --   recomputed in the same way as for any gp_Ax2). 
        -- Raises ConstructionError if the direction of A1 is parallel to the direction of
        --  the "XAxis" of the hyperbola.
     raises ConstructionError
      
     is static;


  SetLocation (me : in out; P : Pnt)   is static;
        ---C++: inline
        --- Purpose : Modifies this hyperbola, by redefining its local coordinate
        -- system so that its origin becomes P.
  


  SetMajorRadius (me : in out; MajorRadius : Real)
        ---C++: inline
        --- Purpose:
        -- Modifies the major  radius of this hyperbola.
        -- Exceptions
        -- Standard_ConstructionError if MajorRadius is negative.
     raises ConstructionError
     is static;


  SetMinorRadius (me : in out; MinorRadius : Real)
        ---C++: inline
        --- Purpose:
        -- Modifies the minor  radius of this hyperbola.
        -- Exceptions
        -- Standard_ConstructionError if MinorRadius is negative. 
     raises ConstructionError
     is static;


  SetPosition (me : in out; A2 : Ax2)   is static;
        ---C++: inline
        --- Purpose : Modifies this hyperbola, by redefining its local coordinate
        -- system so that it becomes A2.


  Asymptote1 (me)   returns Ax1
        ---C++: inline
	--- Purpose :
	--  In the local coordinate system of the hyperbola the equation of
	--  the hyperbola is (X*X)/(A*A) - (Y*Y)/(B*B) = 1.0 and the
        --  equation of the first asymptote is Y = (B/A)*X
        --  where A is the major radius and B is the minor radius. Raises ConstructionError if MajorRadius = 0.0
     raises ConstructionError
     is static;


  Asymptote2 (me)   returns Ax1
        ---C++: inline
	--- Purpose :
	--  In the local coordinate system of the hyperbola the equation of
	--  the hyperbola is (X*X)/(A*A) - (Y*Y)/(B*B) = 1.0 and the
        --  equation of the first asymptote is Y = -(B/A)*X.
        --  where A is the major radius and B is the minor radius. Raises ConstructionError if MajorRadius = 0.0
     raises ConstructionError
     is static;


  Axis (me)  returns Ax1  is static;
        ---C++: inline
        --- Purpose : Returns the axis passing through the center,
        -- and normal to the plane of this hyperbola.
    	---C++: return const&

  ConjugateBranch1 (me)  returns Hypr  is static;
        ---C++: inline
	--- Purpose :
	--  Computes the branch of hyperbola which is on the positive side of the 
	--  "YAxis" of <me>.


  ConjugateBranch2 (me)  returns Hypr  is static;
        ---C++: inline
	--- Purpose :
	--  Computes the branch of hyperbola which is on the negative side of the 
	--  "YAxis" of <me>.


  Directrix1 (me)  returns Ax1   is static;
        ---C++: inline
        --- Purpose :
        --  This directrix is the line normal to the XAxis of the hyperbola
        --  in the local plane (Z = 0) at a distance d = MajorRadius / e 
        --  from the center of the hyperbola, where e is the eccentricity of
        --  the hyperbola.
        --  This line is parallel to the "YAxis". The intersection point
        --  between the directrix1 and the "XAxis" is the "Location" point
        --  of the directrix1. This point is on the positive side of the
        --  "XAxis".


  Directrix2 (me)   returns Ax1  is static;
        ---C++: inline
        --- Purpose :
        --  This line is obtained by the symmetrical transformation 
        --  of "Directrix1" with respect to the "YAxis" of the hyperbola.


  Eccentricity (me)   returns Real
        ---C++: inline
	--- Purpose :
	--  Returns the excentricity of the hyperbola (e > 1).
	--  If f is the distance between the location of the hyperbola
	--  and the Focus1 then the eccentricity e = f / MajorRadius. Raises DomainError if MajorRadius = 0.0
     raises DomainError
     is static;


  Focal (me)  returns Real  is static;
        ---C++: inline
	--- Purpose :
	--  Computes the focal distance. It is the distance between the
        --  the two focus of the hyperbola.


  Focus1 (me)   returns Pnt  is static;
        ---C++: inline
	--- Purpose :
	--  Returns the first focus of the hyperbola. This focus is on the
        --  positive side of the "XAxis" of the hyperbola.


  Focus2 (me)   returns Pnt  is static;
        ---C++: inline
        --- Purpose :
	--  Returns the second focus of the hyperbola. This focus is on the
        --  negative side of the "XAxis" of the hyperbola.


  Location (me)    returns Pnt   is static;
        ---C++: inline
        --- Purpose :
        --  Returns  the location point of the hyperbola. It is the
        --  intersection point between the "XAxis" and the "YAxis".
    	---C++: return const&


  MajorRadius (me)  returns Real is static;
        ---C++: inline
	--- Purpose :
	--  Returns the major radius of the hyperbola. It is the radius
	--  on the "XAxis" of the hyperbola.


  MinorRadius (me)   returns Real  is static;
        ---C++: inline
	--- Purpose :
	--  Returns the minor radius of the hyperbola. It is the radius
	--  on the "YAxis" of the hyperbola.


  OtherBranch (me)   returns Hypr is static;
        ---C++: inline
        --- Purpose :
	--  Returns the branch of hyperbola obtained by doing the 
	--  symmetrical transformation of <me> with respect to the 
	--  "YAxis"  of <me>.


  Parameter (me)  returns Real
        ---C++: inline
        --- Purpose :
        --  Returns p = (e * e - 1) * MajorRadius where e is the 
        --  eccentricity of the hyperbola.
        --- Raises DomainError if MajorRadius = 0.0
     raises DomainError
     is static;


  Position (me)   returns Ax2   is static;
        --- Purpose : Returns the coordinate system of the hyperbola.
        ---C++: inline
        ---C++: return const&


  XAxis (me)  returns Ax1    is static;
        ---C++: inline
        --- Purpose : Computes an axis, whose
        -- -   the origin is the center of this hyperbola, and
        -- -   the unit vector is the "X Direction" 
        --   of the local coordinate system of this hyperbola.
        -- These axes are, the major axis (the "X
        -- Axis") and  of this hyperboReturns the "XAxis" of the hyperbola.


  YAxis (me)  returns Ax1    is static;
        ---C++: inline
        --- Purpose :      Computes an axis, whose
        -- -   the origin is the center of this hyperbola, and
        -- -   the unit vector is the "Y Direction"
        --   of the local coordinate system of this hyperbola. 
        -- These axes are the minor axis (the "Y Axis") of this hyperbola

    

  Mirror (me : in out; P : Pnt)          is static;

  Mirrored (me; P : Pnt)   returns Hypr  is static;
        --- Purpose :
        --  Performs the symmetrical transformation of an hyperbola with 
        --  respect  to the point P which is the center of the symmetry.

  Mirror (me : in out; A1 : Ax1)          is static;

  Mirrored (me; A1 : Ax1)   returns Hypr  is static;


        --- Purpose :
        --  Performs the symmetrical transformation of an hyperbola with 
        --  respect to an axis placement which is the axis of the symmetry.

     
  Mirror (me : in out; A2 : Ax2)         is static;

  Mirrored (me; A2 : Ax2)  returns Hypr  is static;
        --- Purpose :
        --  Performs the symmetrical transformation of an hyperbola with
        --  respect to a plane. The axis placement A2 locates the plane 
        --  of the symmetry (Location, XDirection, YDirection).


  Rotate (me : in out; A1 : Ax1; Ang : Real)         is static;
        ---C++: inline
  Rotated (me; A1 : Ax1; Ang : Real)   returns Hypr  is static;
        ---C++: inline
        --- Purpose :
        --  Rotates an hyperbola. A1 is the axis of the rotation.
        --  Ang is the angular value of the rotation in radians.



  Scale (me : in out; P : Pnt; S : Real)         is static;
        ---C++: inline

  Scaled (me; P : Pnt; S : Real)   returns Hypr  is static;
        ---C++: inline
        --- Purpose : 
        --  Scales an hyperbola. S is the scaling value.

  

  Transform (me : in out; T : Trsf)          is static;
        ---C++: inline

  Transformed (me; T : Trsf)   returns Hypr   is static;
        ---C++: inline
        --- Purpose :
        --  Transforms an hyperbola with the transformation T from 
        --  class Trsf.



  Translate (me : in out; V : Vec)         is static;
        ---C++: inline

  Translated (me; V : Vec)  returns Hypr   is static;
        ---C++: inline
        --- Purpose :
        --  Translates an hyperbola in the direction of the vector V.
        --  The magnitude of the translation is the vector's magnitude.


  Translate(me : in out; P1, P2 : Pnt)          is static;
        ---C++: inline

  Translated (me; P1, P2 : Pnt)   returns Hypr  is static;
        ---C++: inline
        --- Purpose :
        --  Translates an hyperbola from the point P1 to the point P2.


fields

     pos         : Ax2;
     majorRadius : Real;
     minorRadius : Real;


end;

