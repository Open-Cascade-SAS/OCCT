-- Created on: 1993-01-09
-- Created by: CKY / Contract Toubro-Larsen ( SIVA )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ToroidalSurface from IGESSolid  inherits IGESEntity

        ---Purpose: defines ToroidalSurface, Type <198> Form Number <0,1>
        --          in package IGESSolid
        --          This entity is defined by the center point, the axis
        --          direction and the major and minor radii. In case of
        --          parametrised surface a reference direction is provided.

uses

        Point           from IGESGeom,
        Direction       from IGESGeom,
        Pnt             from gp

is

        Create returns ToroidalSurface;

        -- Specific Methods pertaining to the class

        Init (me        : mutable;
              aCenter   : Point;
              anAxis    : Direction;
              majRadius : Real;
              minRadius : Real;
              Refdir    : Direction);
        ---Purpose : This method is used to set the fields of the class
        --           ToroidalSurface
        --       - aCenter   : the center point coordinates
        --       - anAxis    : the direction of the axis
        --       - majRadius : the major radius
        --       - minRadius : the minor radius
        --       - Refdir    : the reference direction (parametrised)
        --                     default Null for unparametrised surface

        Center(me) returns Point;
        ---Purpose : returns the center point coordinates of the surface

        TransformedCenter(me) returns Pnt;
        ---Purpose : returns the center point coordinates of the surface
        -- after applying TransformationMatrix

        Axis(me) returns Direction;
        ---Purpose : returns the direction of the axis

        MajorRadius(me) returns Real;
        ---Purpose : returns the major radius of the surface

        MinorRadius(me) returns Real;
        ---Purpose : returns the minor radius of the surface

        ReferenceDir(me) returns Direction;
        ---Purpose : returns the reference direction (parametrised surface)
        -- Null is returned if the surface is not parametrised

        IsParametrised(me) returns Boolean;
        ---Purpose : Returns True if the surface is parametrised, else False

fields

--
-- Class    : IGESSolid_ToroidalSurface
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class ToroidalSurface.
--
-- Reminder : A ToroidalSurface instance is defined by :
--            This entity is defined by the center point, the axis
--            direction and the major and minor radii. In case of
--            parametrised surface a reference direction is provided.
--

        theCenter      : Point;
            -- the center point coordinates of the surface

        theAxis        : Direction;
            -- the direction of the axis

        theMajorRadius : Real;
            -- the major radius of the surface

        theMinorRadius : Real;
            -- the minor radius of the surface

        theRefDir      : Direction;
            -- the reference direction of the surface (parametrised)

end ToroidalSurface;
