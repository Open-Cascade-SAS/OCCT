-- Created on: 2009-04-06
-- Created by: Sergey ZARITCHNY
-- Copyright (c) 2009-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


deferred class Pattern from TDataXtd inherits Attribute from TDF

	---Purpose: a general pattern model

uses 
     Array1OfTrsf from TDataXtd,
     LabelList    from TDF,
     GUID         from Standard

is

    GetID (myclass)   
    ---C++: return const &  
    returns GUID from Standard;    
   
    ID(me)
    	returns GUID from Standard
	is redefined static;
	---Purpose: Returns the ID of the attribute.
	--          
	---C++: return const &

    PatternID(me)
    	returns GUID from Standard
	is deferred;
	---Purpose: Returns the ID of the attribute.
	--          
	---C++: return const &

    NbTrsfs(me)
    returns Integer from Standard
    is deferred;
        ---Purpose: Give the number of transformation

    ComputeTrsfs(me; Trsfs : in out Array1OfTrsf from TDataXtd)
    is deferred;
        ---Purpose: Give the transformations

end Pattern;


