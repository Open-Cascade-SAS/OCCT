-- File:	StepToGeom_MakeToroidalSurface.cdl
-- Created:	Mon Jun 14 16:23:51 1993
-- Author:	Martine LANGLOIS
---Copyright:	 Matra Datavision 1993

class MakeToroidalSurface from StepToGeom

    ---Purpose: This class implements the mapping between class
    --          ToroidalSurface from StepGeom which describes a
    --          toroidal_surface from Prostep and ToroidalSurface from Geom 
  
uses ToroidalSurface from Geom,
     ToroidalSurface from StepGeom
     
is 

    Convert ( myclass; SS : ToroidalSurface from StepGeom;
                       CS : out ToroidalSurface from Geom )
    returns Boolean from Standard;
    
end MakeToroidalSurface;
