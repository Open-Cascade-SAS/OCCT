-- File:        OffsetCurve3d.cdl
-- Created:     Mon Dec  4 12:02:28 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWOffsetCurve3d from RWStepGeom

	---Purpose : Read & Write Module for OffsetCurve3d

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     OffsetCurve3d from StepGeom,
     EntityIterator from Interface

is

	Create returns RWOffsetCurve3d;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable OffsetCurve3d from StepGeom);

	WriteStep (me; SW : in out StepWriter; ent : OffsetCurve3d from StepGeom);

	Share(me; ent : OffsetCurve3d from StepGeom; iter : in out EntityIterator);

end RWOffsetCurve3d;
