-- Created on: 2001-04-05
-- Created by: Peter KURNEV
-- Copyright (c) 2001-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Tools3D from BOPTools

	---Purpose:  
	--  The class contains handy static functions 
	--  dealing with the topology 

uses  
    Pln   from gp, 
    Dir   from gp, 
    Pnt   from gp,   
    Pnt2d from gp,  
    
    Surface from Geom,
    
    Shape from TopoDS, 
    Wire  from TopoDS, 
    Face  from TopoDS,  
    Edge  from TopoDS,
    Solid from TopoDS,
     
    ShapeEnum   from TopAbs,     
    Orientation from TopAbs, 
    State       from TopAbs, 

    ListOfShape from TopTools, 
    Context     from IntTools, 

    IndexedDataMapOfShapeListOfShape from TopTools

is  

    SubShapesAmount        (myclass;  
    	    	    aS:  Shape from TopoDS; 
    	    	    aT:  ShapeEnum from TopAbs) 
    	returns Integer from Standard ;  
    	---Purpose:   
    	-- Returns amount of sub-shapes of type <aT> 
    	-- for the shape <aS> 
    	--
    IsConvexWire            (myclass;   
    	    	    aW:  Wire from TopoDS) 
    	returns Boolean from Standard ;   
    	---Purpose:   
    	-- Returns TRUE if  
    	-- amount of the vertices <=  amount of the edges> 
    	-- for the wire <aW> 
    	--

    RemoveSims  (myclass;    
    	    	    aF:  Face from TopoDS; 
    	    	    aContext: Context from IntTools); 
    	---Purpose: 
    	-- Remove seam edges from face <aF> 
    	--
    RemoveSims  (myclass;    
    	    	    aS:  Shape from TopoDS; 
    	    	    aContext: Context from IntTools); 
    	---Purpose: 
    	-- Remove seam edges from all faces of shape <aS> 
    	--
    EdgeOrientation  (myclass;  
		    aEx:  Edge from TopoDS; 	     
    	    	    aF1:  Face from TopoDS;   
    	    	    aF2:  Face from TopoDS) 
    	returns Orientation from TopAbs;   
    	---Purpose: 
    	-- For the draft section edge <aEx> computes orientation 
    	-- in accordance with vector product between normals to 
    	-- the faces <aF1>,  <aF2> 
    	--
    IsSplitToReverse1  (myclass;  
		    aE1:  Edge from TopoDS; 	     
		    aE2:  Edge from TopoDS; 
    	    	    aContext: Context from IntTools) 
    	returns Boolean from Standard;
    	---Purpose:  
    	-- Returns TRUE if direction of the edge  <aE1> is not           	     
    	-- the same as for the edge <aE2>   	     
    	-- (using  projection) 
    	--
    DoSplitSEAMOnFace (myclass;  
		    aSp:  Edge from TopoDS; 	     
		    aF :  Face from TopoDS);
    	---Purpose:  
    	-- Make the edge <aSp> seam edge for the face <aF>               	     
    	--
	
    --modified by NIZHNY-MKK  Mon Feb 17 15:02:01 2003.BEGIN
    DoSplitSEAMOnFace (myclass;  
			theSplit  :  Edge from TopoDS;
			theSeam   :  Edge from TopoDS;
		    	theFace   :  Face from TopoDS;
    	    	    	IsReversed: out Boolean from Standard)
    	returns Boolean from Standard;
    	---Purpose:  
    	-- Make the edge <theSplit> seam edge for the face <theFace>
    	-- It uses pcurves of <theSeam> to make <theSplit> seam edge.
	-- IsReversed is true if pcurves of <theSplit> and <theSeam> are
	-- reversed according to each other.
	-- Returns true if <theSplit> was made seam edge for <theFace>
	--
    --modified by NIZHNY-MKK  Mon Feb 17 15:02:04 2003.END
    IsTouchCase  (myclass;  
		    aEx:  Edge from TopoDS; 	     
    	    	    aF1:  Face from TopoDS;   
    	    	    aF2:  Face from TopoDS) 
    	returns Boolean from Standard; 
    	---Purpose:  
    	-- Returns TRUE if the edge  <aEx> is section edge           	     
    	-- between touching faces  <aF1>, <aF2>    	     
    	--
    GetTangentToEdge (myclass;  
		    aE:  Edge from TopoDS; 	     
    	    	    aT:  Real from Standard; 
    	    	    aD:out Dir from gp) 
    	returns Boolean from Standard;   
    	---Purpose:   
    	-- Computes tangent (3D) for the edge <aE>  
    	-- at parameter <aT>           
    	-- Returns TRUE if the edge <aE> is not degenerated. 
    	--
    GetTangentToEdge (myclass;  
		    aE:  Edge from TopoDS; 	     
    	    	    aD:out Dir from gp) 
    	returns Boolean from Standard;    
    	---Purpose:  
    	--- Computes tangent (3D) for the edge <aE>  
    	--- at arbitrary intermediate parameter           
    	--- Returns TRUE if the edge <aE> is not degenerated. 
    	---
    GetNormalToFaceOnEdge (myclass;  
		    aE:  Edge from TopoDS; 	     
    	    	    aF:  Face from TopoDS;   
    	    	    aT:  Real from Standard; 
    	    	    aD:out Dir from gp); 
    	---Purpose:  
    	--- Computes normal to the face <aF> for the point on the edge <aE>  
    	--- at parameter <aT>           
    	---
    GetNormalToFaceOnEdge (myclass;  
		    aE:  Edge from TopoDS; 	     
    	    	    aF:  Face from TopoDS;   
    	    	    aD:out Dir from gp); 	 
    	---Purpose:  
    	--- Computes normal to the face <aF> for the point on the edge <aE>  
    	--- at arbitrary intermediate parameter 
    	---
    GetBiNormal (myclass;  
		    aE:  Edge from TopoDS; 	     
    	    	    aF:  Face from TopoDS; 
                    aT:  Real from Standard;    				 
    	    	    aD:out Dir from gp);  
    	---Purpose:   
    	--- Computes binormal to the face <aF> for the point on the edge <aE>  
    	--- at parameter <aT>           
    	---
    GetBiNormal (myclass;  
		    aE:  Edge from TopoDS; 	     
    	    	    aF:  Face from TopoDS;   
    	    	    aD:out Dir from gp); 
    	---Purpose:   
    	--- Computes binormal to the face <aF> for the point on the edge <aE>  
    	--- at arbitrary intermediate parameter            
    	---
    IsSplitToReverse(myclass;  
		    aE :  Edge from TopoDS; 
		    aSp:  Edge from TopoDS) 
    	returns Boolean from Standard; 
    	---Purpose:  
    	--- Returns TRUE if direction of the edge  <aE1> is not           	     
    	--- the same as for the edge <aE2>   	     
    	---
    GetAdjacentFace (myclass;  
		    aF :  Face from TopoDS;
		    aE :  Edge from TopoDS; 
		    aEFMap: IndexedDataMapOfShapeListOfShape from TopTools; 
		    anAdjF:out Face from TopoDS) 
	returns Boolean from Standard;  
    	---Purpose: 
    	--- Get face <anAdjF> that  is adjacent to the face <aF> through 
    	--- the edge <aE>  (using map EF <aEFMap>) 
    	--- Returns FALSE if adjacent face is not found 
    	---
    IsKeepTwice  (myclass;  
		    aF1   :  Face from TopoDS;
		    aF2   :  Face from TopoDS;
		    aF2Adj:  Face from TopoDS;
		    aSpEF2:  Edge from TopoDS) 
	returns Boolean from Standard;  
    	---Purpose: 
    	--- Returns TRUE if pair of faces <aF2> and <aF2Adj> 
    	--- that are adjacent faces through the edge <aSpEF2> 
    	--- crosses the face <aF1> by <aSpEF2> 
    	---
    SenseFlag    (myclass;  
		    aNF1   :  Dir from gp;
		    aNF2   :  Dir from gp) 
	returns Integer from Standard;   
    	---Purpose: 
    	--- Returns 1  if scalar product aNF1* aNF2>0.   
    	--- Returns 0  if directions aNF1 aNF2 coinside  
    	--- Returns -1 if scalar product aNF1* aNF2<0.      
    	---
    GetNormalToSurface    (myclass;  
		    aS:  Surface from Geom; 
		    U :  Real from Standard;
		    V :  Real from Standard; 
    	    	    aD:out Dir from gp)
	returns Boolean from Standard;   
    	---Purpose:  
    	--- Compute normal <aD> to surface <aS> in point (U,V)  
    	--- Returns TRUE if directions aD1U, aD1V coinside 
    	---
    GetPlanes     (myclass;  
		    aSp :  Edge from TopoDS;
		    aE2 :  Edge from TopoDS; 
		    aEFMap2: IndexedDataMapOfShapeListOfShape from TopTools; 
    	    	    aE1 :  Edge from TopoDS; 
    	    	    aF1 :  Face from TopoDS; 
    	    	    aST1:out State from TopAbs; 
    	    	    aContext: Context from IntTools); 
    	---Purpose: 
    	--- Internal usage 
    	---
    Orientation  (myclass;  
		    aE :  Edge from TopoDS; 
    	    	    aF :  Face from TopoDS) 
    	returns Orientation from TopAbs;  
    	---Purpose: 
    	--- Get the orientation for the edge <aE> on the face <aF> 
    	--- Returns  TopAbs_INTERNAL if  the edge <aE> is not found 
    	--- on the face <aF> 
    	---
    SignDistance (myclass; 
     	    	    aP :  Pnt  from  gp; 
    	    	    aPL:  Pln  from  gp) 
	 returns Real from Standard; 
    	---Purpose: 
    	--- Computes signed distance between the 3D-point <aP> 
    	--- and the plane <aPL>.   
	---
	--  Warning:
    	--- The distance is not divided by sqrt(A*A+B*B+C*C) 
    	---
    GetApproxNormalToFaceOnEdge (myclass;  
		    aE:  Edge from TopoDS; 	     
    	    	    aF:  Face from TopoDS;   
    	    	    aT:  Real from Standard;  
    	    	    aPx:out Pnt from gp;
    	    	    aD:out Dir from gp); 
    	---Purpose:  
    	--- Computes normal to the face <aF> for the 3D-point that 
    	--- belonds to the edge <aE> at parameter <aT>. 
    	--  Output: 
    	--- aPx  -  the 3D-point where the normal computed 
    	--- aD   -  the normal; 
    	---
	--  Warning:
    	--- The normal is computed not exactly in the point on the 
    	--- edge, but in point that is near to the edge towards to 
    	--- the face material (so, we'll have approx. normal) 
    	---
    PointNearEdge   (myclass;   
     	    	    aE   :  Edge from TopoDS; 	     
    	    	    aF   :  Face from TopoDS;   
        	    aT   :  Real from Standard;  
	    	    aDt2D:  Real from Standard;  
		    aP2D :out Pnt2d from  gp; 
    	    	    aPx  :out Pnt from gp);  
    	---Purpose: 
    	--- Compute the point <aPx>,  (<aP2D>)  that is near to  
    	--- the edge <aE>   at parameter <aT>  towards to the  
    	--- material of the face <aF>. The value of shifting in 
    	--- 2D is <aDt2D> 
    	---
    PointNearEdge   (myclass;   
     	    	    aE:  Edge from TopoDS; 	     
    	    	    aF:  Face from TopoDS;   
    	    	    aT:  Real from Standard;  
		    aP2D:out Pnt2d from  gp; 
    	    	    aPx:out Pnt from gp);  
    	---Purpose: 
    	--- Computes the point <aPx>,  (<aP2D>)  that is near to  
    	--- the edge <aE>   at parameter <aT>  towards to the  
    	--- material of the face <aF>. The value of shifting in 
    	--  2D is  dt2D=BOPTools_Tools3D::MinStepIn2d()
    	---
    PointNearEdge   (myclass;   
     	    	    aE:  Edge from TopoDS; 	     
    	    	    aF:  Face from TopoDS;   
		    aP2D:out Pnt2d from  gp; 
    	    	    aPx:out Pnt from gp);   
    	---Purpose: 
    	--- Compute the point <aPx>,  (<aP2D>)  that is near to  
    	--- the edge <aE>   at arbitrary  parameter  towards to the  
    	--- material of the face <aF>. The value of shifting in 
    	--  2D is  dt2D=BOPTools_Tools3D::MinStepIn2d()
    	---
    PointToCompare (myclass; 
    		    aP1: Pnt from gp;	    
    		    aP2: Pnt from gp; 
                    aF:  Face from TopoDS;     		    				 
    		    aPx:out Pnt from gp; 
    	    	    aContext:  Context from IntTools);  
    	---Purpose: 
    	--- For 3D-point <aP1> find projection point <aPx> on the face <aF>. 
    	--- If the distance  (<aP1>, <aPx>) > TolF => 
    	--- For 3D-point <aP2> find projection point <aPx> on the face <aF>.    
    	--- If the distance  (<aP2>, <aPx>) > TolF => returns <aP1> 
    	---
    GetPlane       (myclass;  
		    aSp :  Edge from TopoDS;
    	    	    aE1 :  Edge from TopoDS; 
    	    	    aF1 :  Face from TopoDS; 
    	    	    aF2 :  Face from TopoDS; 
    	    	    aST:out State from TopAbs; 
    	    	    aContext: Context from IntTools); 
    	---Purpose:  
    	--- Compute 3D-state for the point on the split edge <aSp>  
    	--- (with base edge <aE1> and the face <aF1>) comparing with 
    	--- the face <aF2> 
    	---
    GetPointState  (myclass;  
		    aSp    :  Edge from TopoDS;
    	    	    aEF2   :  Edge from TopoDS; 
    	    	    aF2Adj :  Face from TopoDS; 
    	    	    aF1    :  Face from TopoDS; 
    	    	    aST:out State from TopAbs);  
    	---Purpose:  
    	--- Compute 3D-state for the point on the split edge <aSp>  
    	--- (with base edge <aEF2> and the adjacent face <aF2Adj>) comparing with 
    	--- the face <aF1> 
    	---
    	 
    OrientEdgeOnFace  (myclass;  
		    aE    :  Edge from TopoDS;
    	    	    aF    :  Face from TopoDS;  
    	    	    aER   : out  Edge from TopoDS); 
    	---Purpose:  
    	--- Get the edge <aER> from the face <aF> that is the same as   
    	--- the edge <aE>    
    	---

    OrientTouchEdgeOnF1  (myclass;    
    	    	    aSp:  Edge from TopoDS; 	     
    	    	    aEx:  Edge from TopoDS; 	     
    	    	    aF1:  Face from TopoDS;   
    	    	    aF2:  Face from TopoDS) 
    	returns Orientation from TopAbs;    
    	---Purpose: 
    	--- Computes orientation for the split edge <aSp>   
    	--- [with base edge <aEx> and face <aF2>] on the 
    	--- face <aF1> 
    	---
    GetSeams  (myclass;  
    	    	    aF    :  Face from TopoDS;  
    	    	    aSimm1   : out  Edge from TopoDS;
    	    	    aSimm2   : out  Edge from TopoDS); 
    	---Purpose:  
    	--- Get seam edges <aSimm1>, <aSimm2> for the face <aF> 
    	---
    GetSeam   (myclass;  
    	    	    aF    :  Face from TopoDS;  
    	    	    aS1:  Edge from TopoDS;
    	    	    aS2: out  Edge from TopoDS);   	
    	---Purpose:  
    	--- Get opposite seam edge <aS2> for the face <aF> with 
    	--- known  seam edge <aS1>  
    	---
    IsValidArea   (myclass;   
    	    	    aF            :  Face from TopoDS; 
    	    	    aNegativeFlag :  out Boolean from Standard) 
    	returns  Boolean from Standard;  
    	---Purpose:  
    	--- Check validity of the area of face <aF>.  
    	--- Returns TRUE if the Abs. value of the area 
    	--- is greater than  1.e-16 
    	---
    MinStepIn2d(myclass) 
    	returns  Real from Standard;  
    	---Purpose:  
    	--- Returns simple step value that is used in 2D-computations 
    	--- = 1.e-5 
    	---
    IsEmptyShape(myclass; 
    	            aS:  Shape from TopoDS) 
	returns Boolean from Standard; 
    	---Purpose: 
    	--- Returns TRUE if the shape <aS> does not contain 
    	--- geometry information  (e.g. empty compound) 
    	---
    InvertShape(myclass; 
    	            aS   :    Shape from TopoDS; 
    	            aSInv:out Shape from TopoDS);  
    	---Purpose:  
    	--- Change orientations to opposite for the shape <aS> 
    	--- and all its sub-shapes. Returns <aSInv>        
    	---
    GetStatePartIN2D(myclass; 	 
	     aSp    :Edge from TopoDS; 
	     aEF1   :Edge from TopoDS; 
	     aF1    :Face from TopoDS; 	
	     aF2    :Face from TopoDS; 
    	     aContext:  Context from IntTools)
    	returns  State from TopAbs;  
    	---Purpose: 
    	--- Used in touch case          
    	--- Compute the 3D-state for the point on the split 
    	--- edge <aSp> (with base edge <aEF1> on face <aF1>) 
    	--- comparing with <aF2>.   
    	--- Used in touch case  <aF1>/<aF2> 
    	---
    CheckSameDomainFaceInside(myclass; theFace1: Face from TopoDS;
    	    	    	    	       theFace2: Face from TopoDS;
    	    	    	    	       theContext: Context from IntTools)
    	returns Boolean from Standard;

    ComputeFaceState(myclass; theFace: Face from TopoDS;
    	    	    	      theRef : Solid from TopoDS;
    	    	    	      theContext: Context from IntTools;
			      theState: out State from TopAbs)
    	returns Boolean from Standard;

    TreatedAsAnalytic(myclass; aTx    :Real from Standard; 
	    		       aPx    :Pnt  from gp;    
	    	    	       aEx    :Edge from TopoDS; 
    	    	    	       aFx    :Face from TopoDS; 
    	     	    	       aE1    :Edge from TopoDS; 
	     	    	       aF1    :Face from TopoDS;   
             	    	       aTolTangent:Real from Standard; 	      
             	    	       aTolRadius :Real from Standard; 	      
    	     	    	       aState  :out State from TopAbs;     	
    	     	    	       aContext: Context from IntTools)
    	returns  Boolean from Standard;  

    TreatedAsAnalytic (myclass; aFx    :Face from TopoDS; 
    	     	    	    	aSpE1  :Edge from TopoDS; 
    	    	    	    	aF1    :Face from TopoDS; 
    	     	    	    	aTolTangent:Real from Standard; 	      
             	    	    	aTolRadius :Real from Standard;  
    	     	    	    	aState  :out State from TopAbs;     	
    	     	    	    	aContext: Context from IntTools)
    	returns  Boolean from Standard;   

    HasAnalyticSurfaceType (myclass; aF: Face from TopoDS)  
    	returns  Boolean from Standard; 

end Tools3D;



