-- Created on: 1996-08-27
-- Created by: Philippe MANGIN
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class Approx from AppBlend


	---Purpose: Bspline approximation of a surface.

uses Array2OfPnt             from TColgp,
     HArray2OfPnt            from TColgp,
     Array2OfReal            from TColStd,
     HArray2OfReal           from TColStd,
     Array1OfReal            from TColStd,
     HArray1OfReal           from TColStd,
     Array1OfInteger         from TColStd,
     HArray1OfInteger        from TColStd,
     Array1OfPnt2d           from TColgp

raises NotDone     from StdFail,
       DomainError from Standard,
       OutOfRange  from Standard

is

    IsDone(me)
        returns Boolean from Standard	
	is deferred;


    SurfShape(me; UDegree,VDegree  : out Integer from Standard;
                  NbUPoles,NbVPoles: out Integer from Standard;
                  NbUKnots,NbVKnots: out Integer from Standard)
    	raises NotDone from StdFail
    	is deferred;


    Surface(me; TPoles          : out Array2OfPnt from TColgp;
    	        TWeights        : out Array2OfReal from TColStd;
		TUKnots,TVKnots : out Array1OfReal from TColStd;
		TUMults,TVMults : out Array1OfInteger from TColStd)
    	raises NotDone from StdFail
    	is deferred;


    UDegree(me)
    
    	returns Integer from Standard
    	raises NotDone from StdFail
	is deferred;


    VDegree(me)
    
    	returns Integer from Standard
    	raises NotDone from StdFail
	is deferred;


    SurfPoles(me)
    
    	returns Array2OfPnt from TColgp
	---C++: return const&

	raises NotDone from StdFail
	is deferred;


    SurfWeights(me)
    
    	returns Array2OfReal from TColStd
	---C++: return const&

	raises NotDone from StdFail
	is deferred;


    SurfUKnots(me)
    
    	returns Array1OfReal from TColStd
	---C++: return const&

	raises NotDone from StdFail
	is deferred;


    SurfVKnots(me)
    
    	returns Array1OfReal from TColStd
	---C++: return const&

	raises NotDone from StdFail
	is deferred;


    SurfUMults(me)
    
    	returns Array1OfInteger from TColStd
	---C++: return const&

	raises NotDone from StdFail
	is deferred;


    SurfVMults(me)
    
    	returns Array1OfInteger from TColStd
	---C++: return const&

	raises NotDone from StdFail
	is deferred;


    NbCurves2d(me)
    
    	returns Integer from Standard	
	raises NotDone from StdFail
	is deferred;


    Curves2dShape(me; Degree,NbPoles,NbKnots: out Integer from Standard)
    
    	raises NotDone from StdFail,
	       DomainError from Standard

        is deferred;
	
	
    Curve2d(me; Index: Integer from Standard;
                TPoles   : out Array1OfPnt2d from TColgp;
		TKnots   : out Array1OfReal from TColStd;
		TMults   : out Array1OfInteger from TColStd)
		
    	raises NotDone     from StdFail,
	       OutOfRange  from Standard,
	       DomainError from Standard

    	is deferred;     


    Curves2dDegree(me)
    
    	returns Integer from Standard	
	raises NotDone from StdFail,
	       DomainError from Standard
	is deferred;
	
	
    Curve2dPoles(me; Index: Integer from Standard)
    
    	returns Array1OfPnt2d from TColgp
	---C++: return const&
	
	raises NotDone     from StdFail,
	       OutOfRange  from Standard,
	       DomainError from Standard
	is deferred;
	

    Curves2dKnots(me)
    
    	returns Array1OfReal from TColStd
	---C++: return const&

	raises NotDone from StdFail,
	       DomainError from Standard
	is deferred;


    Curves2dMults(me)
    
    	returns Array1OfInteger from TColStd
	---C++: return const&

	raises NotDone from StdFail,
	       DomainError from Standard
	is deferred;
	
    TolReached(me; Tol3d, Tol2d : out Real from Standard)
	raises NotDone from StdFail
	is deferred; 
	 
    TolCurveOnSurf(me; Index  :  Integer  from Standard) 
	returns  Real from Standard  
	raises NotDone from StdFail
        is deferred;    
                    
    ---C++: alias "  Standard_EXPORT virtual ~AppBlend_Approx();"

end Approx;
