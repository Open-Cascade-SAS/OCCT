-- Created on: 1993-01-21
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class WireExplorer from BRepTools

	---Purpose: The WireExplorer is a tool to explore the edges of
	--          a wire in a connection order.
	--          
	--          i.e. each edge is connected to the previous one by
	--          its origin.
	--      If a wire is not closed returns only a segment of edges which
-- length depends on started in exploration edge. If wire has
-- singularities (for example, loops) WireExplorer can return not all
-- edges in a wire. it depends on type of singularity.

uses

    Orientation from TopAbs,
    Wire        from TopoDS,
    Edge        from TopoDS,
    Vertex      from TopoDS,
    Face        from TopoDS,
    DataMapOfShapeListOfShape from TopTools,
    MapOfShape                from TopTools
raises
    DomainError  from Standard,
    NoSuchObject from Standard,
    NoMoreObject from Standard

is
    Create returns WireExplorer from BRepTools;
---Purpose: Constructs an empty explorer (which can be initialized using Init)
    
    Create(W : Wire from TopoDS ) returns WireExplorer from BRepTools
	---Purpose: IInitializes an exploration  of the wire <W>. 
    raises DomainError from Standard;
    
    Create(W : Wire from TopoDS;
    	   F : Face from TopoDS) returns WireExplorer from BRepTools
	---Purpose: Initializes an exploration  of the wire <W>.
	--          F is used to select the edge connected to the 
	--          previous in the parametric representation of <F>.
    raises DomainError from Standard;

    Init(me : in out; W  : Wire from TopoDS)
	---Purpose: Initializes an exploration of the wire <W>.
    raises DomainError from Standard
    is static;
    
    Init(me : in out; W  : Wire from TopoDS;
    	    	      F  : Face from TopoDS)
	---Purpose: Initializes an exploration of the wire <W>.
	--          F is used to select the edge connected to the 
	--          previous in the parametric representation of <F>.
	--          
    raises DomainError from Standard
    is static;
    
    More(me) returns Boolean
	---Purpose: Returns True if there  is a current  edge.
    is static;
    
    Next(me : in out)
	---Purpose: Proceeds to the next edge.
    raises
	NoMoreObject from Standard 
    is static;
    
    Current(me) returns Edge from TopoDS
	---Purpose: Returns the current edge. 
    raises
    	NoSuchObject from Standard
	---C++: return const &
    is static;
    
    Orientation(me) returns Orientation from TopAbs
	---Purpose: Returns an Orientation for the current edge.
    is static;
    
    CurrentVertex(me) returns Vertex from TopoDS
	---Purpose: Returns the vertex connecting the current  edge to
	--          the previous one.
    raises
    	NoSuchObject from Standard
	--          
	---C++: return const &
    is static;
    
   Clear(me : in out)
	---Purpose: Clears the content of the explorer.
    is static;
    
fields
    myMap    : DataMapOfShapeListOfShape from TopTools;
    myEdge   : Edge   from TopoDS;
    myVertex : Vertex from TopoDS;
    myFace   : Face   from TopoDS;
    myDoubles: MapOfShape from TopTools;
    myReverse: Boolean from Standard; 
    myTolU   : Real  from  Standard; 
    myTolV   : Real  from  Standard; 

end WireExplorer;
