-- Created on: 1995-06-14
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class FaceEdgeFiller from TopOpeBRep

uses

    Shape                      from TopoDS,
    FaceEdgeIntersector              from TopOpeBRep,
    HDataStructure                   from TopOpeBRepDS,
    DataStructure                               from TopOpeBRepDS,
    Interference                     from TopOpeBRepDS,
    ListOfInterference               from TopOpeBRepDS,    
    ListIteratorOfListOfInterference from TopOpeBRepDS,
    Point                            from TopOpeBRepDS
    
is 

    Create returns FaceEdgeFiller from TopOpeBRep;
    
    Insert(me : in out;
    	   F,E : Shape from TopoDS;
    	   FEINT : in out FaceEdgeIntersector from TopOpeBRep;
	   HDS : HDataStructure from TopOpeBRepDS)
    is static;

    -- -------
    -- private
    -- -------

    ScanInterfList(me; 
    	IT : in out ListIteratorOfListOfInterference from TopOpeBRepDS;
	DSP : Point from TopOpeBRepDS;
	BDS : DataStructure from TopOpeBRepDS)
    ---Purpose: 
    -- Search, among a list of interferences accessed by the iterator
    -- <IT>, a geometry <G> whose 3D point is identical to the 3D point
    -- of the TheDSPoint <DSP>.
    -- returns True if such an interference has been found, False else.
    -- if True, iterator It points (by the Value() method) on the first 
    -- interference accessing an identical 3D point.
	
    returns Boolean from Standard
    is static private;

    GetGeometry(me ; 
         IT : in out ListIteratorOfListOfInterference from TopOpeBRepDS;
	 EI : FaceEdgeIntersector from TopOpeBRep;
	 G  : in out Integer from Standard;
    	 DS : DataStructure from TopOpeBRepDS)
    ---Purpose:
    -- Search for an interference in list <IT> which 3D geometry 
    -- equals 3D geometry of the current intersection of <EI>.
    -- The search is performed by ScanInterfList.
    -- if found, set <G> to the geometry of the interference found.
    -- returns found.
	
    returns Boolean from Standard
    is static private;

    MakeGeometry(me ; EI : in out FaceEdgeIntersector from TopOpeBRep;
    	    	      DS  : in out DataStructure from TopOpeBRepDS)
    returns Integer from Standard
    is static private;

    GetGeometry(me ; L   : ListOfInterference from TopOpeBRepDS;
		     DSP : Point from TopOpeBRepDS;
		     G   : in out Integer from Standard;
    	    	     DS  : in out DataStructure from TopOpeBRepDS)
    ---Purpose:
    -- Get the geometry of a DS point <DSP>.
    -- First, search it with ScanInterfList (previous method).
    -- if found, set <G> to the geometry of the interference found.
    -- else, add the point <DSP> in the <DS> and set <G> to the 
    -- value of the new geometry such created.
    -- 
    -- returns the value of ScanInterfList().
	
    returns Boolean from Standard
    is static private;


    StoreInterference(me; 
    	    	      I   : Interference from TopOpeBRepDS;
    	    	      LI  : in out ListOfInterference from TopOpeBRepDS;
		      BDS : in out DataStructure from TopOpeBRepDS)
    ---Purpose: 
    -- Add interference <I> to list <LI>.
    -- Add <I> to the interference list of <I> geometry (via <BDS>).
    is static private;
        
end FaceEdgeFiller from TopOpeBRep;
