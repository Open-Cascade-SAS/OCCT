-- Created on: 2000-10-20
-- Created by: Julia DOROVSKIKH
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MidPointRelation from AIS inherits Relation from AIS

	---Purpose: presentation of equal distance to point myMidPoint

uses
    ExtendedString        from TCollection,
    Projector             from Prs3d,
    Presentation          from Prs3d,
    PresentationManager3d from PrsMgr,
    Selection             from SelectMgr,
    Dir                   from gp,
    Pnt                   from gp,
    Lin                   from gp,
    Circ                  from gp,
    Elips                 from gp,
    Plane                 from Geom,
    Transformation        from Geom,
    Shape                 from TopoDS

is
    Create(aSymmTool   : Shape from TopoDS;
    	   FirstShape  : Shape from TopoDS;
    	   SecondShape : Shape from TopoDS;
	   aPlane      : Plane from Geom)
    returns mutable MidPointRelation from AIS;

    IsMovable(me) returns Boolean from Standard 
    ---C++: inline       
    is redefined;        

    SetTool(me: mutable; aMidPointTool : Shape from TopoDS);
    ---C++: inline

    GetTool(me)
    ---C++: inline
    ---C++: return const &
    returns Shape from TopoDS;

-- Methods from PresentableObject
    Compute(me: mutable;
  	    aPresentationManager: PresentationManager3d from PrsMgr;
    	    aPresentation       : mutable Presentation from Prs3d;
    	    aMode               : Integer from Standard= 0) 
    is redefined static private;

    Compute(me: mutable;
    	    aProjector   : Projector from Prs3d;
            aPresentation: mutable Presentation from Prs3d)
    is redefined static private;     

    Compute(me: mutable;
    	    aProjector    : Projector from Prs3d;
    	    aTrsf         : Transformation from Geom;
	    aPresentation : mutable Presentation from Prs3d)
    is redefined;
    ---Purpose: Computes the presentation according to a point of view
    --          given by <aProjector>. 
    --          To be Used when the associated degenerated Presentations 
    --          have been transformed by <aTrsf> which is not a Pure
    --          Translation. The HLR Prs can't be deducted automatically
    --          WARNING :<aTrsf> must be applied
    --           to the object to display before computation  !!!

-- Methods from SelectableObject
    ComputeSelection(me         : mutable;
    	    	     aSelection : mutable Selection from SelectMgr;
    	    	     aMode      : Integer from Standard)is private;

-- Computation private methods
    ComputeFaceFromPnt(me: mutable; aprs : mutable Presentation from Prs3d; first : Boolean from Standard)
    is private;

    ComputeEdgeFromPnt(me: mutable; aprs : mutable Presentation from Prs3d; first : Boolean from Standard)
    is private;

    ComputeVertexFromPnt(me: mutable; aprs : mutable Presentation from Prs3d; first : Boolean from Standard)
    is private;

   
    ComputePointsOnLine(me: mutable; aLin : Lin from gp;
    	    	    	    	     first : Boolean from Standard)
    is private;

    ComputePointsOnLine(me: mutable; pnt1,pnt2 : Pnt from gp;
    	    	    	    	     first : Boolean from Standard)
    is private;

    ComputePointsOnCirc(me: mutable; aCirc : Circ from gp; pnt1,pnt2 : Pnt from gp;
    	    	    	    	     first : Boolean from Standard)
    is private;

    ComputePointsOnElips(me: mutable; anEll : Elips from gp; pnt1,pnt2 : Pnt from gp;
    	    	    	    	      first : Boolean from Standard)
    is private;
    ---Purpose: ComputePointsOn... methods set myFAttach, myFirstPnt and myLastPnt
    -- from the following initial data: curve, end points, myMidPoint.
    -- End points (pnt1 & pnt2) and curve define the trimmed curve.
    -- If end points are equal, curve is not trimmed (line - special case).
    -- 
    --     .------. pnt2
    --    /        \
    --   .  circle  . myLastPnt
    --   |          |
    --   . pnt1     . myFAttach
    --    \   arc  /          . myMidPoint
    --     .______. myFirstPnt
fields
    myTool     : Shape from TopoDS;
    myMidPoint : Pnt   from gp; -- point of symmetry

    myFAttach  : Pnt   from gp; -- position on myFShape to be connected with myMidPoint by segment
    myFirstPnt1 : Pnt   from gp; -- points on myFShape,
    myFirstPnt2 : Pnt   from gp; -- defining a segment of it to be drawn

    mySAttach  : Pnt   from gp; -- position on mySShape to be connected with myMidPoint by segment
    mySecondPnt1  : Pnt   from gp; -- points on mySShape,
    mySecondPnt2  : Pnt   from gp; -- defining a segment of it to be drawn

end MidPointRelation;
