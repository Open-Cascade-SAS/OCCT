-- File:	StepRepr_AssemblyComponentUsage.cdl
-- Created:	Mon Jul  3 19:47:50 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class AssemblyComponentUsage from StepRepr
inherits ProductDefinitionUsage from StepRepr

    ---Purpose: Representation of STEP entity AssemblyComponentUsage

uses
    HAsciiString from TCollection,
    ProductDefinition from StepBasic

is
    Create returns AssemblyComponentUsage from StepRepr;
	---Purpose: Empty constructor

    Init (me: mutable; aProductDefinitionRelationship_Id: HAsciiString from TCollection;
                       aProductDefinitionRelationship_Name: HAsciiString from TCollection;
                       hasProductDefinitionRelationship_Description: Boolean;
                       aProductDefinitionRelationship_Description: HAsciiString from TCollection;
                       aProductDefinitionRelationship_RelatingProductDefinition: ProductDefinition from StepBasic;
                       aProductDefinitionRelationship_RelatedProductDefinition: ProductDefinition from StepBasic;
                       hasReferenceDesignator: Boolean;
                       aReferenceDesignator: HAsciiString from TCollection);
	---Purpose: Initialize all fields (own and inherited)

    ReferenceDesignator (me) returns HAsciiString from TCollection;
	---Purpose: Returns field ReferenceDesignator
    SetReferenceDesignator (me: mutable; ReferenceDesignator: HAsciiString from TCollection);
	---Purpose: Set field ReferenceDesignator
    HasReferenceDesignator (me) returns Boolean;
	---Purpose: Returns True if optional field ReferenceDesignator is defined

fields
    theReferenceDesignator: HAsciiString from TCollection; -- optional
    defReferenceDesignator: Boolean; -- flag "is ReferenceDesignator defined"

end AssemblyComponentUsage;
