-- Created on: 1993-01-26
-- Created by: Laurent PAINNOT
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package Approx 

     ---Purpose: Tis package provides algorithms approximating a set of
     --          points or curves with the possibility of dividing into
     --          one or many bezier curves.
     --          It also provides an instantiation for approximating
     --          a continous function f(t) into one or many curves. 
     
uses AdvApprox, 
     AppCont, 
     AppParCurves, 
     math, 
     gp,
     GeomAbs,
     Geom,
     Geom2d,
     Adaptor3d,
     Adaptor2d,
     TColStd, 
     TColGeom, 
     TColgp, 
     TCollection,  
     Standard, 
     StdFail


is

enumeration ParametrizationType is
    ChordLength,
    Centripetal,
    IsoParametric
end;    

enumeration Status is
    PointsAdded,
    NoPointsAdded,
    NoApproximation
end;
    
    
---------------------------------------------
---Algorithms for Bezier curves construction:
---------------------------------------------


   generic class ComputeLine, MyGradient;

   generic class ComputeCLine;

----------------------------------------------
---Algorithms for BSpline curves construction:
----------------------------------------------


    generic class BSplComputeLine, MyBSplGradient, MyGradientbis;

----------------------------------------------
---Algorithms for BSpline Surface construction:
----------------------------------------------
										   class  SweepApproximation; 
										   deferred  class  SweepFunction;
-----------------------------------------------------------------
--- Transformation of connecting MultiCurves into a MultiBSpCurve
-----------------------------------------------------------------


    class MCurvesToBSpCurve;

------------------------------------------------
---Algorithms  for  PCurve  approximation:
------------------------------------------------
    class  CurveOnSurface;  
    class  Curve3d;     
    class  Curve2d; 
------------------------------------------------
---Algorithms  for  PCurve  approximation:
------------------------------------------------
    class  CurvilinearParameter;  
    class  CurvlinFunc;
--------------------------
--- instantiate classes:
--------------------------

    imported SequenceOfHArray1OfReal;


-----------------------------------------------------------------
--- the folowing classes approximate a continous function f(t) in 
--- one or many bezier curves.
-----------------------------------------------------------------

    class FitAndDivide instantiates ComputeCLine from Approx
    	(Function from AppCont);

    class FitAndDivide2d instantiates ComputeCLine from Approx
    	(Function from AppCont);

    class SameParameter from Approx ;

    imported Array1OfAdHSurface;
    imported transient class HArray1OfAdHSurface;
    imported Array1OfGTrsf2d;
 
    imported transient class HArray1OfGTrsf2d; 
			    
    --    class ApproxPoints from Approx ;
    --    class ApproxPoints  from Approx ;
    --      this approximates a series of points
    --   Boundary conditions can be given as well
    --   a given parameterisation
    --   
 
end Approx;
