-- Created on: 1994-10-28
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class EdgeVertexInterference from TopOpeBRepDS 
    inherits ShapeShapeInterference from TopOpeBRepDS

    ---Purpose: An interference with a parameter.

uses

    Transition from TopOpeBRepDS,
    Config     from TopOpeBRepDS,
    Kind       from TopOpeBRepDS,    	
    OStream    from Standard    
    
is

    Create(T  : Transition from TopOpeBRepDS;
	   ST : Kind from TopOpeBRepDS;
	   S  : Integer from Standard;
	   G  : Integer from Standard;
      	   GIsBound : Boolean from Standard;
    	   C  : Config from TopOpeBRepDS;
	   P  : Real from Standard)
	   
    returns mutable EdgeVertexInterference from TopOpeBRepDS; 

    	---Purpose: Create an interference of VERTEX <G> on a crossed EDGE E.
    	--  
    	--  if support type <ST> == EDGE : <S> is edge E
    	--                          FACE : <S> is the face with bound E. 
    	--  <T> is the transition along the edge, crossing the crossed edge.
    	--   E  is the crossed edge.
    	--  <GIsBound> indicates if <G> is a bound of the edge.
    	--  <P> is the parameter of <G> on the edge.
    	--  
    	--  interference is stored in the list of interfs of the edge.
    	--  


    Create(T : Transition from TopOpeBRepDS;
	   S : Integer from Standard;
	   G : Integer from Standard;
      	   GIsBound : Boolean from Standard;
    	   C : Config from TopOpeBRepDS;
	   P : Real from Standard) 
	   
    	---Purpose: Create an interference of VERTEX <G> on crossed EDGE <S>.
    	--          
    	--  <T> is the transition along the edge, crossing the crossed edge.
    	--  <S> is the crossed edge.
    	--  <GIsBound> indicates if <G> is a bound of the edge.
    	--  <C> indicates the geometric configuration between
    	--        the edge and the crossed edge.
    	--  <P> is the parameter of <G> on the edge.
    	--  
    	--  interference is stored in the list of interfs of the edge.
    	--  

    returns mutable EdgeVertexInterference from TopOpeBRepDS; 
	    
    Parameter(me) returns Real from Standard
    is static;
    
    Parameter(me : mutable; P : Real from Standard)
    is static;

    Dump(me; OS : in out OStream from Standard) returns OStream
    is redefined;
    ---C++: return &
    
fields

    myParam : Real from Standard;

end EdgeVertexInterference from TopOpeBRepDS;
