-- Created by: DCB
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class PlotterParameter from PlotMgt inherits TShared from MMgt

uses
  FStream                 from Aspect,
  Plotter                 from PlotMgt,
  TypeOfPlotterParameter  from PlotMgt,
  HSequenceOfAsciiString  from TColStd,
  AsciiString             from TCollection,
  File                    from OSD

is
  -------------------------
  -- Category: Constructors
  -------------------------
  Create (
    aName  : AsciiString from TCollection
  ) returns mutable PlotterParameter from PlotMgt;
  ---Purpose: Create the class instance WITH undefined TYPE

  -----------------------------------------------
  -- Category: Methods to change class definition
  -----------------------------------------------
  Save (me: mutable; aFile: in out File from OSD)
  returns Boolean from Standard;
  ---Purpose:

  SetState (me: mutable; aState: Boolean from Standard);
  ---Purpose:

  SetType (me: mutable; aType: TypeOfPlotterParameter from PlotMgt);
  ---Purpose:

  ProcessParamVal (me: mutable;
    aParamSign :     CString from Standard;
    aFlag      :     Integer from Standard;
    aValue     : out AsciiString from TCollection
  ) is private;

  CheckListValue (me: mutable
  ) returns Boolean from Standard is private;
  ---Purpose:

  Normalize (me: mutable)
  is protected;
  ---Purpose:

  ----------------------------
  -- Category: Inquire methods
  ----------------------------
  SValue (me; aValue: out AsciiString from TCollection);
  ---Purpose:

  BValue (me)
  returns Boolean from Standard;
  ---Purpose:

  IValue (me)
  returns Integer from Standard;
  ---Purpose:

  RValue (me)
  returns Real from Standard;
  ---Purpose:

  LValues (me; aList: out HSequenceOfAsciiString from TColStd);
  ---Purpose:

  MValue (me
  ) returns HSequenceOfAsciiString from TColStd;
  ---Purpose:

  Name (me)
  returns AsciiString from TCollection;
  ---Purpose:

  OldName (me)
  returns AsciiString from TCollection;
  ---Purpose:

  Description (me : mutable)
  returns HSequenceOfAsciiString from TColStd
  is protected;
  ---Purpose:
  ---C++: return &

  NeedToBeSaved (me)
  returns Boolean from Standard;
  ---Purpose:

  Dump (me);
  ---Purpose:

  PutCommandInfo (me; outStream: FStream from Aspect);
  ---Purpose: Used to put parameter's information in a cmd file
  -- used in PlotterDriver's Spool method.

  ----------------------------------------
  -- Category: Methods to modify parameter
  ----------------------------------------
  SetSValue (me: mutable; aValue: AsciiString from TCollection);
  ---Purpose:

  SetBValue (me: mutable; aValue: Boolean from Standard);
  ---Purpose:

  SetIValue (me: mutable; aValue: Integer from Standard);
  ---Purpose:

  SetRValue (me: mutable; aValue: Real from Standard);
  ---Purpose:

  SetMValue (me: mutable; aMap: HSequenceOfAsciiString from TColStd);
  ---Purpose:

fields
  myName           : AsciiString            from TCollection;
  myOldName        : AsciiString            from TCollection;
  myType           : TypeOfPlotterParameter from PlotMgt;
  myIndex          : Integer                from Standard;
  myState          : Boolean                from Standard;
  myConfigState    : Boolean                from Standard;
  myIsModified     : Boolean                from Standard;
  --------------------------------------------------------
  myFlags          : Integer                from Standard;
  myDialog         : AsciiString            from TCollection;
  myMinValue       : AsciiString            from TCollection;
  myMaxValue       : AsciiString            from TCollection;
  myValues         : AsciiString            from TCollection;
  myDefValue       : AsciiString            from TCollection;
  myMapLength      : Integer                from Standard;
  myMap            : HSequenceOfAsciiString from TColStd;

  myDescription    : HSequenceOfAsciiString from TColStd;

friends
  class Plotter from PlotMgt

end PlotterParameter from PlotMgt;
