-- Created on: 1993-02-19
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



package BRepAdaptor 

	---Purpose: The BRepAdaptor package provides classes to access 
	--          the geometry of the BRep models.
	--          
	--          OverView of classes
	--          
	--          * Surface :  Provides the methods  of Surface from
	--          Adpator on a Face.
	--          
	--          *  Curve  : Provides  the  methods of  Curve  from
	--          Adaptor3d on an Edge.
	--          
	--          * Curve2d : Provides  the methods of  Curve2d from
	--          Adaptor2d on an Edge on a Face.
	--          

uses
    gp, 
    TCollection,
    TColgp,
    TColStd,
    GeomAbs,
    Adaptor3d,
    Adaptor2d,
    Geom,
    Geom2d,
    GeomAdaptor,
    Geom2dAdaptor,
    TopoDS,
    BRep

is

    class Surface;
	---Purpose: Transforms a Face in a Surface from Adaptor3d.
	
    class Curve;
	---Purpose: Transforms an Edge in a Curve from Adaptor3d.

    class Curve2d;
	---Purpose: Transforms an Edge   on a Face  in  a Curve2d from
	--          Adaptor2d. 

    class  CompCurve; 
    	---Purpose: Transforms a Wire in a Curve from Adaptor3d.
    	
    class HSurface instantiates GenHSurface from Adaptor3d
    	(Surface from BRepAdaptor);

    class HCurve instantiates GenHCurve from Adaptor3d
    	(Curve from BRepAdaptor);

    class HCurve2d instantiates GenHCurve2d from Adaptor2d
    	(Curve2d from BRepAdaptor); 
	 
    class HCompCurve instantiates GenHCurve from Adaptor3d
    	(CompCurve from BRepAdaptor); 
	 
    class Array1OfCurve 
    	instantiates Array1 from TCollection (Curve from BRepAdaptor); 
	 
    class HArray1OfCurve
    	instantiates HArray1 from TCollection (Curve from BRepAdaptor,
    	    	    	    	Array1OfCurve from BRepAdaptor);

end BRepAdaptor;
