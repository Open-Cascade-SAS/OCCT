-- Created on: 1992-08-21
-- Created by: Christophe MARION
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Intersection from HLRAlgo

	---Purpose: Describes  an intersection  on   an edge to  hide.
	--          Contains a parameter and   a state (ON =   on  the
	--          face, OUT = above the face, IN = under the Face)

uses
    Integer     from Standard,
    Real        from Standard,
    ShortReal   from Standard,
    Orientation from TopAbs,
    State       from TopAbs

is
    Create returns Intersection from HLRAlgo;

    Create(Ori    : Orientation from TopAbs;
           Lev    : Integer     from Standard;
           SegInd : Integer     from Standard;
           Ind    : Integer     from Standard;
           P      : Real        from Standard;
           Tol    : ShortReal   from Standard;
           S      : State       from TopAbs)
    returns Intersection from HLRAlgo;
    
    Orientation(me : in out; Ori : Orientation from TopAbs)
	---C++: inline
    is static;

    Orientation(me) returns Orientation from TopAbs
	---C++: inline
    is static;
    
    Level(me : in out; Lev : Integer from Standard)
	---C++: inline
    is static;

    Level(me) returns Integer from Standard
	---C++: inline
    is static;
    
    SegIndex(me : in out; SegInd : Integer from Standard)
	---C++: inline
    is static;

    SegIndex(me) returns Integer from Standard
	---C++: inline
    is static;
    
    Index(me : in out; Ind : Integer from Standard)
	---C++: inline
    is static;

    Index(me) returns Integer from Standard
	---C++: inline
    is static;
    
    Parameter(me : in out; P : Real from Standard)
	---C++: inline
    is static;

    Parameter(me) returns Real from Standard
	---C++: inline
    is static;
    
    Tolerance(me : in out; T : ShortReal from Standard)
	---C++: inline
    is static;
    
    Tolerance(me) returns ShortReal from Standard
	---C++: inline
    is static;
    
    State(me : in out; S : State from TopAbs)
	---C++: inline
    is static;

    State(me) returns State from TopAbs
	---C++: inline
    is static;

fields
    myOrien    : Orientation from TopAbs;
    mySegIndex : Integer     from Standard;
    myIndex    : Integer     from Standard;
    myLevel    : Integer     from Standard;
    myParam    : Real        from Standard;
    myToler    : ShortReal   from Standard;
    myState    : State       from TopAbs;

end Intersection;
