-- File:	StepFEA_SymmetricTensor43dMember.cdl
-- Created:	Tue Jan 14 10:53:27 2003
-- Author:	data exchange team
--		<det@petrox.nnov.matra-dtv.fr>
---Copyright:	 Matra Datavision 2003

class SymmetricTensor43dMember from StepFEA inherits SelectArrReal from StepData
    
    ---Purpose: Representation of member for  STEP SELECT type SymmetricTensor43d

is
    Create returns SymmetricTensor43dMember from StepFEA;
    ---Purpose: Empty constructor

    HasName (me) returns Boolean  is redefined;
    ---Purpose: Returns True if has name

    Name (me) returns CString  is redefined;
    ---Purpose: Returns set name

    SetName (me : mutable; name : CString)  returns Boolean  is redefined;
    ---Purpose: Set name

    Matches (me; name : CString) returns Boolean  is redefined;
    ---Purpose : Tells if the name of a SelectMember matches a given one;

fields

    mycase : Integer;                                                                                                         

end SymmetricTensor43dMember;
