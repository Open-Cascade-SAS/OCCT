-- Created on: 1997-01-22
-- Created by: Prestataire Michael ALEONARD
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SymmetricPresentation from DsgPrs
    	---Purpose: A framework to define display of symmetry between shapes.
uses
    Presentation from Prs3d,
    Pnt  from gp,
    Dir  from gp,
    Lin  from gp,
    Circ from gp,
    Drawer from Prs3d,
    ExtendedString from TCollection
    	
is  
    Add( myclass; aPresentation: Presentation from Prs3d;
    	    	  aDrawer: Drawer from Prs3d;
	       	  AttachmentPoint1: Pnt from gp;
		  AttachmentPoint2: Pnt from gp;
		  aDirection1: Dir from gp;  
		  aAxis: Lin from gp;
		  OffsetPoint: Pnt from gp);
	---Purpose: Adds the points OffsetPoint, AttachmentPoint1,
    	-- AttachmentPoint2, the direction aDirection1 and the
    	-- axis anAxis to the presentation object aPresentation.
    	-- The display attributes of the symmetry are defined by
    	-- the attribute manager aDrawer.
    	-- This syntax is used for display of symmetries between two segments.
		  
     
    Add( myclass; aPresentation: Presentation from Prs3d;
    	    	  aDrawer: Drawer from Prs3d;
	       	  AttachmentPoint1: Pnt from gp;
		  AttachmentPoint2: Pnt from gp; 
		  aCircle1: Circ from gp;
		  aAxis: Lin from gp;
		  OffsetPoint: Pnt from gp);
	---Purpose: Adds the points OffsetPoint, AttachmentPoint1,
    	-- AttachmentPoint2, the direction aDirection1 the circle
    	-- aCircle1 and the axis anAxis to the presentation
    	-- object aPresentation.
    	-- The display attributes of the symmetry are defined by
    	-- the attribute manager aDrawer.
    	-- This syntax is used for display of symmetries between two arcs.
	  
    Add( myclass; aPresentation: Presentation from Prs3d;
    	    	  aDrawer: Drawer from Prs3d;
	       	  AttachmentPoint1: Pnt from gp;
		  AttachmentPoint2: Pnt from gp; 
	          aAxis: Lin from gp;
	          OffsetPoint: Pnt from gp);
	---Purpose: Adds the points OffsetPoint, AttachmentPoint1,
    	-- AttachmentPoint2 and the axis anAxis to the
    	-- presentation object aPresentation.
    	-- The display attributes of the symmetry are defined by
    	-- the attribute manager aDrawer.
    	-- This syntax is used for display of symmetries between two vertices.
		  
end SymmetricPresentation;









