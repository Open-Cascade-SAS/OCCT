-- Created on: 1997-07-28
-- Created by: Pierre CHALAMET
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Texture1Dsegment from Graphic3d

inherits Texture1D from Graphic3d

  ---Purpose:  This class provides the implementation
  -- of a 1D texture applyable along a segment.
  -- You might use the SetSegment() method
  -- to set the way the texture is "streched" on facets.

uses

  NameOfTexture1D from Graphic3d,
  AsciiString     from TCollection

is

  Create (theFileName : AsciiString from TCollection) returns mutable Texture1Dsegment from Graphic3d;
  ---Purpose: Creates a texture from a file

  Create (theNOT : NameOfTexture1D from Graphic3d) returns mutable Texture1Dsegment from Graphic3d;
  ---Purpose: Creates a texture from a predefined texture name set.

  SetSegment (me : mutable;
              theX1, theY1, theZ1 : ShortReal from Standard;
              theX2, theY2, theZ2 : ShortReal from Standard);
  ---Purpose: Sets the texture application bounds. Defines the way
  -- the texture is stretched across facets.
  -- Default values are <0.0, 0.0, 0.0> , <0.0, 0.0, 1.0>

  --
  -- inquire methods
  --
  Segment (me;
           theX1, theY1, theZ1 : out ShortReal from Standard;
           theX2, theY2, theZ2 : out ShortReal from Standard);
  ---Purpose: Returns the values of the current segment X1, Y1, Z1 , X2, Y2, Z2.

fields

  myX1, myY1, myZ1 : ShortReal from Standard;
  myX2, myY2, myZ2 : ShortReal from Standard;
      
end  Texture1Dsegment;
