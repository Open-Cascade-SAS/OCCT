-- Created on: 1992-05-05
-- Created by: Remi GILET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package GCE2d

uses gp,
     Geom2d,
     gce,
     StdFail


    ---Level : Public. 
    --  All methods of all  classes will be public.



is

private deferred class Root;

---------------------------------------------------------------------------
--          Constructions of 2d geometrical elements from Geom2d.
---------------------------------------------------------------------------

class MakeLine;
    	---Purpose: Makes a Line from Geom2d.

class MakeCircle;
    	---Purpose: Makes a Circle from Geom2d.

class MakeHyperbola;
    	---Purpose: Makes an hyperbola from Geom2d.

class MakeEllipse;
    	---Purpose: Makes an Ellipse from Geom2d.

class MakeParabola;
    	---Purpose: Makes a parabola from Geom2d.

class MakeSegment;
    	---Purpose: Makes a segment of Line (TrimmedCurve from Geom2d).

class MakeArcOfCircle;
    	---Purpose: Makes an arc of circle (TrimmedCurve from Geom2d).

class MakeArcOfEllipse;
    	---Purpose: Makes an arc of ellipse (TrimmedCurve from Geom2d).

class MakeArcOfParabola;
    	---Purpose: Makes an arc of parabola (TrimmedCurve from Geom2d).

class MakeArcOfHyperbola;
    	---Purpose: Makes an arc of hyperbola (TrimmedCurve from Geom2d).

---------------------------------------------------------------------------
--              Constructions of Transformation from Geom2d.
---------------------------------------------------------------------------

class MakeTranslation;
    	---Purpose: Returns a translation transformation.
 
class MakeMirror;
    	---Purpose: Returns a symmetry transformation. 

class MakeRotation;
    	---Purpose: Returns a rotation transformation.

class MakeScale;
    	---Purpose: Returns a scaling transformation.

    
end GCE2d;



