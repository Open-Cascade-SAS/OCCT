-- Created on: 1992-08-13
-- Created by: Remi LEQUETTE
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package TopBas 

	---Purpose: The  TopBas package  provides  data structure  for
	--          topological algorithms.   THe data  structures are
	--          used to store the intermediary dat and the results
	--          of the algorithms.
	--          
	--          *  Interference, List  :  An Interference  is  the
	--          topological    representation  of an intersection.
	--          The classes are generic in order to be independant
	--          of the data structure.

uses
    Standard,
    TCollection,
    TopAbs

is
    generic class Interference;
	---Purpose: The   Interference  is  the    description  of  an
	--          intersection on a Shape.

    class TestInterference instantiates Interference from TopBas
    	    	    	    (Real    from Standard,
    	    	    	     Integer from Standard);
			    
    class ListOfTestInterference instantiates 
    List from TCollection (TestInterference);

end TopBas;


