-- File:        RatioMeasureWithUnit.cdl
-- Created:     Mon Dec  4 12:02:30 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWRatioMeasureWithUnit from RWStepBasic

	---Purpose : Read & Write Module for RatioMeasureWithUnit

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     RatioMeasureWithUnit from StepBasic,
     EntityIterator from Interface

is

	Create returns RWRatioMeasureWithUnit;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable RatioMeasureWithUnit from StepBasic);

	WriteStep (me; SW : in out StepWriter; ent : RatioMeasureWithUnit from StepBasic);

	Share(me; ent : RatioMeasureWithUnit from StepBasic; iter : in out EntityIterator);

end RWRatioMeasureWithUnit;
