-- Created on: 2002-12-15
-- Created by: data exchange team
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class StructuralResponsePropertyDefinitionRepresentation from StepRepr
inherits PropertyDefinitionRepresentation from StepRepr

    ---Purpose: Representation of STEP entity StructuralResponsePropertyDefinitionRepresentation

uses
    PropertyDefinition from StepRepr,
    Representation from StepRepr

is
    Create returns StructuralResponsePropertyDefinitionRepresentation from StepRepr;
	---Purpose: Empty constructor

end StructuralResponsePropertyDefinitionRepresentation;
