-- Created on: 1995-12-04
-- Created by: Stephane MORTAUD
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

--last modifs by rob 29-01-96 : heritage de CompositionFilter


class OrFilter from SelectMgr inherits CompositionFilter from SelectMgr

    	---Purpose: A framework to define an or selection filter.
    	-- This selects one or another type of sensitive entity.
uses

    Filter       from SelectMgr,
    Transient    from Standard,
    EntityOwner  from SelectMgr

is

    Create
    returns mutable OrFilter from SelectMgr;
    	---Purpose: Constructs an empty or selection filter.
    IsOk(me; anobj : EntityOwner from SelectMgr)
    returns Boolean from Standard ;

end OrFilter;
