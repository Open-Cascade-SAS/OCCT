-- Created on: 1993-01-09
-- Created by: CKY / Contract Toubro-Larsen (Kiran)
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class CompositeCurve from IGESGeom  inherits IGESEntity

        ---Purpose: defines IGESCompositeCurve, Type <102> Form <0>
        --          in package IGESGeom
        --          A composite curve is defined as an ordered list of entities
        --          consisting of a point, connect point and parametrised curve
        --          entities (excluding the CompositeCurve entity).

uses

        HArray1OfIGESEntity from IGESData

raises OutOfRange

is

        Create returns mutable CompositeCurve;

        -- Specific Methods pertaining to the class

        Init (me          : mutable;
              allEntities : HArray1OfIGESEntity);
         ---Purpose : This method is used to set the fields of the class
         --           CompositeCurve
         --       - allEntities : Constituent Entities of the composite curve

        NbCurves (me) returns Integer;
        ---Purpose : returns the number of curves contained in the CompositeCurve

        Curve (me; Index : Integer) returns IGESEntity
        raises OutOfRange;
        ---Purpose : returns Component of the CompositeCurve (a curve or a point)
        -- raises exception if Index <= 0 or Index > NbCurves()

fields

--
-- Class    : IGESGeom_CompositeCurve
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class CompositeCurve.
--
-- Reminder : A CompositeCurve instance is defined by :
--            The collection of constituent curves which could
--            be of type point, connect point or parametric curve
--            entities

        theEntities : HArray1OfIGESEntity;

end CompositeCurve;
