-- Created on: 1997-09-18
-- Created by: Christophe MARION
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class BiPoint from BRepMesh

uses
    Address from Standard,
    Real    from Standard,
    Integer from Standard
    
is
    Create
    returns BiPoint from BRepMesh; 
    	---C++: inline
    
    Create(X1,Y1,X2,Y2 : Real    from Standard)
    returns BiPoint from BRepMesh; 
    
    Indices(me) returns Address from Standard
    	---C++: inline
    is static;

    Coordinates(me) returns Address from Standard
    	---C++: inline
    is static;

fields
    myIndices     : Integer from Standard[2];
    myCoordinates : Real    from Standard[6];
    
end BiPoint;
