-- Created on: 1991-07-17
-- Created by: Isabelle GRIGNON
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class FunctionSample from math 

	---Purpose: This class gives a default sample (constant difference
	--          of parameter) for a function defined between
	--          two bound A,B.

raises OutOfRange from Standard

is

    Create(A,B: Real; N: Integer)
    
    	returns FunctionSample from math;


    Bounds(me; A,B: out Real) is virtual;
    
	---Purpose: Returns the bounds of parameters.



    NbPoints(me)
    
	---Purpose: Returns the number of sample points.

    returns Integer
    is static;


    GetParameter(me; Index: Integer)
    
	---Purpose: Returns the value of parameter of the point of 
	--          range Index : A + ((Index-1)/(NbPoints-1))*B.
	--          An exception is raised if Index<=0 or Index>NbPoints.

    returns Real
    raises OutOfRange
    is virtual;



fields

    a: Real;
    b: Real;
    n: Integer;

end FunctionSample;
