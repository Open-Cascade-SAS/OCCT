-- Created on: 1993-11-10
-- Created by: Jean Marc LACHAUME
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Hatching from Geom2dHatch

uses
    ErrorStatus      from HatchGen ,
    PointOnHatching  from HatchGen ,
    PointsOnHatching from HatchGen ,
    Domain           from HatchGen ,
    Domains          from HatchGen , 
    Pnt2d            from gp,
    Curve            from Geom2dAdaptor

raises
    OutOfRange   from Standard

is

     Create
       
       returns Hatching from Geom2dHatch;


    Create (Curve : Curve from Geom2dAdaptor)
    
    	---Purpose: Creates a hatching.

	returns Hatching from Geom2dHatch ;


    Curve (me)
    
    	---Purpose: Returns the curve associated to the hatching.

    	---C++: return const &

        returns Curve from Geom2dAdaptor
        is static ;


    ChangeCurve (me : in out)
    
    	---Purpose: Returns the curve associated to the hatching.

    	---C++: return &

        returns Curve from Geom2dAdaptor
        is static ;


    TrimDone (me : in out ; Flag : Boolean from Standard)

    	---Purpose: Sets the flag about the trimming computations to the
    	--          given value.

    	is static ;


    TrimDone (me)

    	---Purpose: Returns the flag about the trimming computations.

    	returns Boolean from Standard
	is static ;


    TrimFailed (me : in out ; Flag : Boolean from Standard)

    	---Purpose: Sets the flag about the trimming failure to the
    	--          given value.

    	is static ;


    TrimFailed (me)

    	---Purpose: Returns the flag about the trimming failure.

    	returns Boolean from Standard
	is static ;


    IsDone (me : in out ; Flag : Boolean from Standard)

    	---Purpose: Sets the flag about the domains computation to the
    	--          given value.

    	is static ;


    IsDone (me)

    	---Purpose: Returns the flag about the domains computation.

    	returns Boolean from Standard
	is static ;


    Status (me : in out ; Status : ErrorStatus from HatchGen)

    	---Purpose: Sets the error status.

    	is static ;


    Status (me)

    	---Purpose: Returns the error status.

    	returns ErrorStatus from HatchGen
	is static ;


---Category: Points on hatching.

    AddPoint (me : in out ; Point     : PointOnHatching from HatchGen ;
    	    	    	    Confusion : Real            from Standard)
    
    	---Purpose: Adds an intersection point to the hatching.

	is static ;


    NbPoints (me)
    
    	---Purpose: Returns the number of intersection points
    	--          of the hatching.

        returns Integer from Standard
        is static ;


    Point (me ; Index : Integer from Standard)
    
    	---Purpose: Returns the Index-th intersection point of the
    	--          hatching.
    	--          The exception OutOfRange is raised if
    	--          Index < 1 or Index > NbPoints.

    	---C++: return const &

    	returns PointOnHatching from HatchGen
    	raises OutOfRange from Standard
   	is static ;


    ChangePoint (me : in out ; Index : Integer from Standard)
    
    	---Purpose: Returns the Index-th intersection point of the
    	--          hatching.
    	--          The exception OutOfRange is raised if
    	--          Index < 1 or Index > NbPoints.

    	---C++: return &

    	returns PointOnHatching from HatchGen
    	raises OutOfRange from Standard
   	is static ;


    RemPoint (me : in out ; Index : Integer from Standard)
    
    	---Purpose: Removes the Index-th intersection point of the
    	--          hatching.
    	--          The exception OutOfRange is raised if
    	--          Index < 1 or Index > NbPoints.

    	raises OutOfRange from Standard
    	is static ;


    ClrPoints (me : in out)
    
    	---Purpose: Removes all the intersection points of the hatching.

    	is static ;


---Category: Domains.


    AddDomain (me : in out ; Domain : Domain from HatchGen)
    
    	---Purpose: Adds a domain to the hatching.

	is static ;


    NbDomains (me)
    
    	---Purpose: Returns the number of domains of the hatching.

        returns Integer from Standard
        is static ;


    Domain (me ; Index : Integer from Standard)
    
    	---Purpose: Returns the Index-th domain of the hatching.
    	--          The exception OutOfRange is raised if
    	--          Index < 1 or Index > NbDomains.

    	---C++: return const &

    	returns Domain from HatchGen
    	raises OutOfRange from Standard
   	is static ;


    RemDomain (me : in out ; Index : Integer from Standard)
    
    	---Purpose: Removes the Index-th domain of the hatching.
    	--          The exception OutOfRange is raised if
    	--          Index < 1 or Index > NbDomains.

    	raises OutOfRange from Standard
    	is static ;


    ClrDomains (me : in out)
    
    	---Purpose: Removes all the domains of the hatching.

    	is static ;


    ClassificationPoint (me) 
    	---Purpose: Returns a point on the curve. 
    	--          This point will be used for the classification.
    returns Pnt2d from gp
    is static;
       
fields

    myCurve      : Curve from Geom2dAdaptor ;
    myTrimDone   : Boolean          from Standard ;
    myTrimFailed : Boolean          from Standard ;
    myPoints     : PointsOnHatching from HatchGen ;
    myIsDone     : Boolean          from Standard ;
    myStatus     : ErrorStatus      from HatchGen ;
    myDomains    : Domains          from HatchGen ;

end Hatching from Geom2dHatch ;
