-- Created by: DAUTRY Philippe
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

--      	---------------------------

---Version:	0.0
--Version	Date		Purpose
--		0.0	Sep 17 1997	Creation


class XLinkStorageDriver from MDocStd
    inherits ASDriver from MDF

	---Purpose: Tool used to translate a transient XLink into a
	--          persistent one.

uses

    SRelocationTable from MDF,
    Attribute        from TDF,
    Attribute        from PDF, 
    MessageDriver    from CDM

is

    Create(theMessageDriver : MessageDriver from CDM) -- Version 0
    returns XLinkStorageDriver from MDocStd;

    VersionNumber(me) returns Integer from Standard;
	---Purpose: Returns the version number from which the driver
	--          is available: 0.

    SourceType(me) returns Type from Standard;
	---Purpose: Returns the type: XLink from TXLink.

    NewEmpty (me)
    returns Attribute from PDF;


    Paste(me;
    	  aSource     :         Attribute        from TDF;
    	  aTarget     : Attribute        from PDF;
    	  aRelocTable :         SRelocationTable from MDF);
	  
	  
end XLinkStorageDriver;
