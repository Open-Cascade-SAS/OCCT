-- Created on: 1995-10-24
-- Created by: Mister rmi
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PolygonOnClosedSurface from PBRep

    inherits PolygonOnSurface from PBRep
    
    	---Purpose: Representation by two 2d polygons in the parametric
	--          space of a surface.

uses Polygon2D           from PPoly,
     Surface             from PGeom,
     Location            from PTopLoc



is
    Create(P1: Polygon2D from PPoly;
    	   P2: Polygon2D from PPoly;
    	   S:  Surface   from PGeom;
	   L:  Location  from PTopLoc)
    returns mutable PolygonOnClosedSurface from PBRep;
    
    IsPolygonOnClosedSurface(me) returns Boolean
    	---Purpose: returns True.
    is redefined;

    Polygon2(me) returns any Polygon2D from PPoly;

    
fields

    myPolygon2: Polygon2D from PPoly;

end PolygonOnClosedSurface;
