-- Created on: 1993-07-05
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Update:      Frederic MAUPAS



deferred class CurveRepresentation from PBRep inherits Persistent

	---Purpose: Root class for the curve representations.

uses
    Location from PTopLoc


is

    Initialize(L : Location from PTopLoc);
    	---Level: Internal 

    Location(me) returns Location from PTopLoc
    is static;
    	---Level: Internal 
    
    Next(me) returns CurveRepresentation from PBRep
    is static;
    	---Level: Internal 
		
    Next(me : mutable; N :  CurveRepresentation from PBRep)
    is static;
    	---Level: Internal 

    ------------------------------------------------------
    -- What kind of representation : used to speed Mapping
    ------------------------------------------------------

    IsCurve3D(me)               returns Boolean
	 ---Purpose: A 3D curve representation.
    is virtual;

    IsCurveOnSurface(me)        returns Boolean
	---Purpose: A curve in the parametric space of a surface.
    is virtual;

    IsRegularity(me)            returns Boolean
	---Purpose: A continuity between two surfaces.
    is virtual;
    
    IsCurveOnClosedSurface(me)  returns Boolean
	---Purpose: A curve with two parametric   curves  on the  same
	--          surface. 
    is virtual;

    IsGCurve(me) returns Boolean from Standard
    	---Purpose:
    is virtual;
    
    IsPolygon3D(me) returns Boolean
	---Purpose: 
    is virtual;
    
    IsPolygonOnTriangulation(me) returns Boolean
	---Purpose: 
    is virtual;

    IsPolygonOnClosedTriangulation(me) returns Boolean
	---Purpose: 
    is virtual;

    IsPolygonOnSurface(me) returns Boolean
	---Purpose: 
    is virtual;

    IsPolygonOnClosedSurface(me) returns Boolean
	---Purpose: 
    is virtual;
    
    
fields
    
    myLocation : Location from PTopLoc;
    myNext     : CurveRepresentation from PBRep;

end CurveRepresentation;
