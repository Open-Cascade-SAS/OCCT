-- Created on: 1996-04-01
-- Created by: Philippe MANGIN
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

private class EnergyOfMVC from FairCurve  inherits Energy from FairCurve

	---Purpose: Energy Criterium to minimize in MinimalVariationCurve.
	---Category: Private use

uses BattenLaw from FairCurve,  
     DistributionOfTension from FairCurve, 
     DistributionOfSagging from FairCurve,
     DistributionOfJerk    from FairCurve,
     AnalysisCode from FairCurve,
     Vector  from  math,
     Matrix  from math,
     HArray1OfPnt2d from TColgp,
     Array1OfXY  from TColgp,
     Pnt2d from gp,
     HArray1OfReal from TColStd
     
raises DomainError


is
    Create( BSplOrder     : Integer;
            FlatKnots     : HArray1OfReal;
	    Poles         : HArray1OfPnt2d;
    	    ContrOrder1   : Integer;
	    ContrOrder2   : Integer;
	    Law           : BattenLaw;
	    PhysicalRatio : Real;
	    LengthSliding : Real;
	    FreeSliding   : Boolean = Standard_True;
            Angle1        : Real = 0;
            Angle2        : Real = 0;
    	    Curvature1    : Real = 0;
    	    Curvature2    : Real = 0 )
     ---Purpose: Angles corresspond to the Ox axis
     returns  EnergyOfMVC
     raises  DomainError; -- if  PhysicalRatio < 0 or  PhysicalRatio > 1
    
    LengthSliding(me)
    ---Purpose: return  the  lengthSliding = P1P2 + Sliding
    ---C++: inline
    returns  Real;
    
         
    Status(me) 
    ---Purpose: return  the status 
    ---C++: inline
    returns  AnalysisCode;
    
    ComputePoles(me: in out; X: Vector)
    ---Purpose: compute  the  poles wich correspond with the variable X
    is redefined protected; 
    
    Variable(me; X: out Vector)
    ---Purpose: compute the variables <X> wich correspond with the field <MyPoles>
    returns Boolean
    is redefined;  
	
    Compute(me:in out; DerivativeOrder : Integer; Result : out Vector)
        ---Purpose: compute the energy in intermediat format
    returns Boolean 
    is redefined protected;
    
fields
    MyLengthSliding : Real;
    OriginalSliding : Real;
    MyBattenLaw     : BattenLaw;
    MyPhysicalRatio : Real;
    MyTension       : DistributionOfTension;
    MySagging       : DistributionOfSagging;
    MyJerk          : DistributionOfJerk;
    MyStatus        : AnalysisCode;

end EnergyOfMVC;
