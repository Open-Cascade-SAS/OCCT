-- Created on: 1994-09-02
-- Created by: Yves FRICAUD
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

private generic class FuncCurNul from LProp (Curve as any;
                                             Vec   as any; -- as Vec or Vec2d
		     	                     Pnt   as any; -- as Pnt or Pnt2d
		   	                     Dir   as any; -- as Dir or Dir2d Vec  
    	    	    	    	    	     Tool  as any) -- as Tool(Curve, Pnt, Vec)
inherits FunctionWithDerivative from math
	---Purpose: Function used to find the inflections in 2d. 

is
    Create ( C : Curve) returns FuncCurNul from LProp;
    
    Value (me : in out; X : Real; F : out Real)
    	---Purpose: Returns the value for the variable <X>.
    returns Boolean;
    
    Derivative(me : in out; X : Real; D : out Real)
        ---Purpose: Returns the derivative for the variable <X>
    returns Boolean;

    Values(me : in out ; X  : Real; F  : out Real; D  : out Real)    
    	---Purpose: Returns the value of the function and the derivative
    	--          for the variable <X>.
    returns Boolean;    

fields
    theCurve : Curve;
    
end FuncCurNul;

