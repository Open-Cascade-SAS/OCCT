-- Created on: 1992-09-28
-- Created by: Remi GILET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MakeArcOfHyperbola from GCE2d inherits Root from GCE2d
    	---Purpose: Implements construction algorithms for an arc of
    	-- hyperbola in the plane. The result is a Geom2d_TrimmedCurve curve.
    	-- A MakeArcOfHyperbola object provides a framework for:
    	-- -   defining the construction of the arc of hyperbola,
    	-- -   implementing the construction algorithm, and
    	-- -   consulting the results. In particular, the Value
    	--   function returns the constructed arc of hyperbola.
  
uses Pnt2d        from gp,
     Hypr2d       from gp,
     Real         from Standard,
     Boolean      from Standard,
     TrimmedCurve from Geom2d

raises NotDone from StdFail

is

Create(Hypr           : Hypr2d  from gp                      ;
       Alpha1, Alpha2 : Real    from Standard                ;
       Sense          : Boolean from Standard = Standard_True) 
    returns MakeArcOfHyperbola;
    	---Purpose: Makes an arc of Hyperbola (TrimmedCurve from Geom2d) from 
    	--          a Hyperbola between two parameters Alpha1 and Alpha2.

Create(Hypr  : Hypr2d  from gp                      ;
       P     : Pnt2d   from gp                      ;
       Alpha : Real    from Standard                ;
       Sense : Boolean from Standard = Standard_True) 
    returns MakeArcOfHyperbola;
    	---Purpose: Makes an arc of Hyperbola (TrimmedCurve from Geom2d) from 
    	--          a Hyperbola between point <P> and the parameter
        --          Alpha.

Create(Hypr  : Hypr2d  from gp                      ;
       P1    : Pnt2d   from gp                      ;
       P2    : Pnt2d   from gp                      ;
       Sense : Boolean from Standard = Standard_True) 
    returns MakeArcOfHyperbola;
    	---Purpose: Makes an arc of Hyperbola (TrimmedCurve from Geom2d) from 
    	--          a Hyperbola between two points P1 and P2.
    	-- Note: the orientation of the arc of hyperbola is:
    	-- -   the trigonometric sense if Sense is not defined or
    	--   is true (default value), or
    	-- -   the opposite sense if Sense is false.
    	-- - IsDone always returns true.
        
Value(me) returns TrimmedCurve from Geom2d
    raises NotDone
    is static;
    	---C++: return const&
    	---Purpose: Returns the constructed arc of hyperbola.
        ---C++: alias "operator const Handle(Geom2d_TrimmedCurve)& () const { return Value(); }"

fields

    TheArc : TrimmedCurve from Geom2d;
    --The solution from Geom2d.
    
end MakeArcOfHyperbola;
