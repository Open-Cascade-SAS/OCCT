-- Created on: 1998-06-03
-- Created by: data exchange team
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- szv#4 S4163

class WireVertex from ShapeAnalysis 

	---Purpose: Analyzes and records status of vertices in a Wire
    	--           
    	--          The Wire has formerly been loaded in a ShapeExtend_WireData
    	--          For each Vertex, a status and some data can be attached
    	--          (case found, position and parameters)
    	--          Then, these informations can be used to fix problems

uses
    XYZ              from gp,
    HArray1OfXYZ     from TColgp,
    HArray1OfInteger from TColStd,
    HArray1OfReal    from TColStd,
    Wire             from TopoDS,
    WireData         from ShapeExtend

is
    Create returns WireVertex;
    	---Purpose: Empty constructor
	
    Init (me: in out; wire: Wire from TopoDS; preci : Real);

    Init (me: in out; swbd: WireData from ShapeExtend; preci : Real);

    Load (me: in out; wire: Wire from TopoDS);
    	
    Load (me: in out; sbwd: WireData from ShapeExtend);

    SetPrecision (me: in out; preci: Real);
    	---Purpose: Sets the precision for work
    	--          Analysing: for each Vertex, comparison between the end of the
    	--          preceeding edge and the start of the following edge
    	--          Each Vertex rank corresponds to the End Vertex of the Edge of
    	--          same rank, in the ShapeExtend_WireData. I.E. for Vertex <num>,
    	--          Edge <num> is the preceeding one, <num+1> is the following one

    Analyze (me: in out);

    SetSameVertex (me: in out; num: Integer);
    	---Purpose: Records status "Same Vertex" (logically) on Vertex <num>

    SetSameCoords (me: in out; num: Integer);
    	---Purpose: Records status "Same Coords" (at the Vertices Tolerances)

    SetClose (me: in out; num: Integer);
    	---Purpose: Records status "Close Coords" (at the Precision of <me>)

    SetEnd (me: in out; num : Integer;
    	    	        pos : XYZ from gp;
    	    	    	ufol: Real);
    	---Purpose: <num> is the End of preceeding Edge, and its projection on the
    	--          following one lies on it at the Precision of <me>
    	--          <ufol> gives the parameter on the following edge

    SetStart (me: in out; num : Integer;
    	    	          pos : XYZ from gp;
    	    	    	  upre: Real);
    	---Purpose: <num> is the Start of following Edge, its projection on the
    	--          preceeding one lies on it at the Precision of <me>
    	--          <upre> gives the parameter on the preceeding edge

    SetInters (me: in out; num      : Integer;
    	    	    	   pos      : XYZ from gp;
    	    	    	   upre,ufol: Real);
    	---Purpose: <num> is the Intersection of both Edges
    	--          <upre> is the parameter on preceeding edge, <ufol> on
    	--          following edge

    SetDisjoined (me: in out; num: Integer);
    	---Purpose: <num> cannot be said as same vertex


    IsDone (me) returns Boolean;
    	---Purpose: Returns True if analysis was performed, else returns False
	
    Precision (me) returns Real;
    	---Purpose: Returns precision value used in analysis
    
    NbEdges (me) returns Integer;
    	---Purpose: Returns the number of edges in analyzed wire (i.e. the
	--          length of all arrays)
    
    WireData (me) returns WireData from ShapeExtend;
    	---Purpose: Returns analyzed wire
    	---C++ : return const &
	
    Status (me; num: Integer) returns Integer;
    	---Purpose: Returns the recorded status for a vertex
    	--          More detail by method Data
	
    Position (me; num: Integer) returns XYZ from gp;
    
    UPrevious(me; num: Integer) returns Real; --szv#4:S4163:12Mar99 was Interger
    
    UFollowing(me; num: Integer) returns Real; --szv#4:S4163:12Mar99 was Interger
    
    Data(me; num      : Integer;
    	     pos      : out XYZ from gp;
    	     upre,ufol: out Real)
    returns Integer;
    	---Purpose: Returns the recorded status for a vertex
    	--          With its recorded position and parameters on both edges
    	--          These values are relevant regarding the status:
    	--          Status  Meaning   Position  Preceeding  Following
    	--          0       Same       no        no          no
    	--          1       SameCoord  no        no          no
    	--          2       Close      no        no          no
    	--          3       End        yes       no          yes
    	--          4       Start      yes       yes         no
    	--          5       Inters     yes       yes         yes
    	--         -1       Disjoined  no        no          no

    NextStatus (me; stat: Integer; num : Integer = 0) returns Integer;
    	---Purpose: For a given status, returns the rank of the vertex which
    	--          follows <num> and has the same status. 0 if no more
    	--          Acts as an iterator, starts on the first one

    NextCriter(me; crit: Integer; num : Integer = 0) returns Integer;
    	---Purpose: For a given criter, returns the rank of the vertex which
    	--           follows <num> and has the same status. 0 if no more
    	--           Acts as an iterator, starts on the first one
    	--           Criters are:
    	--           0: same vertex (status 0)
    	--           1: a solution exists (status >= 0)
    	--           2: same coords (i.e. same params) (status 0 1 2)
    	--           3: same coods but not same vertex (status 1 2)
    	--           4: redefined coords (status 3 4 5)
    	--          -1: no solution (status -1)

fields

    myWire: WireData from ShapeExtend;
    myStat: HArray1OfInteger from TColStd;
    myPos : HArray1OfXYZ from TColgp;
    myUPre: HArray1OfReal from TColStd;
    myUFol: HArray1OfReal from TColStd;
    myPreci: Real;
    myDone: Boolean;

end WireVertex;
