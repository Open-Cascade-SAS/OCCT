-- File:	PTColStd.cdl
-- Created:	Fri Jul  5 15:49:10 1996
-- Author:	Jean-Louis Frenkel
--		<rmi@pernox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1996


package PTColStd

uses
    Standard,TColStd,TCollection
   ---Category:  reusable class
   --           
is

   class MapPersistentHasher instantiates MapHasher from TCollection(Persistent);

   class DoubleMapOfTransientPersistent  instantiates   
	     DoubleMap from TCollection(Transient from Standard,
      	    	    	    	 Persistent from Standard,
      	    	    	    	 MapTransientHasher from TColStd,
    	    	    	    	 MapPersistentHasher from PTColStd);  

   class TransientPersistentMap instantiates 
   DataMap from TCollection(Transient from Standard,
                            Persistent from Standard,
	       	            MapTransientHasher from TColStd);
    
   class PersistentTransientMap instantiates
   DataMap from TCollection(Persistent from Standard,
                             Transient from Standard,
                             MapPersistentHasher from PTColStd);

end PTColStd;
