-- Created on: 1999-04-30
-- Created by: data exchange team
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ShapeDivideContinuity from ShapeUpgrade inherits ShapeDivide from ShapeUpgrade

	---Purpose: API Tool for converting shapes with C0 geometry into C1 ones

uses
    
    Shape from TopoDS,
    Shape from GeomAbs,
    FaceDivide from ShapeUpgrade

is
    Create returns ShapeDivideContinuity from ShapeUpgrade;
    
    Create (S: Shape from TopoDS)
    returns ShapeDivideContinuity from ShapeUpgrade;
    	---Purpose: Initialize by a Shape.
    
    SetTolerance(me: in out; Tol: Real);
    	---Purpose: Sets tolerance.
    
    SetTolerance2d(me: in out; Tol: Real);
    	---Purpose: Sets tolerance.
    
    SetBoundaryCriterion (me: in out; Criterion: Shape from GeomAbs = GeomAbs_C1);
    	---Purpose: 
        --  Defines a criterion of continuity for the boundary (all the
        --  Wires)
        --  
        --  The possible values are C0, G1, C1, G2, C2, C3, CN The
        --  default is C1 to respect the Cas.Cade Shape Validity.  G1
        --  and G2 are not authorized.
	
    SetPCurveCriterion (me: in out; Criterion: Shape from GeomAbs = GeomAbs_C1);
    	---Purpose: 
        --  Defines a criterion of continuity for the boundary (all the
        --  pcurves of Wires)
        --  
        --  The possible values are C0, G1, C1, G2, C2, C3, CN The
        --  default is C1 to respect the Cas.Cade Shape Validity.  G1
        --  and G2 are not authorized.
    
    SetSurfaceCriterion (me: in out; Criterion: Shape from GeomAbs = GeomAbs_C1);
    	---Purpose: 
        --  Defines a criterion of continuity for the boundary (all the
        --  Wires)
        --  
        --  The possible values are C0, G1, C1, G2, C2, C3, CN The
        --  default is C1 to respect the Cas.Cade Shape Validity.  G1
        --  and G2 are not authorized.
    
    ---Level: Internal
    
    GetSplitFaceTool (me) returns FaceDivide from ShapeUpgrade
    is redefined protected;
    	---Purpose: Returns the tool for dividing faces.
    
fields

    myCurve3dCriterion: Shape from GeomAbs;
    myCurve2dCriterion: Shape from GeomAbs;
    mySurfaceCriterion : Shape from GeomAbs;
    myTolerance3d: Real;
    myTolerance2d: Real;

end ShapeDivideContinuity;
