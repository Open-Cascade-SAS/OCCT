-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class NamedUnit from StepBasic 

inherits TShared from MMgt


  -- N.B : EXPRESS Complexe SUBTYPE Declaration :

  -- ANDOR ( ONEOF ( si_unit conversion_based_unit ) ONEOF ( length_unit plane_angle_unit ) ) 

uses

	DimensionalExponents from StepBasic
is

	Create returns mutable NamedUnit;
	---Purpose: Returns a NamedUnit

	Init (me : mutable;
	      aDimensions : mutable DimensionalExponents from StepBasic) is virtual;

	-- Specific Methods for Field Data Access --

	SetDimensions(me : mutable; aDimensions : mutable DimensionalExponents) 
    	is virtual;

	Dimensions (me) returns mutable DimensionalExponents
    	is virtual;

fields

	dimensions : DimensionalExponents from StepBasic;

end NamedUnit;
