-- Created on: 2000-05-10
-- Created by: Andrey BETENEV
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1

class ExternallyDefinedGeneralProperty from StepAP214
inherits GeneralProperty from StepBasic

    ---Purpose: Representation of STEP entity ExternallyDefinedGeneralProperty

uses
    HAsciiString from TCollection,
    SourceItem from StepBasic,
    ExternalSource from StepBasic,
    ExternallyDefinedItem from StepBasic

is
    Create returns ExternallyDefinedGeneralProperty from StepAP214;
	---Purpose: Empty constructor

    Init (me: mutable; aGeneralProperty_Id: HAsciiString from TCollection;
                       aGeneralProperty_Name: HAsciiString from TCollection;
                       hasGeneralProperty_Description: Boolean;
                       aGeneralProperty_Description: HAsciiString from TCollection;
                       aExternallyDefinedItem_ItemId: SourceItem from StepBasic;
                       aExternallyDefinedItem_Source: ExternalSource from StepBasic);
	---Purpose: Initialize all fields (own and inherited)

    ExternallyDefinedItem (me) returns ExternallyDefinedItem from StepBasic;
	---Purpose: Returns data for supertype ExternallyDefinedItem
    SetExternallyDefinedItem (me: mutable; ExternallyDefinedItem: ExternallyDefinedItem from StepBasic);
	---Purpose: Set data for supertype ExternallyDefinedItem

fields
    theExternallyDefinedItem: ExternallyDefinedItem from StepBasic; -- supertype

end ExternallyDefinedGeneralProperty;
