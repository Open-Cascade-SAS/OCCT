-- Created on: 1992-09-23
-- Created by: Christian CAILLET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ExternalSources  from IFGraph  inherits GraphContent

    	---Purpose : this class gives entities which are Source of entities of
    	--           a sub-part, but are not contained by this sub-part

uses Transient, EntityIterator, Graph

is

    Create (agraph : Graph) returns ExternalSources;
    ---Purpose : creates empty ExternalSources, ready to work

    GetFromEntity (me : in out; ent : any Transient);
    ---Purpose : adds an entity and its shared ones to the list

    GetFromIter (me : in out; iter : EntityIterator);
    ---Purpose : adds a list of entities (as an iterator) with shared ones

    ResetData (me : in out);
    ---Purpose : Allows to restart on a new data set

    	-- --   Results   -- --
    	--   More-Next-Value give External Source entities

    Evaluate (me : in out) is redefined;
    ---Purpose : Evaluates external sources of a set of entities

    IsEmpty(me : in out) returns Boolean;
    ---Purpose : Returns True if no External Source are found
    --           It means that we have a "root" set
    --           (performs an Evaluation as necessary)

fields

    thegraph : Graph;

end ExternalSources;
