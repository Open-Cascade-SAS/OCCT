-- Created on: 2009-04-06
-- Created by: Sergey ZARITCHNY
-- Copyright (c) 2009-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Plane from TDataXtd inherits Attribute from TDF

    	
	---Purpose: The basis to define a plane attribute.
    	--  Warning:  Use TDataXtd_Geometry  attribute  to retrieve  the
	--          gp_Pln of the Plane attribute

uses Attribute       from TDF,
     Label           from TDF,
     GUID            from Standard,
     Label           from TDF,
     Plane           from Geom,
     Pln             from gp,
     DataSet         from TDF,
     RelocationTable from TDF

is    

    ---Purpose: class methods
    --          =============
   
    GetID (myclass)    
    	---C++: return const & 
    returns GUID from Standard;
    	---Purpose:
    	-- Returns the GUID for plane attributes.

    Set (myclass ; label : Label from TDF)    
    	---Purpose:  Finds or creates the plane attribute defined by
    	-- the label label.
    	-- Warning
    	-- If you are creating the attribute with this syntax, a
    	-- planar face should already be associated with label.
    returns Plane from TDataXtd;    

    Set (myclass ; label : Label from TDF; P : Pln from gp)
    	---Purpose: Finds,  or creates,  a Plane  attribute  and sets <P>  as
    	--          generated the associated NamedShape.
    returns Plane from TDataXtd;    


    ---Purpose: Plane methods
    --         =============    

    Create
    returns mutable Plane from TDataXtd;  
    
    ---Category: TDF_Attribute methods
    --           =====================
    
    ID (me)  
    	---C++: return const & 
    returns GUID from Standard;

    Restore (me: mutable; With : Attribute from TDF);

    NewEmpty (me)
    returns mutable Attribute from TDF;

    Paste (me; Into : mutable Attribute from TDF;
	       RT   : mutable RelocationTable from TDF);  

    Dump (me; anOS : in out OStream from Standard)
    	returns OStream from Standard
    	is redefined;
	---C++: return &

end Plane;


