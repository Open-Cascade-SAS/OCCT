-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class OrientedEdge from StepShape 

inherits Edge from StepShape 

uses

	Boolean from Standard, 
	Vertex from StepShape, 
	HAsciiString from TCollection
is

	Create returns mutable OrientedEdge;
	---Purpose: Returns a OrientedEdge
	

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aEdgeElement : mutable Edge from StepShape;
	      aOrientation : Boolean from Standard) is virtual;

	-- Specific Methods for Field Data Access --

	SetEdgeElement(me : mutable; aEdgeElement : mutable Edge);
	EdgeElement (me) returns mutable Edge;
	SetOrientation(me : mutable; aOrientation : Boolean);
	Orientation (me) returns Boolean;
	SetEdgeStart(me : mutable; aEdgeStart : mutable Vertex) is redefined;
	EdgeStart (me) returns mutable Vertex is redefined;
	SetEdgeEnd(me : mutable; aEdgeEnd : mutable Vertex) is redefined;
	EdgeEnd (me) returns mutable Vertex is redefined;

fields

	edgeElement : Edge from StepShape;
	orientation : Boolean from Standard;

 -- 
 -- NB : field <edge_start> inherited from classe <edge> is redeclared.
 --      it shall appears in a physical file as a *.
 --

 -- 
 -- NB : field <edge_end> inherited from classe <edge> is redeclared.
 --      it shall appears in a physical file as a *.
 --

end OrientedEdge;
