-- Created on: 1995-02-13
-- Created by: Mister rmi
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Modified by ROB : Wed Oct 98 
--               Add One Method : RecomputeSelection 
--               Modification of Update Method (just computes the 
--               flagged selections)


class SelectionManager from SelectMgr inherits TShared from MMgt

  ---Purpose: A framework to manage selection from the point of
      -- view of viewer selectors. These can be added and
      -- removed, and selection modes can be activated and
      -- deactivated. In addition, objects may be known to all
      -- selectors or only to some.

uses
    AsciiString              from TCollection,
    ViewerSelector           from SelectMgr,
    SelectableObject         from SelectMgr,
    CString                  from Standard,
    MapOfTransient           from TColStd,
    TypeOfUpdate             from SelectMgr,
    DataMapOfObjectSelectors from SelectMgr
    

is


    Create returns SelectionManager from SelectMgr;
    --- Purpose: Constructs an empty selection manager object.

    ---Category: Management of the view selectors


    Add (me          : mutable;
         theSelector : ViewerSelector from SelectMgr)
      is static;
          ---Purpose: Adds the viewer selector theSelector to the list of known items.
    
    Remove (me          : mutable;
            theSelector : ViewerSelector from SelectMgr)
      is static;
    ---Purpose: Removes viewer selector theSelector from the list of known items.
    
    Contains (me;
              theSelector : ViewerSelector from SelectMgr)
      returns Boolean
      is static;
    ---Purpose: Returns true if the manager contains the viewer selector theSelector in a list of known items.

    Contains (me;
              theObject : SelectableObject from SelectMgr)
      returns Boolean
      is static;
    ---Purpose: Returns true if the manager contains the selectable object theObject.





    Load (me        : mutable;
          theObject : SelectableObject from SelectMgr;
          theMode   : Integer = -1)
      is static;
    ---Purpose: Loads and computes selection mode theMode (if it is not equal to -1) in global context and adds selectable
    -- object to BVH tree. If the object theObject has an already calculated selection with mode theMode and it was removed,
    -- the selection will be recalculated.

    Load (me          : mutable;
          theObject   : SelectableObject from SelectMgr;
          theSelector : ViewerSelector from SelectMgr;
          theMode     : Integer = -1)
      is static;
    ---Purpose: Loads and computes selection mode theMode (if it is not equal to -1) and adds selectable object to BVH tree.
    -- Does not perform check of existance of theObject in global context before addition, but adds theSelector to local context.


    Remove (me        : mutable;
            theObject : SelectableObject from SelectMgr)
      is static;
    ---Purpose: Removes selectable object theObject from all viewer selectors it was added to previously, removes it from all contexts
    -- and clears all computed selections of theObject.


    Remove (me          : mutable;
            theObject   : SelectableObject from SelectMgr;
            theSelector : ViewerSelector from SelectMgr)
      is static;
    ---Purpose: Removes theObject from theSelector, does not clear selections and unbind theObject from context maps.





    Activate (me          : mutable;
              theObject   : SelectableObject from SelectMgr;
              theMode     : Integer = 0;
              theSelector : ViewerSelector from SelectMgr = NULL)
      is static;
    ---Purpose: Activates the selection mode theMode in the selector theSelector for the selectable object anObject.
    -- By default, theMode is equal to 0. If theSelector is set to default (NULL), the selection with the mode theMode
    -- will be activated in all the viewers available.

    Deactivate (me          : mutable;
                theObject   : SelectableObject from SelectMgr;
                theMode     : Integer = -1;
                theSelector : ViewerSelector from SelectMgr = NULL);
    ---Purpose: Deactivates mode theMode of theObject in theSelector. If theMode value is set to default (-1), all
    -- avtive selection modes will be deactivated. Likewise, if theSelector value is set to default (NULL), theMode
    -- will be deactivated in all viewer selectors.

    
    IsActivated (me;
                 theObject   : SelectableObject from SelectMgr;
                 theMode     : Integer = -1;
                 theSelector : ViewerSelector from SelectMgr = NULL)
      returns Boolean from Standard;
    ---Purpose: Returns true if the selection with theMode is active for the selectable object theObject and selector theSelector.
    -- If all parameters are set to default values, it returns it there is any active selection in any known viewer selector for
    -- object theObject.





    ClearSelectionStructures (me          : mutable;
                              theObj      : SelectableObject from SelectMgr;
                              theMode     : Integer from Standard = -1;
                              theSelector : ViewerSelector from SelectMgr = NULL)
         is static;
    ---Purpose: Removes sensitive entities from all viewer selectors
    -- after method Clear() was called to the selection they belonged to
    -- or it was recomputed somehow.

    RestoreSelectionStructures (me          : mutable;
                                theObj      : SelectableObject from SelectMgr;
                                theMode     : Integer from Standard = -1;
                                theSelector : ViewerSelector from SelectMgr = NULL)
         is static;
    ---Purpose: Re-adds newely calculated sensitive  entities of recomputed selection
    -- defined by mode theMode to all viewer selectors contained that selection.





    RecomputeSelection (me         : mutable;
                        theObject  : SelectableObject from SelectMgr;
                        theIsForce : Boolean from Standard  = Standard_False;
                        theMode    : Integer from Standard = -1);
    ---Purpose: Recomputes activated selections of theObject for all known viewer selectors according to theMode specified.
    -- If theMode is set to default (-1), then all activated selections will be recomputed. If theIsForce is set to true,
    -- then selection mode theMode for object theObject will be recomputed regardless of its activation status.


    Update (me         : mutable;
            theObject  : SelectableObject from SelectMgr;
            theIsForce : Boolean from Standard = Standard_True)
      is static;
    ---Purpose: Updates all selections of theObject in all viewer selectors according to its current update status.
    -- If theIsForce is set to true, the call is equal to recomputation.

    Update (me          : mutable;
            theObject   : SelectableObject from SelectMgr;
            theSelector : ViewerSelector from SelectMgr;
            theIsForce  : Boolean from Standard = Standard_True)
      is static;
    ---Purpose: Updates all selections of theObject in specified viewer selector according to its current update status.
    -- If theIsForce is set to true, the call is equal to recomputation.





    SetUpdateMode (me        : mutable;
                   theObject : SelectableObject from SelectMgr;
                   theType   : TypeOfUpdate from SelectMgr)
      is static;
    ---Purpose: Sets type of update of all selections of theObject to the given theType.


    SetUpdateMode (me        : mutable;
                   theObject : SelectableObject from SelectMgr;
                   theMode   : Integer from Standard;
                   theType   : TypeOfUpdate    from SelectMgr)
      is static;
    ---Purpose: Sets type of update of selection with theMode of theObject to the given theType.





    loadMode (me          : mutable;
              theObject   : SelectableObject from SelectMgr;
              theMode     : Integer;
              theSelector : ViewerSelector from SelectMgr = NULL)
      is static private;
    ---Purpose: Loads and creates selection structures for object theObject with mode theMode in specified
    -- viewer selector theSelector. If theSelector is set to default value (NULL), the selection mode
    -- created will be added to all known viewer selectors.

    rebuildSelectionStructures (me          : mutable;
                                theSelector : ViewerSelector from SelectMgr = NULL)
      is static private;
    ---Purpose: Internal function that marks 1st level BVH of the object theObj as
    -- outdated.





fields

    -- myselectors : selectors dedicated to one particular view;
    -- myglobal    : objects which will be selectable in all the views
    -- mylocal     : objects with the selectors where they are selectable


    mySelectors : MapOfTransient           from TColStd;
    myGlobal    : MapOfTransient           from TColStd;
    myLocal     : DataMapOfObjectSelectors from SelectMgr;


end SelectionManager;



