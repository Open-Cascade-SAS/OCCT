-- Created on: 1995-04-05
-- Created by: Christophe MARION
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Projector from HLRTest inherits Drawable3D from Draw
	---Purpose: 

uses
    OStream,
    Display     from Draw,
    Interpretor from Draw,
    Projector   from HLRAlgo

is
    Create(P : Projector from HLRAlgo)
    returns mutable Projector from HLRTest; 
    
    Projector(me) returns Projector from HLRAlgo;
	---C++: return const &
	---C++: inline

    DrawOn(me; dis : in out Display from Draw);
	---Purpose: Does nothhing,
    
    Copy(me) returns mutable Drawable3D from Draw
	---Purpose: For variable copy.
    is redefined;
	
    Dump(me; S : in out OStream)
	---Purpose: For variable dump.
    is redefined;

    Whatis(me; I : in out Interpretor from Draw)
	---Purpose: For variable whatis command. Set  as a result  the
	--          type of the variable.
    is redefined;

fields
    myProjector : Projector from HLRAlgo;

end Projector;
