-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class WeekOfYearAndDayDate from StepBasic 

inherits Date from StepBasic 

uses

	Integer from Standard, 
	Boolean from Standard
is

	Create returns WeekOfYearAndDayDate;
	---Purpose: Returns a WeekOfYearAndDayDate


	Init (me : mutable;
	      aYearComponent : Integer from Standard) is redefined;

	Init (me : mutable;
	      aYearComponent : Integer from Standard;
	      aWeekComponent : Integer from Standard;
	      hasAdayComponent : Boolean from Standard;
	      aDayComponent : Integer from Standard) is virtual;

	-- Specific Methods for Field Data Access --

	SetWeekComponent(me : mutable; aWeekComponent : Integer);
	WeekComponent (me) returns Integer;
	SetDayComponent(me : mutable; aDayComponent : Integer);
	UnSetDayComponent (me:mutable);
	DayComponent (me) returns Integer;
	HasDayComponent (me) returns Boolean;

fields

	weekComponent : Integer from Standard;
	dayComponent : Integer from Standard;   -- OPTIONAL can be NULL
	hasDayComponent : Boolean from Standard;

end WeekOfYearAndDayDate;
