-- Created on: 1993-04-28
-- Created by: Laurent PAINNOT
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



deferred generic class TheSurfTool from AppCont(Surf as any)

    ---Purpose: Template for describing a continuous surface.


uses Pnt           from gp,
     Vec           from gp

is


    D0(myclass; S: Surf; U, V: Real; Pt: out Pnt);
    	---Purpose: returns the point of the surface at <U, V>.


    D1(myclass; S: Surf; U, V: Real; Pt: out Pnt; V1U, V1V: out Vec);
    	---Purpose: returns the derivative and the point values of the surface
    	--          at the parameters <U, V> .

end TheSurfTool;
