-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class BoxedHalfSpace from StepShape 

inherits HalfSpaceSolid from StepShape 

uses

	BoxDomain from StepShape, 
	HAsciiString from TCollection, 
	Surface from StepGeom, 
	Boolean from Standard
is

	Create returns mutable BoxedHalfSpace;
	---Purpose: Returns a BoxedHalfSpace


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aBaseSurface : mutable Surface from StepGeom;
	      aAgreementFlag : Boolean from Standard) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aBaseSurface : mutable Surface from StepGeom;
	      aAgreementFlag : Boolean from Standard;
	      aEnclosure : mutable BoxDomain from StepShape) is virtual;

	-- Specific Methods for Field Data Access --

	SetEnclosure(me : mutable; aEnclosure : mutable BoxDomain);
	Enclosure (me) returns mutable BoxDomain;

fields

	enclosure : BoxDomain from StepShape;

end BoxedHalfSpace;
