-- File:	ShapeFix_ComposeShell.cdl
-- Created:	Mon Apr 26 19:04:10 1999
-- Author:	Andrey BETENEV
--		<abv@doomox.nnov.matra-dtv.fr>
---Copyright:	 Matra Datavision 1999


class ComposeShell from ShapeFix inherits Root from ShapeFix

	---Purpose: This class is intended to create a shell from the composite
	--          surface (grid of surfaces) and set of wires.
	--          It may be either division of the supporting surface of the 
        --          face, or creating a shape corresponding to face on composite
	--          surface which is missing in CAS.CADE but exists in some other 
        --          systems.
	--
	--          It splits (if necessary) original face to several ones by
	--          splitting lines which are joint lines on a supplied grid of
	--          surfaces (U- and V- isolines of the  composite surface).
	--          There are two modes of work, which differ in the way of 
	--          handling faces on periodic surfaces:
	--
	--        - if ClosedMode is False (default), when splitting itself is
	--          done as if surface were not periodic. The periodicity of the 
	--          underlying surface is taken into account by duplicating splitting
	--          lines in the periodic direction, as necessary to split all
	--          the wires (whole parametrical range of a face)
	--          In this mode, some regularization procedures are performed
	--          (indexation of splitted segments by patch numbers), and it is 
        --          expected to be more reliable and robust in case of bad shapes
	--
	--        - if ClosedMode is True, when everything on a periodic surfaces
        --          is considered as modulo period. This allows to deal with wires
	--          which are closed in 3d but not in 2d, with wires which may be
        --          shifted on several periods in 2d etc. However, this mode is 
        --          less reliable since some regularizations do not work for it.
	--
	--          The work is made basing on pcurves of the edges. These pcurves
	--          should already exist (for example, in the case of division of 
	--          existing face), then they are taken as is. The existing pcurves
	--          should be assigned to one surface (face) for all edges,
	--          this surface (face) will be used only for accessing pcurves,
	--          and it may have any geometry.
    	--
        --          All the modifications are recorded in the context tool
        --          (ShapeBuild_ReShape).

uses
    Lin2d    from gp,
    Curve    from Geom2d,
    Surface  from Geom,
    Location from TopLoc,
    Edge     from TopoDS,
    Face     from TopoDS,
    Shape    from TopoDS, 
    Status   from ShapeExtend,
    WireData from ShapeExtend,
    CompositeSurface from ShapeExtend,
    WireSegment      from ShapeFix,
    Orientation      from TopAbs,
    SequenceOfReal        from TColStd,
    SequenceOfInteger     from TColStd,
    SequenceOfShape       from TopTools,
    SequenceOfWireSegment from ShapeFix,
    TransferParameters    from ShapeAnalysis
is
    Create returns ComposeShell from ShapeFix;
        ---Purpose: Creates empty tool.
    
    Init (me: mutable; Grid: CompositeSurface from ShapeExtend;
    	    	       L   : Location from TopLoc;
                       Face: Face from TopoDS;
    	    	       Prec: Real);
        ---Purpose: Initializes with composite surface, face and precision.
	--          Here face defines both set of wires and way of getting
	--          pcurves. Precision is used (together with tolerance of edges)
	--          for handling subtle cases, such as tangential intersections.

    ClosedMode (me: mutable) returns Boolean;
    	---Purpose: Returns (modifiable) flag for special 'closed'
	--          mode which forces ComposeShell to consider
	--          all pcurves on closed surface as modulo period.
	--          This can reduce reliability, but allows to deal
	--          with wires closed in 3d but open in 2d (missing seam)
	--          Default is False
	---C++: return &
		      
    Perform (me: mutable) 
    returns Boolean is virtual;
        ---Purpose: Performs the work on already loaded data.

    SplitEdges (me: mutable);
    	---Purpose: Splits edges in the original shape by grid.
	--          This is a part of Perform() which does not produce any
        --          resulting shape; the only result is filled context
	--          where splittings are recorded.
	--
	--          NOTE: If edge is splitted, it is replaced by wire, and 
	--          order of edges in the wire corresponds to FORWARD orientation
	--          of the edge.
    
    Result (me) returns Shape from TopoDS;
        ---Purpose: Returns resulting shell or face (or Null shape if not done)
    	---C++: return const &
    
    Status (me; status: Status from ShapeExtend) returns Boolean;
        ---Purpose: Queries status of last call to Perform()
	-- OK   : nothing done (some kind of error)
	-- DONE1: splitting is done, at least one new face created
	-- DONE2: splitting is done, several new faces obtained
	-- FAIL1: misoriented wire encountered (handled)
	-- FAIL2: recoverable parity error
	-- FAIL3: edge with no pcurve on supporting face
	-- FAIL4: unrecoverable algorithm error (parity check)
    
    ---Protected methods:
    
    LoadWires (me; seqw: out SequenceOfWireSegment from ShapeFix)
    is protected;
    	---Purpose: Fill sequence of wire segments by wires from myFace
	--          (pre-loaded). It performs reorder so that edges in segments
	--          are well-ordered. The context is applied to all wires
	--          before using them.
    
    ComputeCode (me: mutable; wire  : WireData from ShapeExtend;
			      line  : Lin2d from gp;
		    	      begInd: Integer;
		    	      endInd: Integer;
       		    	      begPar: Real;
		    	      endPar: Real;
    	    	    	      IsInternal : Boolean = Standard_False)
    returns Integer is protected;
    	---Purpose: Analyze tangencies and compute orientation code for wire segment 
    	--          between two intersections: tells if segment is on left or right side 
	--          of cutting line, or tangent to it (by several points recomputed to 3d, 
	--          distance is compared with tolerance of corresponding edge).

    SplitWire (me: mutable; wire    : in out WireSegment from ShapeFix;
    	    	            indexes : in out SequenceOfInteger from TColStd;
		            values  : SequenceOfReal    from TColStd;
    	    	            vertices: out SequenceOfShape from TopTools;
			    segcodes: SequenceOfInteger from TColStd;
			    cutbyu  : Boolean;
			    cutindex: Integer)
    returns WireSegment from ShapeFix is protected;
    	---Purpose: Splits edges in the wire by given indices of edges and 
	--          parameters on them. Returns resulting wire and vertices 
	--          corresponding to splitting parameters. If two consequtive
	--          splitting points are too near one to another (with tolerance 
	--          of edge), edge is divided in single point. In the same way,
	--          splitting which is too near to end of edge, is not applied
	--          (end vertex is returned instead).
	--
	--          NOTE: If edge is splitted, it is replaced by wire, and 
	--          order of edges in the wire corresponds to FORWARD orientation
	--          of the edge.
	
    SplitByLine (me: mutable; wire           : in out WireSegment from ShapeFix;
    	    	              line           : Lin2d from gp;
			      cutbyu  : Boolean;
			      cutindex: Integer;
		     	      SplitLinePar   : out SequenceOfReal from TColStd;
		     	      SplitLineCode  : out SequenceOfInteger from TColStd;
		      	      SplitLineVertex: out SequenceOfShape from TopTools)
    returns Boolean is protected;
        ---Purpose: Split edges in the wire by cutting line.
	--          Wires with FORWARD or REVERSED orientation are considered
	--          as closed.
	--
	--          All modifications (splitting) are recorded in context, 
        --          except splitting of wires marked as EXTERNAL
	--          (they are supposed to be former cutting lines).
	--
	--          Method fills sequences of parameters of intersection points 
	--          of cutting line with all edges, their types, and corresponding
	--          vertices (including ones created during splitting edges).
    
    SplitByLine (me: mutable; seqw: in out SequenceOfWireSegment from ShapeFix;
                              line: Lin2d from gp;
			      cutbyu  : Boolean;
			      cutindex: Integer)
    is protected;
        ---Purpose: Split edges in the sequence of wires by cutting line.
	--          Wires with FORWARD or REVERSED orientation are considered
	--          as closed.
	--
	--          Parts of cutting line which get inside the face (defined by 
        --          parity check of intersections with all wires) are added 
        --          into that sequence (with orientation EXTERNAL). Each part
	--          is represented by one-edge wire segment with no 3d curve.
	--          They share common vertices with all wires they intersect.
        --          
	--          All modifications (splitting) are recorded in context, 
        --          except splitting of wires marked as EXTERNAL
	--          (they are supposed to be former cutting lines).
    
    SplitByGrid (me: mutable; seqw: in out SequenceOfWireSegment from ShapeFix)
    is protected;
        ---Purpose: Split initial set of (closed) wires by grid of lines corresponding 
	--          to joints between patches on the composite surface.
	--          Parts of joint lines which get inside the face are also added
	--          into the sequence as wires with orientation EXTERNAL.
	--          They share common vertices with all wires they intersect.
	--          All modifications (splitting) are recorded in context, 
        --          except splitting of joint edge itself and wires marked as
	--          EXTERNAL (they supposed to be another joint edges).
    
    BreakWires (me: mutable; seqw: in out SequenceOfWireSegment from ShapeFix)
    is protected;
        ---Purpose: Break wires into open wire segments by common vertices
	--          (splitting points), so that each segment is either closed and 
	--          not touching others, or touches others at ends (have common 
	--          vertices). 
        --          After that, each wire segment lies on its own patch of grid.
    
    CollectWires (me: mutable; wires: out SequenceOfWireSegment from ShapeFix;
    	    	               seqw : in out SequenceOfWireSegment from ShapeFix )
    is protected;
        ---Purpose: Collect set of wire segments (already splitted) into closed 
	--          wires. This is done by traversing all the segments in allowed
	--          directions, starting only from the REVERSED and FORWARD and
	--          taking EXTERNAL as necessary in fork points. Forks are detected
	--          by common vertices. In fork point, most left way is seleccted
        --          among all possible ways.
  
    MakeFacesOnPatch (me; faces: out SequenceOfShape from TopTools;
    	    	    	  surf : Surface from Geom;
			  loops: in out SequenceOfShape from TopTools)
    is protected;
    	---Purpose: Creates new faces on one path of grid. It dispatches given loops
	--          (wires) into one or several faces depending on their mutual
	--          position.
    
    DispatchWires (me; faces  : out SequenceOfShape from TopTools;
    	    	       wires  : in out SequenceOfWireSegment from ShapeFix);
        ---Purpose: Creates new faces from the set of (closed) wires. Each wire 
	--          is put on corresponding patch in the composite surface,
	--          and all pcurves on the initial (pseudo)face are reassigned to
	--          that surface. If several wires are one inside another, single
	--          face is created.
    
    SetTransferParamTool(me: mutable; TransferParam : TransferParameters from ShapeAnalysis);
    ---Purpose: Sets tool for transfer parameters from 3d to 2d and vice versa.
	
    GetTransferParamTool(me) returns TransferParameters from ShapeAnalysis; 
    ---Purpose: Gets tool for transfer parameters from 3d to 2d and vice versa.

fields

    myGrid     : CompositeSurface from ShapeExtend;
    myLoc      : Location from TopLoc;
    myFace     : Face from TopoDS;  -- underlying face for pcurves (real or pseudo)
    myOrient   : Orientation from TopAbs is protected;  -- orientation of face
    myResult   : Shape from TopoDS is protected;
    myStatus   : Integer is protected;
    myUResolution: Real;  -- summary resolution on grid (minimum on patches)
    myVResolution: Real;
    myTransferParamTool: TransferParameters from ShapeAnalysis;
    myInvertEdgeStatus : Boolean;
    myClosedMode       : Boolean;
    myUClosed  : Boolean;
    myVClosed  : Boolean;
    myUPeriod  : Real;
    myVPeriod  : Real;
    
end ComposeShell;
