-- Created on: 1997-10-28
-- Created by: Roman BORISOV
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Curve2d from Approx 

	---Purpose: Makes  an  approximation  for  HCurve2d  from  Adaptor3d

uses
    HCurve2d    from  Adaptor2d, 
    Shape  from  GeomAbs, 
    BSplineCurve  from  Geom2d 
    
is
  Create(C2D  :  HCurve2d    from  Adaptor2d; 
    	 First, 
	 Last, 		      
         TolU,  TolV  :  Real; 
	 Continuity  :  Shape  from  GeomAbs; 
         MaxDegree  :  Integer  ; 
         MaxSegments  :  Integer) 
	      
     returns  Curve2d;	 
      
    IsDone(me) returns Boolean from Standard;
    
    HasResult(me) returns  Boolean from Standard;
   
    Curve(me) 
    returns  BSplineCurve  from  Geom2d; 
     
    MaxError2dU(me) returns  Real;  
    MaxError2dV(me) returns  Real;
    
fields
   
  myCurve            : BSplineCurve  from  Geom2d; 
  myIsDone           : Boolean       from  Standard;   
  myHasResult        : Boolean       from  Standard; 
  myMaxError2dU      : Real          from  Standard; 
  myMaxError2dV      : Real          from  Standard; 
  
end Curve2d;
