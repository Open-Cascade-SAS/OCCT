-- Created on: 1999-03-10
-- Created by: data exchange team
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PresentedItemSelect from StepAP214 
inherits SelectType from StepData
	
uses
     ProductDefinition from StepBasic,
     ProductDefinitionRelationship from StepBasic


is

    Create returns PresentedItemSelect;
	---Purpose : Returns a PresentedItemSelect SelectType

    CaseNum (me; ent : Transient) returns Integer;
	---Purpose: Recognizes a PresentedItemSelect Kind Entity that is :
	--  1 -> ProductDefinition,
	--  2 -> ProductDefinitionRelationship,
	--        0 else

    ProductDefinitionRelationship (me) returns any ProductDefinitionRelationship;
    ---Purpose : returns Value as a ProductDefinitionRelationship (Null if another type)

    ProductDefinition (me) returns any ProductDefinition;
    ---Purpose : returns Value as a ProductDefinition (Null if another type)

end PresentedItemSelect;
