-- File:        Approval.cdl
-- Created:     Fri Dec  1 11:11:13 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class Approval from StepBasic 

inherits TShared from MMgt

uses

	ApprovalStatus from StepBasic, 
	HAsciiString from TCollection
is

	Create returns mutable Approval;
	---Purpose: Returns a Approval

	Init (me : mutable;
	      aStatus : mutable ApprovalStatus from StepBasic;
	      aLevel : mutable HAsciiString from TCollection) is virtual;

	-- Specific Methods for Field Data Access --

	SetStatus(me : mutable; aStatus : mutable ApprovalStatus);
	Status (me) returns mutable ApprovalStatus;
	SetLevel(me : mutable; aLevel : mutable HAsciiString);
	Level (me) returns mutable HAsciiString;

fields

	status : ApprovalStatus from StepBasic;
	level : HAsciiString from TCollection;

end Approval;
