-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class DateAndTimeAssignment from StepBasic 

inherits TShared from MMgt

uses

	DateAndTime from StepBasic, 
	DateTimeRole from StepBasic
is

	Init (me : mutable;
	      aAssignedDateAndTime : mutable DateAndTime from StepBasic;
	      aRole : mutable DateTimeRole from StepBasic) is virtual;

	-- Specific Methods for Field Data Access --

	SetAssignedDateAndTime(me : mutable; aAssignedDateAndTime : mutable DateAndTime);
	AssignedDateAndTime (me) returns mutable DateAndTime;
	SetRole(me : mutable; aRole : mutable DateTimeRole);
	Role (me) returns mutable DateTimeRole;

fields

	assignedDateAndTime : DateAndTime from StepBasic;
	role : DateTimeRole from StepBasic;

end DateAndTimeAssignment;
