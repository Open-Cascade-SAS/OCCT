-- Created on: 1991-10-10
-- Created by: Jean Claude VAUTHIER
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.






class EllipseToBSplineCurve   from Convert   inherits ConicToBSplineCurve

        --- Purpose :
        --  This algorithm converts a ellipse into a rational B-spline curve.
        --  The ellipse is represented an Elips2d from package gp with
        --  the parametrization :
        --  P (U) = 
        --  Loc + (MajorRadius * Cos(U) * Xdir + MinorRadius * Sin(U) * Ydir)
        --  where Loc is the center of the ellipse, Xdir and Ydir are the 
        --  normalized directions of the local cartesian coordinate system of
        --  the ellipse. The parametrization range is U [0, 2PI].
        --- KeyWords :
        --  Convert, Ellipse, BSplineCurve, 2D .

uses Elips2d              from gp,
     ParameterisationType from Convert

raises DomainError from Standard

is

  Create (E : Elips2d;
    	   Parameterisation : ParameterisationType from Convert 
    	    = Convert_TgtThetaOver2 )   returns EllipseToBSplineCurve;
        --- Purpose : The equivalent B-spline curve has the same orientation
        --  as the ellipse E.


  Create (E : Elips2d; U1, U2 : Real;
           Parameterisation : ParameterisationType from Convert 
    	    = Convert_TgtThetaOver2 )   returns EllipseToBSplineCurve
        --- Purpose : 
        --  The ellipse E is limited between the parametric values U1, U2.
        --  The equivalent B-spline curve is oriented from U1 to U2 and has
        --  the same orientation as E.
     raises DomainError;
        --- Purpose :
        --  Raised if U1 = U2 or U1 = U2 + 2.0 * Pi



end EllipseToBSplineCurve;

