-- Created by: Peter KURNEV
-- Copyright (c) 2010-2014 OPEN CASCADE SAS
-- Copyright (c) 2007-2010 CEA/DEN, EDF R&D, OPEN CASCADE
-- Copyright (c) 2003-2007 OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN, CEDRAT,
--                         EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class BuilderFace from BOPAlgo 
    	inherits BuilderArea from BOPAlgo 
	 
	---Purpose: The algorithm to build faces from set of edges  

uses    
    Orientation from TopAbs,
    Face from TopoDS,
    BaseAllocator from BOPCol 
--raises

is 
    Create  
    	returns BuilderFace from BOPAlgo; 
    ---C++: alias "Standard_EXPORT virtual ~BOPAlgo_BuilderFace();" 
      
    Create (theAllocator: BaseAllocator from BOPCol)  
    	returns BuilderFace from BOPAlgo;  
	
    SetFace(me:out; 
            theFace:Face from TopoDS);  
    ---Purpose: Sets the face generatix  
	 
    Face(me) 
    ---Purpose: Returns the face generatix   
    	returns Face from TopoDS; 
    ---C++:  return const &
		 
    Perform(me:out)  
    	---Purpose:  Performs the algorithm 
    	is redefined;  
	 
    PerformShapesToAvoid(me:out) 
	---Purpose:  Collect the edges that 
	--           a) are internal        	 
	--           b) are the same and have different orientation         	 
    	is redefined protected; 
	 
    PerformLoops(me:out) 
	---Purpose: Build draft wires 
        --          a)myLoops - draft wires that consist of  
        --                       boundary edges 
	--          b)myLoopsInternal - draft wires that contains 
	--                               inner edges 
    	is redefined protected;  
	 
    PerformAreas(me:out)   
    	---Purpose: Build draft faces that contains boundary edges 
    	is redefined protected;  

    PerformInternalShapes(me:out)   
    	---Purpose: Build finalized faces with internals   
    	is redefined protected;  
     
    CheckData(me:out) 
	is redefined protected;   
     
    Orientation(me) 
    	returns Orientation from TopAbs; 
 
fields  
    myFace : Face from TopoDS is protected;     
    myOrientation: Orientation from TopAbs is protected;   	      
 
end BuilderFace; 

