-- Created on: 1996-12-16
-- Created by: Christian CAILLET
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Field    from StepData

    ---Purpose : Defines a generally defined Field for STEP data : can be used
    --           either in any kind of entity to implement it or in free format
    --           entities in a "late-binding" mode
    --           A field can have : no value (or derived), a single value of
    --           any kind, a list of value : single or double list
    --           
    --           When a field is set, this defines its new kind (Integer etc..)
    --           A single value is immediately set. A list of value is, firstly
    --           declared as for a kind (Integer String etc), then declared as
    --           a list with its initial size, after this its items are set
    --           Also it can be set in once if the HArray is ready 

uses Transient, HAsciiString, CString,
     HArray1OfInteger from TColStd, HArray1OfReal from TColStd,
     HArray1OfTransient from TColStd, HArray1OfHAsciiString from Interface,
     Logical from StepData, SelectMember from StepData

is

    Create returns Field;
    ---Purpose : Creates a Field, empty ("no value defined")

    Create (other : Field; copy : Boolean = Standard_False)  returns Field;
    ---Purpose : Creates a Field from another one. If <copy> is True, Handled
    --           data (Select,String,List, not entities) are copied

    CopyFrom (me : in out; other : Field);
    ---Purpose : Gets the copy of the values of another field

    Clear (me : in out; kind : Integer = 0);
    ---Purpose : Clears the field, to set it as "no value defined"
    --           Just before SetList, predeclares it as "any"
    --           A Kind can be directly set here to declare a type

    	-- Setting a Single Value, or predeclaring a list

    SetDerived (me : in out);
    ---Purpose : Codes a Field as derived (no proper value)

    SetInt (me : in out; val : Integer);
    ---Purpose : Directly sets the Integer value, if its Kind matches
    --           Integer, Boolean, Logical, or Enum (does not change Kind)

    SetInteger (me : in out; val : Integer = 0);
    ---Purpose : Sets an Integer value (before SetList* declares it as Integer)

    SetBoolean (me : in out; val : Boolean = Standard_False);
    ---Purpose : Sets a Boolean value (or predeclares a list as boolean)

    SetLogical (me : in out; val : Logical = StepData_LFalse);
    ---Purpose : Sets a Logical Value (or predeclares a list as logical)

    SetReal    (me : in out; val : Real = 0.0);
    ---Purpose : Sets a Real    Value (or predeclares a list as Real);

    SetString  (me : in out; val : CString = "");
    ---Purpose : Sets a String  Value (or predeclares a list as String)
    --           Does not redefine the Kind if it is alread String or Enum

    SetEnum    (me : in out; val : Integer = -1; text : CString = "");
    ---Purpose : Sets an Enum Value (as its integer counterpart)
    --           (or predeclares a list as Enum)
    --           If <text> is given , also sets its textual expression
    --           <val> negative means unknown (known values begin at 0)

    SetSelectMember (me : in out; val : SelectMember);
    ---Purpose : Sets a SelectMember (for Integer,Boolean,Enum,Real,Logical)
    --           Hence, the value of the field is accessed through this member

    SetEntity  (me : in out; val : Transient);
    ---Purpose : Sets an Entity Value

    SetEntity  (me : in out);
    ---Purpose : Predeclares a list as of entity

    SetList  (me : in out; size : Integer; first : Integer = 1);
    ---Purpose : Declares a field as a list, with an initial size
    --           Initial lower is defaulted as 1, can be defined
    --           The list starts empty, typed by the last Set*
    --           If no Set* before, sets it as "any" (transient/select)

    SetList2 (me : in out; siz1, siz2 : Integer; f1,f2 : Integer = 1);
    ---Purpose : Declares a field as an homogeneous square list, with initial\
    --           sizes, and initial lowers

    Set (me : in out; val : Transient);
    ---Purpose : Sets an undetermined value : can be String, SelectMember,
    --           HArray(1-2) ... else, an Entity
    --           In case of an HArray, determines and records its size(s)

    	-- Setting List Items : Single List

    ClearItem  (me : in out; num : Integer);
    ---Purpose : Declares an item of the list as undefined
    --           (ignored if list not defined as String,Entity or Any)

    SetInt     (me : in out; num : Integer; val : Integer; kind : Integer);
    ---Purpose : Internal access to an Integer Value for a list, plus its kind

    SetInteger (me : in out; num : Integer; val : Integer);
    ---Purpose : Sets an Integer Value for a list (rank num)
    --           (recognizes a SelectMember)

    SetBoolean (me : in out; num : Integer; val : Boolean);

    SetLogical (me : in out; num : Integer; val : Logical);

    SetEnum    (me : in out; num : Integer; val : Integer; text: CString = "");
    ---Purpose : Sets an Enum Value (Integer counterpart), also its text
    --           expression if known (if list has been set as "any")

    SetReal    (me : in out; num : Integer; val : Real);

    SetString  (me : in out; num : Integer; val : CString);

    SetEntity  (me : in out; num : Integer; val : Transient);

    	-- Quering Value
    	-- For a Single field, n1 and n2 are ignored
    	-- For a Single List, n1 is considered and n2 is ignored

    IsSet (me; n1, n2 : Integer = 1) returns Boolean;

    ItemKind (me; n1, n2 : Integer = 1) returns Integer;
    ---Purpose : Returns the kind of an item in a list or double list
    --           It is the kind of the list, except if it is "Any", in such a
    --           case the true kind is determined and returned

    Kind     (me; type : Boolean = Standard_True) returns Integer;  -- enum ?
    ---Purpose : Returns the kind of the field
    --           <type> True (D) : returns only the type itself
    --           else, returns the complete kind

    Arity    (me) returns Integer;  -- 0:single  1:list  2:list2

    Length   (me; index : Integer = 1) returns Integer;  -- for index 1 or 2
    --  True Length, not simply the reserved one

    Lower    (me; index : Integer = 1) returns Integer;  -- for index 1 or 2

    	-- Single :

    Int (me) returns Integer;  -- the field Integer itself

    Integer  (me; n1, n2 : Integer = 1) returns Integer;

    Boolean  (me; n1, n2 : Integer = 1) returns Boolean;

    Logical  (me; n1, n2 : Integer = 1) returns Logical;

    Real     (me; n1, n2 : Integer = 1) returns Real;

    String   (me; n1, n2 : Integer = 1) returns CString;

    Enum     (me; n1, n2 : Integer = 1) returns Integer;

    EnumText (me; n1, n2 : Integer = 1) returns CString;  -- "" if unknown

    Entity   (me; n1, n2 : Integer = 1) returns Transient;

    Transient (me) returns Transient;  -- the fields itself

fields

    thekind : Integer;
    theint  : Integer;
    thereal : Real;
    theany  : Transient;

end Field;
