-- Created on: 1992-09-29
-- Created by: Didier PIFFAULT
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



generic class InterferencePolyhedron from Intf
    (Polyhedron1  as any;
     ToolPolyhe1  as any;
     Polyhedron2  as any;
     ToolPolyhe2  as any)     -- as ToolPolyhedron(Polyhedron)
    inherits Interference from Intf

	---Purpose: Computes the  interference between two polyhedra or the
	--          self interference of a polyhedron.

uses    Pnt               from gp,
        XYZ               from gp,
    	Box               from Bnd,
    	SectionPoint      from Intf,
    	SeqOfSectionPoint from Intf,
    	SectionLine       from Intf,
    	SeqOfSectionLine  from Intf,
    	TangentZone       from Intf,
    	SeqOfTangentZone  from Intf

is

-- Interface :

    Create          returns InterferencePolyhedron from Intf;
    ---Purpose: Constructs an empty interference of Polyhedron.

    Create         (Obje1  : in Polyhedron1;
    	    	    Obje2  : in Polyhedron2) 
    	            returns InterferencePolyhedron from Intf;
    ---Purpose: Constructs  and computes  an  interference between  the two
    --          Polyhedra.

    Create         (Obje   : in Polyhedron1) 
    	            returns InterferencePolyhedron from Intf;
    ---Purpose: Constructs  and  computes   the self   interference  of   a
    --          Polyhedron.

    Perform        (me     : in out;
    	    	    Obje1  : in Polyhedron1;
    	    	    Obje2  : in Polyhedron2);
    ---Purpose: Computes the interference between the two Polyhedra.

    Perform        (me     : in out;
    	    	    Obje   : in Polyhedron1);
    ---Purpose: Computes the self interference of a Polyhedron.

-- Implementation :

    Interference   (me     : in out;
    	    	    Obje1  : in Polyhedron1)
    	    	    is private;
    Interference   (me     : in out;
    	    	    Obje1  : in Polyhedron1;
     	    	    Obje2  : in Polyhedron2)
    	    	    is private;
    ---Purpose: Compares the bounding volumes between the facets of <Obje1>
    --          and the facets of <Obje2> and intersects the facets when the
    --          bounding volumes have a common part.

    Intersect      (me     : in out;
		    TriF   : in Integer from Standard;
    	    	    Obje1  : in Polyhedron1;
		    TriS   : in Integer from Standard;
    	    	    Obje2  : in Polyhedron2)
    	    	    is private;
    ---Purpose: Computes  the intersection between    the  facet <Tri1>  of
    --          <FirstPol> and the facet <Tri2> of <SecondPol>.

    TangentZoneValue
    	    	   (me;
    	    	    TheTZ  : in out TangentZone from Intf;
		    Obje1  : Polyhedron1;
		    Tri1   : Integer from Standard;
    	    	    Obje2  : Polyhedron2;
    	    	    Tri2   : Integer from Standard)
		    returns Boolean from Standard
    	    	    is private;
    ---Purpose: Computes the  zone of tangence between the  facet <Tri1> of
    --          <FirstPol> and the facet <Tri2> of <SecondPol>.

    CoupleCharacteristics (me: in out;
            FirstPol: Polyhedron1;
            SeconPol: Polyhedron2) is private;
fields
    OI       : Integer from Standard[3]; -- index des sommets de l objet
    TI       : Integer from Standard[3]; -- index des sommets du tool
    dpOpT    : Real from Standard[3, 3]; -- distance point Objet - point Tool
    dpOeT    : Real from Standard[3, 3]; -- distance point Objet - edge  Tool
    deOpT    : Real from Standard[3, 3]; -- distance edge  Objet - point Tool
    voo      : XYZ from gp[3];           -- vecteur point point Obje
    vtt      : XYZ from gp[3];           -- vecteur point point Tool
    Incidence: Real from Standard;       -- angle entre les deux plans

end InterferencePolyhedron;
