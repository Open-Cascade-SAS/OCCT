-- Created on: 1992-08-24
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package IntSurf 

	---Purpose: This package provides resources for
	--          all the packages concerning the intersection
	--          between surfaces. 

        ---Level: Internal
        --
        -- All the methods of all the classes of this package are Internal.
        -- 


uses Standard, MMgt, StdFail, GeomAbs, TCollection, gp, TColgp

is

    class PntOn2S;
    
    imported Allocator;
    
    imported SequenceOfPntOn2S;

    class Couple;

    imported SequenceOfCouple;
    
    
    class LineOn2S;
    
    class Quadric;
    
    class QuadricTool;
    
    class PathPoint;
    
    imported SequenceOfPathPoint;

    class PathPointTool;
    
    class InteriorPoint;
    
    imported SequenceOfInteriorPoint;
    
    class InteriorPointTool;

    class Transition;    

    --amv    
    imported ListOfPntOn2S;
    imported ListIteratorOfListOfPntOn2S;
    
    enumeration TypeTrans is In, Out, Touch, Undecided;
    
    enumeration Situation is Inside, Outside, Unknown;


    MakeTransition(TgFirst,TgSecond: Vec from gp; Normal: Dir from gp;
                   TFirst,TSecond: out Transition from IntSurf);

	---Purpose: Computes the transition of the intersection point
	--          between the two lines.
	--          TgFirst is the tangent vector of the first line.
	--          TgSecond is the tangent vector of the second line.
	--          Normal is the direction used to orientate the cross
	--          product TgFirst^TgSecond.
	--          TFirst is the transition of the point on the first line.
	--          TSecond is the transition of the point on the second line.


end IntSurf;
