-- Created on: 1999-03-11
-- Created by: data exchange team
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SweptFaceSolid from StepShape 
inherits SolidModel from StepShape
	
uses
    	HAsciiString from TCollection,
    	FaceSurface from StepShape

is
    	Create returns mutable SweptFaceSolid;
	---Purpose: Returns a SweptFaceSolid


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aSweptArea : mutable FaceSurface from StepShape) is virtual;

	-- Specific Methods for Field Data Access --

	SetSweptFace(me : mutable; aSweptArea : mutable FaceSurface from StepShape) is virtual;
	SweptFace (me) returns mutable FaceSurface from StepShape is virtual;

    	
fields
    	sweptArea :  FaceSurface from StepShape;
	    	
end SweptFaceSolid;
