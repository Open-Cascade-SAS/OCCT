-- Created on: 2000-10-23
-- Created by: Pavel TELKOV
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



package XDEDRAW 

    ---Purpose: Provides DRAW commands for work with DECAF data structures

uses
    Draw

is

    class Shapes;
    	---Purpose: Provides functions for work with shapes and assemblies

    class Colors;
    	---Purpose: Provides functions for work with colors

    class Layers;
    	---Purpose: Provides functions for work with layers

    class Props;
    	---Purpose: Provides functions for work with geometric properties  
	
    class Common; 
    	---Purpose: Provides common commands for work XDE

    Init (di: in out Interpretor from Draw);
    	---Purpose: Initializes all the functions

    Factory (theDI : out Interpretor from Draw);
    ---Purpose: Loads all Draw commands of  TKXDEDRAW. Used for plugin.

end XDEDRAW;
