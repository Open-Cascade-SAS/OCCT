-- Created on: 2014-11-13
-- Created by: Maxim YAKUNIN
-- Copyright (c) 2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class FixSmallSolid from ShapeFix inherits Root from ShapeFix

	---Purpose: Fixing solids with small size

uses
    Shape   from TopoDS,
    ReShape from ShapeBuild
    
is
    Create returns FixSmallSolid;
    ---Purpose: Construct

    SetFixMode (me: mutable; theMode: Integer);
    ---Purpose: Set working mode for operator:
    -- - theMode = 0 use both WidthFactorThreshold and VolumeThreshold parameters
    -- - theMode = 1 use only WidthFactorThreshold parameter
    -- - theMode = 2 use only VolumeThreshold parameter
    
    SetVolumeThreshold (me: mutable; theThreshold: Real = -1.0);
    ---Purpose: Set or clear volume threshold for small solids

    SetWidthFactorThreshold (me: mutable; theThreshold: Real = -1.0);
    ---Purpose: Set or clear width factor threshold for small solids

    Remove(me; theShape: Shape from TopoDS; theContext: ReShape from ShapeBuild)
    returns Shape from TopoDS;
    ---Purpose: Remove small solids from the given shape
    
    Merge (me; theShape: Shape from TopoDS; theContext: ReShape from ShapeBuild)
    returns Shape from TopoDS;
    ---Purpose: Merge small solids in the given shape to adjacent non-small ones

    IsThresholdsSet (me) returns Boolean is private;

    IsSmall (me; theSolid: Shape from TopoDS) returns Boolean is private;

    IsUsedWidthFactorThreshold (me) returns Boolean is private;

    IsUsedVolumeThreshold (me) returns Boolean is private;

fields

    myFixMode              : Integer;
    myVolumeThreshold      : Real;
    myWidthFactorThreshold : Real;

end FixSmallSolid;
