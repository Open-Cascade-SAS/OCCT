-- Created on: 1994-05-31
-- Created by: Christian CAILLET
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class DispPerSingleView  from IGESSelect  inherits Dispatch

    ---Purpose : This type of dispatch defines sets of entities attached to
    --           distinct single views. This information appears in the
    --           Directory Part. Drawings are taken into account too,
    --           because of their frames (proper lists of annotations)
    --           
    --           Remaining data concern entities not attached to a single view.


uses AsciiString from TCollection, EntityIterator, Graph, SubPartsIterator,
     ViewSorter

is

    Create returns mutable DispPerSingleView;
    ---Purpose : Creates a DispPerSingleView

    Label (me) returns AsciiString from TCollection;
    ---Purpose : Returns as Label, "One File per single View or Drawing Frame"

    	    -- --    Evaluation    -- --

    Packets (me; G : Graph; packs : in out SubPartsIterator);
    ---Purpose : Computes the list of produced Packets. Packets are computed
    --           by a ViewSorter (SortSingleViews with also frames).

    CanHaveRemainder (me) returns Boolean  is redefined;
    ---Purpose : Returns True, because of entities attached to no view.

    Remainder (me; G : Graph) returns EntityIterator  is redefined;
    ---Purpose : Returns Remainder which is a set of Entities.
    --           It is supposed to be called once Packets has been called.

fields

    thesorter : ViewSorter;

end DispPerSingleView;
