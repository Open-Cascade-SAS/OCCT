-- Created on: 2008-12-10
-- Created by: Pavel TELKOV
-- Copyright (c) 2008-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class DimTol from PXCAFDoc inherits  Attribute from PDF

	---Purpose: 
uses
    Integer       from Standard,
    HAsciiString  from PCollection,
    HArray1OfReal from PColStd
is
    Create returns mutable DimTol from PXCAFDoc;

    Create (theKind : Integer from Standard;
    	    theVal  : HArray1OfReal from PColStd;
    	    theName : HAsciiString from PCollection;
    	    theDescr: HAsciiString from PCollection)
    returns mutable DimTol from PXCAFDoc;
    
    GetKind (me) returns Integer from Standard;

    GetVal (me) returns HArray1OfReal from PColStd;

    GetName (me) returns HAsciiString from PCollection;

    GetDescription (me) returns HAsciiString from PCollection;

    Set (me : mutable; theKind : Integer from Standard;
    	    	       theVal  : HArray1OfReal from PColStd;
    	    	       theName : HAsciiString from PCollection;
    	    	       theDescr: HAsciiString from PCollection);
    
fields

    myKind : Integer from Standard;
    myVal  : HArray1OfReal from PColStd;
    myName : HAsciiString from PCollection;
    myDescr: HAsciiString from PCollection;

end DimTol from PXCAFDoc;
