-- Created on: 1992-06-22
-- Created by: Gilles DEBARBOUILLE
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Quantity from Units 

inherits

    TShared from MMgt 


	---Purpose: This  class stores  in its  field all the possible
	--          units of all the unit systems for a given physical
	--          quantity. Each unit's  value  is  expressed in the
	--          S.I. unit system.

uses

    UnitsSequence from Units,
    Dimensions    from Units,
    HAsciiString  from TCollection,
    AsciiString   from TCollection

is

    Create(aname          : CString ;
           adimensions    : Dimensions    from Units ;
           aunitssequence : UnitsSequence from Units)
    
    ---Level: Internal 
    
    ---C++: inline
    
    ---Purpose: Creates  a new Quantity  object with <aname> which  is
    --          the name of the physical quantity, <adimensions> which
    --          is the physical dimensions, and <aunitssequence> which
    --          describes all the units known for this quantity.
    
    returns mutable Quantity from Units;
    
    Name(me) returns AsciiString from TCollection
    
    ---Level: Internal 
    
    ---C++: inline
    
    ---Purpose: Returns in a AsciiString from TCollection the name of the quantity.
    
    is static;
    
    Dimensions(me) returns any Dimensions from Units
    
    ---Level: Internal 
    
    ---C++: inline
    
    ---Purpose: Returns the physical dimensions of the quantity.
    
    is static;
    
    Sequence(me) returns any UnitsSequence from Units
    
    ---Level: Internal 
    
    ---C++: inline
    
    ---Purpose: Returns <theunitssequence>, which  is the  sequence of
    --          all the units stored for this physical quantity.
    
    is static;
    
    IsEqual(me ; astring : CString) returns Boolean
    
    ---Level: Internal 
    
--    ---C++: alias "friend Standard_EXPORT Standard_Boolean operator ==(const Handle(Units_Quantity)&,const Standard_CString);"
    
    ---Purpose: Returns True if the name of the Quantity <me> is equal 
    --          to <astring>, False otherwise.
    
    is static;
    
    Dump(me ; ashift , alevel : Integer)
    
    ---Level: Internal 
    
    ---Purpose: Useful for debugging.
    
    is static;

fields

    thename          : HAsciiString  from TCollection;
    thedimensions    : Dimensions    from Units;
    theunitssequence : UnitsSequence from Units;

end Quantity;
