-- Created on: 1999-01-14
-- Created by: Xuan PHAM PHU
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class face from TopOpeBRepTool

uses
    Wire from TopoDS,
    Face from TopoDS
is
    Create returns face from TopOpeBRepTool;
    Init (me : in out; W : Wire from TopoDS; Fref : Face from TopoDS) 
    returns Boolean;
    -- Builds face f for <myW> on <Fref>, 
    -- updates <myfinite> to true if f is finite,
    -- <myFfinite> is finite.
    -- returns false if the compute fails
    W(me) returns Wire from TopoDS;
    ---C++: return const &
    
    IsDone(me)  returns Boolean;    
    
    Finite(me)  returns Boolean;    
    Ffinite(me) returns Face from TopoDS; 
    ---C++: return const &   
    RealF(me)   returns Face from TopoDS;
    -- Raises if !IsDone
    
fields
    myW       : Wire from TopoDS;
    myfinite  : Boolean;
    myFfinite : Face from TopoDS;
    
end face;
