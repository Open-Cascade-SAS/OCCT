-- Created by: DAUTRY Philippe
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

--      	-------------------

---Version:	0.0
--Version	Date		Purpose
--		0.0	Sep  8 1998	Creation

class ClosureTool from TDF

	---Purpose: This class provides services to build the closure
	--          of an information set.
	--          
	--          You can set closure options by using IDFilter
	--          (to select or exclude specific attribute IDs) and
	--          CopyOption objects and by giving to Closure
	--          method.
	--          


uses

    Boolean             from Standard,
    Label               from TDF,
    Attribute           from TDF,
    DataSet             from TDF,
    RelocationTable     from TDF,
    AttributeMap        from TDF,
    LabelMap            from TDF,
    IDFilter            from TDF,
    ClosureMode         from TDF

-- raises

is

    Closure(myclass;
    	aDataSet : mutable DataSet from TDF);
	---Purpose: Builds the transitive closure of label and
	--          attribute sets into <aDataSet>.

    Closure(myclass;
    	aDataSet : mutable DataSet from TDF;
    	aFilter  : IDFilter from TDF;
    	aMode    : ClosureMode from TDF);
	---Purpose: Builds the transitive closure of label and
	--          attribute sets into <aDataSet>. Uses <aFilter> to
	--          determine if an attribute has to be taken in
	--          account or not. Uses <aMode> for various way of
	--          closing.


    -- ----------------------------------------------------------------------
    -- 
    -- Private methods
    -- 
    -- ----------------------------------------------------------------------

    Closure(myclass;
    	    aLabel   : Label        from TDF;
	    aLabMap  : in out LabelMap     from TDF;
	    anAttMap : in out AttributeMap from TDF;
    	    aFilter  : IDFilter     from TDF;
    	    aMode    : ClosureMode  from TDF);
	---Purpose: Builds the transitive closure of <aLabel>.


    LabelAttributes(myclass;
    	    	    aLabel   : Label        from TDF;
		    aLabMap  : in out LabelMap     from TDF;
		    anAttMap : in out AttributeMap from TDF;
    	    	    aFilter  : IDFilter     from TDF;
    	    	    aMode    : ClosureMode  from TDF)
    	is private;
	---Purpose: Adds label attributes and dependences.


end ClosureTool;
