-- File:        ShapeRepresentation.cdl
-- Created:     Mon Dec  4 12:02:31 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWShapeRepresentation from RWStepShape

	---Purpose : Read & Write Module for ShapeRepresentation

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     ShapeRepresentation from StepShape,
     EntityIterator from Interface

is

	Create returns RWShapeRepresentation;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable ShapeRepresentation from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : ShapeRepresentation from StepShape);

	Share(me; ent : ShapeRepresentation from StepShape; iter : in out EntityIterator);

end RWShapeRepresentation;
