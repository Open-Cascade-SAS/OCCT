-- File:        PointStyle.cdl
-- Created:     Fri Dec  1 11:11:25 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class PointStyle from StepVisual 

inherits TShared from MMgt

uses

	HAsciiString from TCollection, 
	MarkerSelect from StepVisual, 
	SizeSelect from StepBasic, 
	Colour from StepVisual
is

	Create returns mutable PointStyle;
	---Purpose: Returns a PointStyle

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aMarker : MarkerSelect from StepVisual;
	      aMarkerSize : SizeSelect from StepBasic;
	      aMarkerColour : mutable Colour from StepVisual) is virtual;

	-- Specific Methods for Field Data Access --

	SetName(me : mutable; aName : mutable HAsciiString);
	Name (me) returns mutable HAsciiString;
	SetMarker(me : mutable; aMarker : MarkerSelect);
	Marker (me) returns MarkerSelect;
	SetMarkerSize(me : mutable; aMarkerSize : SizeSelect);
	MarkerSize (me) returns SizeSelect;
	SetMarkerColour(me : mutable; aMarkerColour : mutable Colour);
	MarkerColour (me) returns mutable Colour;

fields

	name : HAsciiString from TCollection;
	marker : MarkerSelect from StepVisual; -- a SelectType
	markerSize : SizeSelect from StepBasic; -- a SelectType
	markerColour : Colour from StepVisual;

end PointStyle;
