-- Created on: 1994-08-26
-- Created by: Frederic MAUPAS
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MakeAxis2Placement2d from GeomToStep inherits Root from GeomToStep

    ---Purpose: This class implements the mapping between classes 
    --          Axis2Placement from Geom and Ax2, Ax22d from gp, and the class
    --          Axis2Placement2d from StepGeom which describes an
    --          axis2_placement_2d from Prostep. 
   
uses Ax2              from gp,
     Ax22d            from gp,
     Axis2Placement   from Geom,
     Axis2Placement2d from StepGeom
     
raises NotDone from StdFail
     
is 

Create ( A : Ax2 from gp ) returns MakeAxis2Placement2d;

Create ( A : Ax22d from gp ) returns MakeAxis2Placement2d;

--Create ( A : Axis2Placement from Geom ) returns MakeAxis2Placement2d;

Value (me) returns Axis2Placement2d from StepGeom
    raises NotDone
    is static;
    ---C++: return const&

fields

    theAxis2Placement2d : Axis2Placement2d from StepGeom;
    	-- TheOP solution from StepGeom
    	
end MakeAxis2Placement2d;


