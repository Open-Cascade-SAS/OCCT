-- Created on: 1991-02-22
-- Created by: Jean Claude Vauthier
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package CPnts 

        --- Purpose :  
        --  This package  contains   the definition  of  the geometric
        --  algorithms   used to  compute  characteristic  points   on
        --  parametrized curves in 3d or 2d space. 
        --  This package defines the external geometric entities, with
        --  their requirements, used in the algorithms.

uses math, gp, StdFail, Adaptor3d  ,  Adaptor2d

is


   imported RealFunction;

   private class MyGaussFunction;

   private class MyRootFunction;

   class  AbscissaPoint;

   class UniformDeflection;

end CPnts;








