-- Created by: Peter KURNEV
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class BOP from BOPAlgo  
    inherits Builder from BOPAlgo
---Purpose: 

uses
    Shape from TopoDS,  
    BaseAllocator from BOPCol,  
    ListOfShape from BOPCol, 
    ListOfShape from TopTools, 
    MapOfShape  from BOPCol,  
    IndexedDataMapOfShapeListOfShape from BOPCol,
    Operation from BOPAlgo, 
    PaveFiller from BOPAlgo 

--raises

is
    Create 
    ---Purpose:  Empty constructor     
    returns BOP from BOPAlgo;  
    ---C++: alias "Standard_EXPORT virtual ~BOPAlgo_BOP();"  
      
    Create (theAllocator: BaseAllocator from BOPCol)
    returns BOP from BOPAlgo; 
	 
    Clear(me:out) 
    is redefined; 
    ---Purpose:  Clears internal fields and arguments   
     
    AddArgument (me:out;  
        theShape: Shape from TopoDS) 
    ---Purpose:  Adds Object argument of the operation     
     is redefined;
	 
    AddTool (me:out;  
        theShape: Shape from TopoDS) 
    ---Purpose:  Adds Tool argument of the operation    	     
    is virtual; 
	 
    Object(me) 
    returns Shape from TopoDS; 
    ---C++: return const &   

    Tool(me) 
    returns Shape from TopoDS; 
    ---C++: return const &   

    SetOperation(me:out;  
        theOperation: Operation from BOPAlgo); 
	 
    Operation(me) 
    returns Operation from BOPAlgo;  
    --
    --  protected methods 
    -- 
    CheckData(me:out) 
    is redefined protected; 

    Prepare(me:out)  
    is redefined protected; 
    ---Purpose:  Provides preparing actions 

    PerformInternal(me:out; 
        thePF:PaveFiller from BOPAlgo) 
    is redefined protected;   
    ---Purpose:  Performs calculations using prepared Filler 
    --           object theDSF          	 
      
    BuildShape(me:out) 
    is protected; 
 
    BuildRC(me:out) 
    is protected; 
 
    BuildSolid(me:out) 
    is protected; 
	 
    BuildSection(me:out) 
    is protected;  
 
    IsBoundSplits(me:out; 
        theS:Shape from TopoDS; 
        theMEF:out IndexedDataMapOfShapeListOfShape from BOPCol)  
    returns Boolean from Standard
    is protected;

    Generated (me:out;  
        theS : Shape from TopoDS)
    ---Purpose: Returns the  list of shapes generated from the
    --          shape theS. 
    returns ListOfShape from TopTools
    is redefined;
    ---C++: return const & 

fields 
    myNbArgs    : Integer from Standard    is protected;
    myOperation : Operation from BOPAlgo   is protected; 
    myArgs      : Shape from TopoDS[2]     is protected;  
    myDims      : Integer from Standard[2] is protected;  
    -- 
    myRC        : Shape from TopoDS        is protected; 
    myTools     : ListOfShape from BOPCol  is protected; 
    myMapTools  : MapOfShape  from BOPCol  is protected;  
    
end BOP;
