-- Created on: 2000-04-18
-- Created by: Andrey BETENEV
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0

class DimensionalCharacteristic from StepShape
inherits SelectType from StepData

    ---Purpose: Representation of STEP SELECT type DimensionalCharacteristic

uses
    DimensionalLocation from StepShape,
    DimensionalSize from StepShape

is
    Create returns DimensionalCharacteristic from StepShape;
	---Purpose: Empty constructor

    CaseNum (me; ent: Transient) returns Integer;
	---Purpose: Recognizes a kind of DimensionalCharacteristic select type
	--          1 -> DimensionalLocation from StepShape
	--          2 -> DimensionalSize from StepShape
	--          0 else

    DimensionalLocation (me) returns DimensionalLocation from StepShape;
	---Purpose: Returns Value as DimensionalLocation (or Null if another type)

    DimensionalSize (me) returns DimensionalSize from StepShape;
	---Purpose: Returns Value as DimensionalSize (or Null if another type)

end DimensionalCharacteristic;
