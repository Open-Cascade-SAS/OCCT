-- Created on: 1991-03-06
-- Created by: Denis Pascal
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



generic class VertexIterator from GraphTools (Graph  as any;
		    		               Vertex as any)
				  
--template class VertexIterator from GraphTools (Graph  as any,
--                                                 Vertex as any)
				  
    ---Purpose: Template class which  defines Signature of an iterator
    --          to visit each adjacent vertex  of a  given one  in the
    --          underlying graph.


raises NoMoreObject from Standard,
       NoSuchObject from Standard

is

    Create (G : Graph; V : Vertex) returns VertexIterator;

    More (me) returns Boolean;
	---Purpose: Returns TRUE if there are other vertices.
       ---Level: Public

    Next(me : in out)
    	--- Purpose : Set the iterator to the next Vertex.
       ---Level: Public
    raises NoMoreObject from Standard;

    Value(me) returns Vertex
	--- Purpose: Returns the vertex value for the current position
	--           of the iterator.
       ---Level: Public
    raises NoSuchObject from Standard;

end VertexIterator;



















