-- File:	Interface_IntList.cdl
-- Created:	Fri May 12 17:48:33 1995
-- Author:	Christian CAILLET
--		<cky@anion>
---Copyright:	 Matra Datavision 1995


class IntList  from Interface

    ---Purpose : This class detains the data which describe a Graph. A Graph
    --           has two lists, one for shared refs, one for sharing refs
    --           (the reverses). Each list comprises, for each Entity of the
    --           Model of the Graph, a list of Entities (shared or sharing).
    --           In fact, entities are identified by their numbers in the Model
    --           or Graph : this gives better performances.
    --           
    --           A simple way to implement this is to instantiate a HArray1
    --           with a HSequenceOfInteger : each Entity Number designates a
    --           value, which is a Sequence (if it is null, it is considered as
    --           empty : this is a little optimisation).
    --           
    --           This class gives a more efficient way to implement this.
    --           It has two lists (two arrays of integers), one to describe
    --           list (empty, one value given immediately, or negated index in
    --           the second list), one to store refs (pointed from the first
    --           list). This is much more efficient than a list of sequences,
    --           in terms of speed (especially for read) and of memory
    --           
    --           An IntList can also be set to access data for a given entity
    --           number, it then acts as a single sequence
    --           
    --           Remark that if an IntList is created from another one, it can
    --           be read, but if it is created without copying, it may not be
    --           edited

uses HArray1OfInteger

is
    Create returns IntList;
    ---Purpose :Creates empty IntList.
    
   
    
    Create (nbe : Integer) returns IntList;
    ---Purpose : Creates an IntList for <nbe> entities

    Create (other : IntList; copied : Boolean) returns IntList;
    ---Purpose : Creates an IntList from another one.
    --           if <copied> is True, copies data
    --           else, data are not copied, only the header object is
    Initialize(me : in out;nbe : Integer);
    ---Purpose :Initialize IntList by number of entities.
    Internals (me; nbrefs : out Integer; ents, refs : out mutable HArray1OfInteger);
    ---Purpose : Returns internal values, used for copying

    NbEntities (me) returns Integer;
    ---Purpose : Returns count of entities to be aknowledged

    SetNbEntities (me : in out; nbe : Integer);
    ---Purpose : Changes the count of entities (ignored if decreased)

    SetNumber (me : in out; number : Integer);
    ---Purpose : Sets an entity number as current (for read and fill)

    Number (me) returns Integer;
    ---Purpose : Returns the current entity number

    List (me; number : Integer; copied : Boolean = Standard_False) returns IntList;
    ---Purpose : Returns an IntList, identical to <me> but set to a specified
    --           entity Number
    --           By default, not copied (in order to be read)
    --           Specified <copied> to produce another list and edit it

    SetRedefined (me : in out; mode : Boolean);
    ---Purpose : Sets current entity list to be redefined or not
    --           This is used in a Graph for redefinition list : it can be
    --           disable (no redefinition, i.e. list is cleared), or enabled
    --           (starts as empty). The original list has not to be "redefined"

    Reservate (me : in out; count : Integer);
    ---Purpose : Makes a reservation for <count> references to be later
    --           attached to the current entity. If required, it increases
    --           the size of array used to store refs. Remark that if count is
    --           less than two, it does nothing (because immediate storing)

    Add (me : in out; ref : Integer);
    ---Purpose : Adds a reference (as an integer value, an entity number) to
    --           the current entity number. Zero is ignored

    Length (me) returns Integer;
    ---Purpose : Returns the count of refs attached to current entity number

    IsRedefined (me; num : Integer = 0) returns Boolean;
    ---Purpose : Returns True if the list for a number (default is taken as
    --           current) is "redefined"  (usefull for empty list)

    Value (me; num : Integer) returns Integer;
    ---Purpose : Returns a reference number in the list for current number,
    --           according to its rank

    Remove (me : in out; num : Integer) returns Boolean;
    ---Purpose : Removes an item in the list for current number, given its rank
    --           Returns True if done, False else

    Clear (me : in out);
    ---Purpose : Clears all data, hence each entity number has an empty list

    AdjustSize (me : in out; margin : Integer = 0);
    ---Purpose : Resizes lists to exact sizes. For list of refs, a positive
    --           margin can be added.

fields

    thenbe   : Integer;
    thenbr   : Integer;
    thenum   : Integer;  -- for current entity number :
    thecount : Integer;
    therank  : Integer;
    theents  : HArray1OfInteger;
    therefs  : HArray1OfInteger;

end IntList;
