-- Created on: 1997-07-28
-- Created by: Pierre CHALAMET
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

deferred class TextureRoot from Graphic3d

inherits TShared from MMgt

    ---Purpose: This is the texture root class enable the dialog with the GraphicDriver 
    -- allows the loading of texture.

uses

    CInitTexture     from Graphic3d,
    GraphicDriver    from Graphic3d,
    StructureManager from Graphic3d,
    TypeOfTexture    from Graphic3d,
    PixMap           from Image,
    Path             from OSD,
    HArray1OfReal    from TColStd

is

    Initialize (theSM       :  StructureManager from Graphic3d;
                thePath     :  CString from Standard;
                theFileName :  CString from Standard;
                theType     :  TypeOfTexture from Graphic3d);
    ---Purpose: Creates a texture from a file	       
    --  Warning: Note that if <FileName> is NULL the texture must be realized
    -- using LoadTexture(image) method.

    Destroy (me);
    ---C++ : alias ~

    --
    -- public methods
    --

    IsDone (me) returns Boolean from Standard;
    ---Level: public
    ---Purpose: Checks if a texture class is valid or not
    -- returns true if the construction of the class is correct

    IsValid (me) returns Boolean from Standard;
    ---Level: public
    ---Purpose: Checks if a texture class is valid or not
    -- returns true if the construction of the class is correct

    Path (me) returns Path from OSD;
    ---Level: public
    ---Purpose:
    -- Returns the full path of the defined texture.
    ---C++: return const &

    Type (me) returns TypeOfTexture from Graphic3d;
    ---Level: public
    ---Purpose:
    -- Returns the texture type.

    LoadTexture (me : mutable; theImage : PixMap from Image) returns Boolean from Standard;
    ---Level: advanced
    ---Purpose:
    -- Updates the current texture from a requested image.

    TextureId (me) returns Integer from Standard;
    ---Level: advanced
    ---Purpose:
    -- returns the Texture ID which references the
    -- texture to use for drawing. Used by the graphic driver.

    GetTexUpperBounds(me) returns HArray1OfReal from TColStd;
    ---Level: advanced
    ---Purpose:
    ---Gets upper bounds of texture coordinates. This is used when sizes
    ---of texture are not equal to the powers of two

    --
    -- private methods
    --

    Update (me) is protected;

fields

    myGraphicDriver  : GraphicDriver from Graphic3d;
    myTexId          : Integer from Standard;
    MyCInitTexture   : CInitTexture from Graphic3d is protected;
    myPath           : Path from OSD;
    myType           : TypeOfTexture from Graphic3d;
    myTexUpperBounds : HArray1OfReal from TColStd;

end TextureRoot;
