-- Created on: 1992-11-18
-- Created by: Christian CAILLET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SelectErrorEntities  from IFSelect  inherits SelectExtract

    ---Purpose : A SelectErrorEntities sorts the Entities which are qualified
    --           as "Error" (their Type has not been recognized) during reading
    --           a File. This does not concern Entities which are syntactically
    --           correct, but with incorrect data (for integrity constraints).

uses AsciiString from TCollection, InterfaceModel

is

    Create returns SelectErrorEntities;
    ---Purpose : Creates a SelectErrorEntities

    Sort (me; rank : Integer; ent : Transient; model : InterfaceModel)
    	returns Boolean;
    ---Purpose : Returns True for an Entity which is qualified as "Error", i.e.
    --           if <model> explicitly knows <ent> (through its Number) as
    --           Erroneous


    ExtractLabel (me) returns AsciiString from TCollection;
    ---Purpose : Returns a text defining the criterium : "Error Entities"

end SelectErrorEntities;
