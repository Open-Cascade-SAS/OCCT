--
-- File:	Graphic3d_VertexC.cdl
-- Created:	Jeudi 22 Aout 1991
-- Author:	NW,JPB,CAL
--
---Copyright:	MatraDatavision 1991,1992,1993
--

class VertexC from Graphic3d inherits Vertex from Graphic3d

	---Version:

	---Purpose: This class allows the creation and update of a point
	--	    with a colour value.

	---Keywords: Vertex, Color, Coordinate, Point

	---Warning:
	---References:

uses

	Color	from Quantity
    	---Purpose: Returns the color of this point.
is

	Create
		returns VertexC from Graphic3d;
    	---Purpose: Constructs an empty point
        
	Create ( AX, AY ,AZ	: Real from Standard;
		 AColor		: Color from Quantity )
		returns VertexC from Graphic3d;
	---Level: Public
	---Purpose: Creates a point with coordinates <AX>, <AY>, <AZ> and
	--	    with colour <AColor>.

	Create ( APoint	: Vertex from Graphic3d;
		 AColor	: Color from Quantity )
		returns VertexC from Graphic3d;
	---Level: Public
	---Purpose: Creates a point situated in <APoint> and
	--	    for which the colour is <AColor>.

	---------------------------------------------------
	-- Category: Methods to modify the class definition
	---------------------------------------------------

	SetColor ( me		: in out;
		   ColorNew	: Color from Quantity )
		is static;
	---Level: Public
	---Purpose: Modifies the colour of the point <me>.
	---Category: Methods to modify the class definition

	----------------------------
	-- Category: Inquire methods
	----------------------------

	Color ( me )
		returns Color from Quantity
		is static;
	---Level: Public
	---Purpose: Returns the colour of the point <me>.
	---Category: Inquire methods

--

fields

--
-- Class	:	Graphic3d_VertexC
--
-- Purpose	:	Declaration of variables specific to points
--
-- Reminder	:	a point is defined by its coordinates and its colour
--

	-- the colour of a point
	MyColor		:	Color from Quantity;

end VertexC;
