-- File:	RWStepShape_RWExtrudedFaceSolid.cdl
-- Created:	Mon Mar 15 15:13:10 1999
-- Author:	data exchange team
--		<det@androx.nnov.matra-dtv.fr>
---Copyright:	 Matra Datavision 1999


class RWExtrudedFaceSolid from RWStepShape 

	---Purpose: Read & Write Module for ExtrudedFaceSolid

uses
     Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     ExtrudedFaceSolid from StepShape,
     EntityIterator from Interface

is
	Create returns RWExtrudedFaceSolid;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable ExtrudedFaceSolid from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : ExtrudedFaceSolid from StepShape);

	Share(me; ent : ExtrudedFaceSolid from StepShape; iter : in out EntityIterator);


end RWExtrudedFaceSolid;
