-- Created on: 1994-09-02
-- Created by: Yves FRICAUD
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



generic class NumericCurInf from LProp (Curve as any;
    	    	    	    	        Vec   as any; -- as Vec or Vec2d
		     	                Pnt   as any; -- as Pnt or Pnt2d
		   	                Dir   as any; -- as Dir or Dir2d Vec  
    	    	    	    	    	Tool  as any) -- as Tool(Curve, Pnt, Vec) 
					
	---Purpose: Computes the locals extremas of curvature and the 
    	--          inflections of a bounded curve in 2d. 

uses
    CurAndInf from LProp
    
private class FCurExt instantiates FuncCurExt from LProp (Curve,Vec,Pnt,Dir,Tool); 
private class FCurNul instantiates FuncCurNul from LProp (Curve,Vec,Pnt,Dir,Tool);

is
    Create;
    
    PerformCurExt (me : in out; C : Curve; Result : in out CurAndInf) 
    	---Purpose: Computes the locals extremas of curvature.
    is static;
    
    PerformInf    (me : in out; C : Curve; Result : in out CurAndInf)
       	---Purpose: Computes the inflections.
    is static;
    
    PerformCurExt (me     : in out; 
    	           C      : Curve ; 
                   UMin   : Real;
    	    	   UMax   : Real;
    	    	   Result : in out CurAndInf) 
    	---Purpose: Computes the locals extremas of curvature.
    	--          in the interval of parmeters [UMin,UMax].
    is static;
    
    PerformInf    (me     : in out;
        	   C      : Curve ; 
                   UMin   : Real;
    	    	   UMax   : Real;
    	    	   Result : in out CurAndInf)
       	---Purpose: Computes the inflections in the interval of 
       	--          parmeters [UMin,UMax].
    is static;
    
    IsDone (me) returns Boolean
	---Purpose: True if the solutions are found.
    is static;
    
fields
    isDone : Boolean from Standard;

end NumericCurInf;
