-- Created on: 1993-01-11
-- Created by: CKY / Contract Toubro-Larsen ( Arun MENON )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class LevelFunction from IGESAppli  inherits IGESEntity

        ---Purpose: defines LevelFunction, Type <406> Form <3>
        --          in package IGESAppli
        --          Used to transfer the meaning or intended use of a level
        --          in the sending system

uses

        HAsciiString from TCollection

is

        Create returns LevelFunction;

        -- Specific Methods pertaining to the class

        Init (me           : mutable;
              nbPropVal    : Integer;
              aCode        : Integer;
              aFuncDescrip : HAsciiString);
        ---Purpose : This method is used to set the fields of the class
        --           LevelFunction
        --       - nbPropVal    : Number of Properties, always = 2
        --       - aCode        : Function Description code
        --                        default = 0
        --       - aFuncDescrip : Function Description
        --                        default = null string

        NbPropertyValues (me) returns Integer;
        ---Purpose : is always 2

        FuncDescriptionCode (me) returns Integer;
        ---Purpose : returns the function description code . Default = 0

        FuncDescription (me) returns HAsciiString from TCollection;
        ---Purpose : returns the function description
        -- Default = null string

fields

--
-- Class    : IGESAppli_LevelFunction
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class LevelFunction.
--
-- Reminder : A LevelFunction instance is defined by :
--            -  Function Description code, default = 0
--            -  Function Description, default = null string

        theNbPropertyValues : Integer;
        theFuncDescripCode  : Integer;
        theFuncDescrip      : HAsciiString;

end LevelFunction;
