-- Created on: 1998-01-14
-- Created by: Philippe MANGIN
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DraftLaw from BRepFill  inherits  Edge3DLaw  from  BRepFill 

	---Purpose: Build Location Law, with a  Wire.

uses 
  LocationDraft  from  GeomFill, 
  Wire   from TopoDS

is    
  Create (Path   :  Wire  from  TopoDS; 
          Law    :  LocationDraft  from  GeomFill)   
  returns DraftLaw from BRepFill;   
   
  CleanLaw(me  :  mutable;  TolAngular  :  Real)  
    ---Purpose: To clean the little discontinuities.          
  is  static;    
    
end DraftLaw;



