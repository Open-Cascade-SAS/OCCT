-- Created on: 1999-10-29
-- Created by: Pavel DURANDIN
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class UndefinedTypeHandler from GeomTools inherits TShared from MMgt

	---Purpose: 

uses

    Curve   from Geom,
    Surface from Geom,
    Curve   from Geom2d,
    OStream,
    IStream

is

    Create returns mutable UndefinedTypeHandler from GeomTools;
    
    -- Curve
    
    PrintCurve(me; C  : Curve from Geom;
    	      	   OS : in out OStream;
		   compact : Boolean = Standard_False) is virtual;
    
    ReadCurve(me; ctype: Integer;
    	    	  IS   : in out IStream;
    	    	  C    : in out Curve from Geom)
    returns IStream is virtual;
    ---C++: return &
    
    --PCurve
    
    PrintCurve2d(me; C  : Curve from Geom2d;
    	    	     OS : in out OStream;
		     compact : Boolean = Standard_False) is virtual;
    
    ReadCurve2d(me; ctype: Integer;
    	    	    IS   : in out IStream;
    	    	    C    : in out Curve from Geom2d)
    returns IStream is virtual;
    ---C++: return &
    
    --Surface
    
    PrintSurface(me; S  : Surface from Geom;
    	    	     OS : in out OStream;
		     compact : Boolean = Standard_False) is virtual;
    
    ReadSurface(me; ctype: Integer;
    	    	    IS   : in out IStream;
    	    	    S    : in out Surface from Geom)
    returns IStream is virtual;
    ---C++: return &
    
end UndefinedTypeHandler;
