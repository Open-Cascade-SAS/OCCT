-- Created on: 1995-12-07
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class PointClassifier from TopOpeBRep

uses 

    State from TopAbs,
    Face from TopoDS,
    Pnt2d from gp,
    TopolTool from BRepTopAdaptor,
    HSurface from BRepAdaptor,
    DataMapOfTopolTool from TopOpeBRep    
    
is

    Create returns PointClassifier from TopOpeBRep;
    
    Init(me:in out) is static;
    
    Load(me:in out;F:Face from TopoDS) is static;

    Classify(me:in out;F:Face from TopoDS;P:Pnt2d from gp;Tol:Real)
    ---Purpose: compute position of point <P> regarding with the face <F>. 
    returns State from TopAbs is static;

    State(me) returns State from TopAbs is static;    

fields

    myTopolTool : TopolTool from BRepTopAdaptor;
    myHSurface : HSurface from BRepAdaptor;
    myTopolToolMap : DataMapOfTopolTool from TopOpeBRep;
    myState : State from TopAbs;
    
end PointClassifier from TopOpeBRep;
