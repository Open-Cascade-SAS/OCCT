-- Created on: 1997-02-12
-- Created by: Alexander BRIVIN
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class PerspectiveCamera from Vrml 

	---Purpose: specifies a PerspectiveCamera node of VRML specifying properties of cameras. 
    	--  A perspective camera defines a perspective projection from a viewpoint. The viewing
       	--  volume for a perspective camera is a truncated right pyramid. 
uses
 
     Vec         from gp, 
     SFRotation  from  Vrml
is
                                                    --  defaults  :
    Create  returns  PerspectiveCamera from Vrml;   --  myPosition(0 0 1) Camera looks along the negative Z-axis
 						    --  myOrientation(0 0 1 0)
						    --  myFocalDistance(5)
						    --  myHeightAngle(0.785398)
    Create  ( aPosition      :  Vec         from  gp; 
    	      aOrientation   :  SFRotation  from  Vrml; 
    	      aFocalDistance :  Real        from  Standard; 
    	      aHeightAngle   :  Real        from  Standard ) 
    	returns  PerspectiveCamera from Vrml; 

    SetPosition ( me : in out;  aPosition : Vec  from  gp );
    Position ( me  )  returns Vec  from  gp;

    SetOrientation ( me : in out;  aOrientation : SFRotation  from  Vrml );
    Orientation ( me )  returns SFRotation  from  Vrml;

    SetFocalDistance ( me : in out;  aFocalDistance : Real  from  Standard );
    FocalDistance ( me )  returns Real  from  Standard;

    SetAngle ( me : in out;  aHeightAngle : Real  from  Standard );
    Angle ( me )  returns  Real  from  Standard;

    Print  ( me;  anOStream: in out OStream from Standard) returns OStream from Standard;
    ---C++:  return  & 

fields
 
    myPosition      :  Vec         from  gp;       -- Location of viewpoint
    myOrientation   :  SFRotation  from  Vrml;     -- Orientation (rotation with respect to (0,0,-1) vector)     
    myFocalDistance :  Real        from  Standard; -- Distance from viewpoint to point of focus.
    myHeightAngle   :  Real        from  Standard; -- Angle (in radians) of field
    	    	    	    	    	    	   -- of  view, in  height  direction
end PerspectiveCamera;
