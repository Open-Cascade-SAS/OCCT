-- File:	TDataXtd_Shape.cdl
-- Created:	Mon Apr  6 18:16:04 2009
-- Author:	Sergey ZARITCHNY
--		<sergey.zaritchny@opencascade.com>
---Copyright:	Open CasCade SA 2009 

class Shape from TDataXtd inherits Attribute from TDF

	---Purpose: A Shape is associated in the framework with :
	--          a NamedShape attribute 


uses Attribute       from TDF,
     Label           from TDF,
     NamedShape      from TNaming,
     GUID            from Standard,
     DataSet         from TDF,
     RelocationTable from TDF,
     Shape           from TopoDS
is    


    ---Purpose: class methods
    --          =============
    
    Find (myclass; current : Label from TDF; S : in out Shape from TDataXtd)
    ---Purpose: try to retrieve a Shape attribute at <current> label
    --           or in  fathers  label of  <current>. Returns True  if
    --          found and set <S>.
    returns Boolean from Standard;
    
    New (myclass; label : Label from TDF)
    ---Purpose: Find, or create, a Shape attribute.  the Shape attribute
    --          is returned. Raises if <label> has attribute.
    returns Shape from TDataXtd;

    Set (myclass; label : Label from TDF; shape : Shape from TopoDS)
    ---Purpose: Create or update associated NamedShape attribute.  the
    --          Shape attribute is returned.
    returns Shape from TDataXtd;    

    Get (myclass; label : Label from TDF)
    ---Purpose:   the Shape from  associated NamedShape attribute
    --            is returned.
    returns Shape from TopoDS;
    
    GetID (myclass)   
    ---C++: return const &  
    returns GUID from Standard;

    ---Purpose: Shape methods
    --          ============

    Create
    returns mutable Shape from TDataXtd;

    
    ---Category: methodes de TDF_Attribute
    --           =========================
 
	
    ID (me)
    ---C++: return const & 
    returns GUID from Standard;

    Restore (me: mutable; with : Attribute from TDF);

    NewEmpty (me)
    returns mutable Attribute from TDF;

    Paste (me; into : mutable Attribute from TDF;
	       RT   : mutable RelocationTable from TDF);       

    References (me; DS : DataSet from TDF) is redefined;   

    Dump(me; anOS : in out OStream from Standard)
    returns OStream from Standard
     is redefined;
	---C++: return &

end Shape;

