-- File:	QAYasaki.cdl
-- Created:	Tue May 21 11:10:01 2002
-- Author:	QA Admin
--		<qa@russox>
---Copyright:	 Matra Datavision 2002

package QAYasaki
     uses Draw
is
    Commands(DI : in out Interpretor from Draw);
end;
