-- File:        SiUnitAndPlaneAngleUnit.cdl
-- Created:     Fri Dec  1 11:11:34 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class SiUnitAndPlaneAngleUnit from StepBasic inherits SiUnit from StepBasic 

	--- This classe is an implementation of EXPRESS
	--  ANDOR Subtype Declaration.
uses

    PlaneAngleUnit from StepBasic, 
    DimensionalExponents from StepBasic, 
    SiPrefix from StepBasic, 
    SiUnitName from StepBasic

is

    Create returns mutable SiUnitAndPlaneAngleUnit;
	---Purpose: Returns a SiUnitAndPlaneAngleUnit

    Init (me: mutable; aDimensions : mutable DimensionalExponents from StepBasic)
    is redefined;

    Init (me: mutable; hasAprefix : Boolean from Standard;
		       aPrefix : SiPrefix from StepBasic;
		       aName : SiUnitName from StepBasic) is redefined;

    -- Specific Methods for Field Data Access --

    SetPlaneAngleUnit(me: mutable; aPlaneAngleUnit: mutable PlaneAngleUnit);
    
    PlaneAngleUnit (me) returns mutable PlaneAngleUnit;

fields

    planeAngleUnit : PlaneAngleUnit from StepBasic;

end SiUnitAndPlaneAngleUnit;
