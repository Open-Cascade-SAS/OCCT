-- File:	Geom_Conic.cdl
-- Created:	Wed Mar 10 09:30:27 1993
-- Author:	JCV
--		<fid@phylox>
-- Copyright:	 Matra Datavision 1993


deferred class Conic from Geom inherits Curve from Geom

    	---Purpose : The abstract class Conic describes the common
    	-- behavior of conic curves in 3D space and, in
    	-- particular, their general characteristics. The Geom
    	-- package provides four concrete classes of conics:
    	-- Geom_Circle, Geom_Ellipse, Geom_Hyperbola and Geom_Parabola.
    	-- A conic is positioned in space with a right-handed
    	-- coordinate system (gp_Ax2 object), where:
    	-- - the origin is the center of the conic (or the apex in
    	--   the case of a parabola),
    	-- - the origin, "X Direction" and "Y Direction" define the
    	--   plane of the conic.
    	-- This coordinate system is the local coordinate
    	-- system of the conic.
    	-- The "main Direction" of this coordinate system is the
    	-- vector normal to the plane of the conic. The axis, of
    	-- which the origin and unit vector are respectively the
    	-- origin and "main Direction" of the local coordinate
    	-- system, is termed the "Axis" or "main Axis" of the conic.
    	-- The "main Direction" of the local coordinate system
    	-- gives an explicit orientation to the conic, determining
    	-- the direction in which the parameter increases along
    	-- the conic. The "X Axis" of the local coordinate system
    	-- also defines the origin of the parameter of the conic.
      

uses  Ax1   from gp, 
      Ax2   from gp, 
      Pnt   from gp, 
      Vec   from gp,
      Shape from GeomAbs


raises ConstructionError from Standard,
       RangeError        from Standard,
       DomainError       from Standard

is

  SetAxis (me : mutable; A1 : Ax1)
    	---Purpose : Changes the orientation of the conic's plane. The normal
    	--  axis to the plane is A1. The XAxis and the YAxis are recomputed.
     raises ConstructionError;
        ---Purpose :
        --  raised if the A1 is parallel to the XAxis of the conic.


  SetLocation (me : mutable; P : Pnt);
        ---Purpose : changes the location point of the conic.


  SetPosition (me : mutable; A2 : Ax2);
        ---Purpose : changes the local coordinate system of the conic.


  Axis (me)  returns Ax1;
        ---Purpose : Returns the "main Axis" of this conic. This axis is
    	-- normal to the plane of the conic.
     

  Eccentricity (me)  returns Real
        ---Purpose :
        --  Returns the eccentricity value of the conic e.
        --  e = 0 for a circle
        --  0 < e < 1 for an ellipse  (e = 0 if MajorRadius = MinorRadius)
        --  e > 1 for a hyperbola
        --  e = 1 for a parabola
      	--  Exceptions
    	-- Standard_DomainError in the case of a hyperbola if
    	-- its major radius is null.
     raises DomainError
     is deferred;


  Location (me)  returns Pnt;
        ---Purpose :
        --  Returns the location point of the conic.
        --  For the circle, the ellipse and the hyperbola it is the center of
        --  the conic. For the parabola it is the Apex of the parabola.


  Position (me)   returns Ax2;
        ---Purpose :
	--  Returns the local coordinates system of the conic.
        --  The main direction of the Axis2Placement is normal to the
        --  plane of the conic. The X direction of the Axis2placement
        --  is in the plane of the conic and corresponds to the origin 
        --  for the conic's parametric value u.
    	---C++: return const&


  XAxis (me)  returns Ax1;
        ---Purpose :
        -- Returns the XAxis of the conic.
        -- This axis defines the origin of parametrization of the conic.
        -- This axis is perpendicular to the Axis of the conic.
        -- This axis and the Yaxis define the plane of the conic.


  YAxis (me)  returns Ax1;
        ---Purpose :
        --  Returns the YAxis of the conic.
        --  The YAxis is perpendicular to the Xaxis.
        --  This axis and the Xaxis define the plane of the conic.
	  

  Reverse (me : mutable);
	---Purpose :
	--  Reverses the direction of parameterization of <me>.
        --  The local coordinate system of the conic is modified.


  ReversedParameter(me; U : Real) returns Real
	---Purpose: Returns the  parameter on the  reversed  curve for
	--          the point of parameter U on <me>.
	--          
  is deferred;


  Continuity (me)   returns Shape from GeomAbs;
        ---Purpose : The continuity of the conic is Cn.
        
  IsCN (me; N : Integer) returns Boolean
        ---Purpose : Returns True. 
     raises RangeError;
        ---Purpose : Raised if N < 0.

fields

  pos : Ax2 is protected;

end;

