-- Created on: 1993-04-06
-- Created by: Philippe DAUTRY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class TrimmedCurve from PGeom2d inherits BoundedCurve from PGeom2d

        ---Purpose :
        --  Defines a portion of a curve limited by two values of 
        --  parameters inside the parametric domain of the curve.
        --  
	---See Also : TrimmedCurve from Geom2d.


uses Curve from PGeom2d

is


  Create returns mutable TrimmedCurve from PGeom2d;
	---Purpose: Creates a TrimmedCurve with default values.
	---Level: Advanced 


  Create (
    	aBasisCurve: Curve from PGeom2d;
    	aFirstU, aLastU: Real from Standard)
     returns mutable TrimmedCurve from PGeom2d;
        ---Purpose : Creates a TrimmedCurve with these field values.
	---Level: Advanced 


  FirstU(me : mutable; aFirstU: Real from Standard);
        ---Purpose : Set the value of the field firstU with <aFirstU>.
	---Level: Advanced 


  FirstU(me) returns Real from Standard;
        ---Purpose : Returns the value of the field firstU.
	---Level: Advanced 


  LastU(me : mutable; aLastU: Real from Standard);
        ---Purpose : Set the value of the field lastU with <aLastU>.
	---Level: Advanced 


  LastU(me) returns Real from Standard;
        ---Purpose : Returns the value of the field lastU.
	---Level: Advanced 


  BasisCurve (me: mutable; aBasisCurve: Curve from PGeom2d);
        ---Purpose : Set the value of the field basisCurve with <aBasisCurve>.
        --  This curve can be a trimmed curve.
	---Level: Advanced 


  BasisCurve (me) returns Curve from PGeom2d;
        ---Purpose : Returns the value of the field basisCurve. 
        --  This curve can be a trimmed curve.
	---Level: Advanced 


fields

    basisCurve : Curve from PGeom2d;
    firstU     : Real from Standard;
    lastU      : Real from Standard;

end;
