-- Created on: 1993-04-06
-- Created by: Philippe DAUTRY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Parabola from PGeom2d  
inherits Conic from PGeom2d

        --- Purpose :
        --  Defines the parabola in the parameterization range  :
        --  ]-infinite,+infinite[
        --  See Also : Parabola from Geom2d.

uses  Ax22d from gp 

is


  Create returns mutable Parabola from PGeom2d;
        ---Purpose : Creates a parabola with default values.
	---Level: Internal 


  Create (aPosition : Ax22d from gp; aFocalLength : Real)
    returns mutable Parabola from PGeom2d;
	---Purpose : Creates a Parabola with <aPosition> and <aFocalLength>
	--         as field values.
	---Level: Internal 


  FocalLength (me : mutable; aFocalLength : Real);
        ---Purpose :   Set the value  of   the  field focalLength with
        --         <aFocalLength>.
	---Level: Internal 


  FocalLength (me)  returns Real;
	---Purpose : Retruns the value of the field focalLength.
	---Level: Internal 


fields

  focalLength : Real;

end;
