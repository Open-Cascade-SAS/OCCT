-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class StyleContextSelect from StepVisual inherits SelectType from StepData

	-- <StyleContextSelect> is an EXPRESS Select Type construct translation.
	-- it gathers : Representation, RepresentationItem, PresentationSet

uses

	Representation from StepRepr,
	RepresentationItem from StepRepr,
	PresentationSet from StepVisual
is

	Create returns StyleContextSelect;
	---Purpose : Returns a StyleContextSelect SelectType

	CaseNum (me; ent : Transient) returns Integer;
	---Purpose: Recognizes a StyleContextSelect Kind Entity that is :
	--        1 -> Representation
	--        2 -> RepresentationItem
	--        3 -> PresentationSet
	--        0 else

	Representation (me) returns any Representation;
	---Purpose : returns Value as a Representation (Null if another type)

	RepresentationItem (me) returns any RepresentationItem;
	---Purpose : returns Value as a RepresentationItem (Null if another type)

	PresentationSet (me) returns any PresentationSet;
	---Purpose : returns Value as a PresentationSet (Null if another type)


end StyleContextSelect;

