-- Created on: 1994-03-23
-- Created by: Bruno DUMORTIER
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package Geom2dAPI

	---Purpose: The  Geom2dAPI  package  provides  an  Application
	--          Programming Interface for the Geometry.
	--          
	--          The API is a set of classes aiming to provide :
	--          
	--          * High level and simple calls  for the most common
	--          operations. 
	--          
	--          *    Keeping   an   access  on    the    low-level
	--          implementation of high-level calls.
	--          
	-- 	    
	-- 	    The API  provides classes to  call the algorithmes
	-- 	    of the Geometry
	-- 	    
	-- 	    * The  constructors  of the classes  provides  the
	-- 	    different constructions methods.
	-- 	    
	-- 	    * The  class keeps as fields the   different tools
	-- 	    used by the algorithmes
	-- 	    
	-- 	    *   The class  provides  a  casting  method to get
	-- 	    automatically the  result  with  a   function-like
	-- 	    call. 
	-- 	    
	-- 	    For example to evaluate the distance <D> between a
	-- 	    point <P> and a curve <C>, one can writes :
	-- 	    
	-- 	        D = Geom2dAPI_ProjectPointOnCurve(P,C);
	-- 	    
	-- 	    or
	-- 	    
	-- 	        Geom2dAPI_ProjectPointOnCurve PonC(P,C);
	-- 	        D = PonC.LowerDistance();
	-- 	    


uses

    Geom2d,
    gp,
    TColgp,
    Extrema,
    Geom2dAdaptor,
    Geom2dInt,
    GeomAbs,
    TColStd,
    Quantity, 
    Approx,
    StdFail
    

is

    ------------------------------------------------------------------
    -- This classes  provides algo  to  evaluate  the distance between
    -- points and curves, curves and curves. 
    ------------------------------------------------------------------

    class ProjectPointOnCurve;

    class ExtremaCurveCurve;
    


    ------------------------------------------------------------------
    -- This classes provides algo to evaluate a curve  passing through
    -- an array of points.
    ------------------------------------------------------------------

    --- Approximation:
    --  
    class PointsToBSpline;
    
    
    --- Interpolation:
    --
    class Interpolate;
    
    
    ------------------------------------------------------------------
    -- This classes provides algo to evaluate an intersection between 
    -- two 2d-Curves.
    ------------------------------------------------------------------

    class InterCurveCurve;


end Geom2dAPI;
