-- Created on: 1997-07-29
-- Created by: Denis PASCAL 
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- modified     Sergey Zaritchny


class Constraint from PDataXtd inherits Attribute from PDF

	---Purpose: 

uses Integer          from Standard,
     Real             from PDataStd,
     HAttributeArray1 from PDF,
     NamedShape       from PNaming
    
is

    Create returns mutable Constraint from  PDataXtd;
    
    
    Create (Type        : Integer          from Standard;
    	    Geometries  : HAttributeArray1 from PDF;
    	    Value       : Real             from PDataStd;
    	    Plane       : NamedShape       from PNaming) 
    returns mutable Constraint from PDataXtd;
    
    
    GetValue (me) returns Real from PDataStd;
    

    GetType (me) returns Integer from Standard;
    
    
    GetGeometries (me) returns HAttributeArray1 from PDF;
    
    
    Set (me : mutable; V : Real from PDataStd);


    SetType (me : mutable; Type : Integer from Standard);
    
    
    SetGeometries (me : mutable; Geometries : HAttributeArray1 from PDF);
    
    SetPlane (me : mutable; plane : NamedShape from PNaming);
    GetPlane (me)
    returns NamedShape from PNaming;
    
    Verified(me:mutable; status : Boolean from Standard);
    Verified(me) 
    returns Boolean from Standard;    

    Inverted(me:mutable; status : Boolean from Standard);
    Inverted(me) 
    returns Boolean from Standard;    

    Reversed(me:mutable; status : Boolean from Standard);
    Reversed(me) 
    returns Boolean from Standard;    
    
fields

    myType       : Integer          from Standard;
    myGeometries : HAttributeArray1 from PDF;
    myValue      : Real             from PDataStd;
    myIsReversed : Boolean          from Standard;
    myIsInverted : Boolean          from Standard;
    myIsVerified : Boolean          from Standard;
    myPlane      : NamedShape       from PNaming;
    
end Constraint;
