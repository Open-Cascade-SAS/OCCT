-- Created on: 2000-01-19
-- Created by: data exchange team
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package XSAlgo 

    ---Purpose: 

uses

    MMgt,
    Geom,
    Geom2d,
    TopoDS,
    ShapeExtend,
    ShapeAnalysis,
    ShapeFix,
    Transfer,
    Message
    
is

    enumeration Caller is
    	---Purpose: Identifies the caller of the algorithm
      DEFAULT,
      IGES,
      STEP
    end Caller;

    class ToolContainer;
    	---Purpose: Returns tools used by AlgoContainer

    class AlgoContainer;
    	---Purpose: Provides initerface to the algorithms from Shape Healing
	--          and others for XSTEP processors.

    
    Init;
    	---Purpose: Creates and initializes default AlgoContainer.
    
    SetAlgoContainer (aContainer: AlgoContainer from XSAlgo);
    	---Purpose: Sets default AlgoContainer

    AlgoContainer returns AlgoContainer from XSAlgo;
    	---Purpose: Returns default AlgoContainer

end XSAlgo;
