-- Created on: 1995-12-04
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package RWStepGeom 

uses

	StepData, Interface, TCollection, TColStd, StepGeom

is


--class ReadWriteModule;

--class GeneralModule;

class RWAxis1Placement;
class RWAxis2Placement2d;
class RWAxis2Placement3d;
class RWBSplineCurve;
class RWBSplineCurveWithKnots;
class RWBSplineSurface;
class RWBSplineSurfaceWithKnots;
class RWBezierCurve;
class RWBezierSurface;
class RWBoundaryCurve;
class RWBoundedCurve;
class RWBoundedSurface;
class RWCartesianPoint;
class RWCartesianTransformationOperator;
class RWCartesianTransformationOperator3d;
class RWCircle;
class RWCompositeCurve;
class RWCompositeCurveOnSurface;
class RWCompositeCurveSegment;
class RWConic;
class RWConicalSurface;
class RWCurve;
class RWCurveBoundedSurface;
class RWCurveReplica;
class RWCylindricalSurface;
class RWDegeneratePcurve;
class RWDegenerateToroidalSurface;
class RWDirection;
class RWElementarySurface;
class RWEllipse;
class RWEvaluatedDegeneratePcurve;
class RWGeometricRepresentationContext;
class RWGeometricRepresentationContextAndGlobalUnitAssignedContext;
-- added by FMA:
class RWGeometricRepresentationContextAndParametricRepresentationContext;
-- added by FMA:
class RWGeomRepContextAndGlobUnitAssCtxAndGlobUncertaintyAssCtx; 
class RWGeometricRepresentationItem;
class RWHyperbola;
class RWIntersectionCurve;
class RWLine;
class RWOffsetCurve3d;
class RWOffsetSurface;
class RWOuterBoundaryCurve;
class RWParabola;
class RWPcurve;
class RWPlacement;
class RWPlane;
class RWPoint;
class RWPointOnCurve;
class RWPointOnSurface;
class RWPointReplica;
class RWPolyline;
class RWQuasiUniformCurve;
class RWQuasiUniformSurface;
class RWRationalBSplineCurve;
class RWRationalBSplineSurface;
class RWRectangularCompositeSurface;
class RWRectangularTrimmedSurface;
class RWReparametrisedCompositeCurveSegment;
class RWSeamCurve;
class RWSphericalSurface;
class RWSurface;
class RWSurfaceCurve;
class RWSurfaceOfLinearExtrusion;
class RWSurfaceOfRevolution;
class RWSurfaceCurveAndBoundedCurve;
class RWSurfacePatch;
class RWSurfaceReplica;
class RWSweptSurface;
class RWToroidalSurface;
class RWTrimmedCurve;
class RWUniformCurve;
class RWUniformSurface;
class RWOrientedSurface; --  Added from AP214 DIS to IS 4.01.2002
class RWVector;

class RWUniformCurveAndRationalBSplineCurve;
class RWBSplineCurveWithKnotsAndRationalBSplineCurve;
class RWQuasiUniformCurveAndRationalBSplineCurve;
class RWBezierCurveAndRationalBSplineCurve;
class RWBSplineSurfaceWithKnotsAndRationalBSplineSurface;
class RWUniformSurfaceAndRationalBSplineSurface;
class RWQuasiUniformSurfaceAndRationalBSplineSurface;
class RWBezierSurfaceAndRationalBSplineSurface;

	---Package Method ---

--	Init;
	---Purpose: enforced the initialisation of the  libraries

end RWStepGeom;
