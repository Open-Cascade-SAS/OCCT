-- Created on: 1991-01-30
-- Created by: Arnaud BOUZY
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class LessThan from Expr

inherits SingleRelation from Expr

uses GeneralExpression from Expr,
    GeneralRelation from Expr,
    AsciiString from TCollection

raises NumericError from Standard

is

    Create(exp1 : GeneralExpression ; exp2 : GeneralExpression)
    ---Purpose: Creates the relation <exp1> < <exp2>.
    returns LessThan;

    IsSatisfied(me)
    returns Boolean;

    Simplified(me)
    ---Purpose: Returns a GeneralRelation after replacement of
    --          NamedUnknowns by an associated expression, and after
    --          values computation.
    returns GeneralRelation
    raises NumericError;
    
    Simplify(me : mutable)
    ---Purpose: Replaces NamedUnknowns by associated expressions,
    --          and computes values in <me>.
    raises NumericError;
    
    Copy(me)
    ---Purpose: Returns a copy of <me> having the same unknowns and functions.
    returns like me;
    
    String(me)
    ---Purpose: returns a string representing <me> in a readable way.
    returns AsciiString;

end LessThan;
