-- Created on: 1991-06-24
-- Created by: Christophe MARION
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- modified by mps (dec 96)  add of  ContinuityCommands



package GeometryTest 

	---Purpose: this  package  provides  commands for  curves  and
	--          surface.
uses
    Draw,
    Standard, 
    GeomliteTest

is

    AllCommands(I : in out Interpretor from Draw);
	---Purpose: defines all geometric commands.
    
    CurveCommands(I : in out Interpretor from Draw);
	---Purpose: defines curve commands.
    
    FairCurveCommands(I : in out Interpretor from Draw);
	---Purpose: defines fair curve commands.
    
    SurfaceCommands(I : in out Interpretor from Draw);
	---Purpose: defines surface commands.

    ConstraintCommands(I : in out Interpretor from Draw);
	---Purpose: defines cosntrained curves commands.
    
    API2dCommands(I : in out Interpretor from Draw);
	---Purpose: defines commands to test the Geom2dAPI
	--          - Intersection
	--          - Extrema
	--          - Projection
	--          - Approximation, interpolation
    
    APICommands(I : in out Interpretor from Draw);
	---Purpose: defines commands to test the Geom2dAPI
	--          - Intersection
	--          - Extrema
	--          - Projection
	--          - Approximation, interpolation
 
    ContinuityCommands(I : in out Interpretor from Draw);
        --- Purpose: defines commands to check local
        --          continuity between curves or surfaces

    PolyCommands(I : in out Interpretor from Draw);
	---Purpose: defines     command  to    test  the    polyhedral
	--          triangulations and the polygons from the Poly package.
    
    TestProjCommands(I : in out Interpretor from Draw);
	---Purpose: defines commands to test projection of geometric objects
    
end GeometryTest;
