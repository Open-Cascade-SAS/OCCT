-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class BooleanOperand from StepShape 

    -- inherits SelectType from StepData

	-- <BooleanOperand> is an EXPRESS Select Type construct translation.
	-- it gathers : SolidModel, HalfSpaceSolid, CsgPrimitive, BooleanResult

uses

	SolidModel,
	HalfSpaceSolid,
	CsgPrimitive,
	BooleanResult
is

    Create returns BooleanOperand;
    ---Purpose : Returns a BooleanOperand SelectType

    SetTypeOfContent(me : in out; aTypeOfContent : Integer);

    TypeOfContent(me) returns Integer;
    	-- 1 : SolidModel,
    	-- 2 : HalfSpaceSolid,
    	-- 3 : CsgPrimitive,
    	-- 4 : BooleanResult

    SolidModel (me) returns any SolidModel;
    ---Purpose : returns Value as a SolidModel (Null if another 
    --         type)

    SetSolidModel(me : in out;
    	    	  aSolidModel : SolidModel from StepShape);

    HalfSpaceSolid (me) returns any HalfSpaceSolid;
    ---Purpose : returns Value as a HalfSpaceSolid (Null if 
    --         another type)

    SetHalfSpaceSolid(me : in out; 
    	    	      aHalfSpaceSolid : HalfSpaceSolid from StepShape);

    CsgPrimitive (me) returns CsgPrimitive;
    ---Purpose : returns Value as a CsgPrimitive (Null if another 
    --           type)
    --           CsgPrimitive is another Select Type

    SetCsgPrimitive(me : in out; 
    	    	    aCsgPrimitive : CsgPrimitive from StepShape);

    BooleanResult (me) returns any BooleanResult;
    ---Purpose : returns Value as a BooleanResult (Null if another 
    --           type)

    SetBooleanResult(me:in out;
    	    	     aBooleanResult : BooleanResult from StepShape);
    
fields

    theSolidModel     : SolidModel     from StepShape;
    theHalfSpaceSolid : HalfSpaceSolid from StepShape;
    theCsgPrimitive   : CsgPrimitive   from StepShape;  -- Select Type
    theBooleanResult  : BooleanResult  from StepShape;
    theTypeOfContent  : Integer        from Standard;

end BooleanOperand;

