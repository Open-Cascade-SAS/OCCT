-- Created on: 1997-12-01
-- Created by: Jean-Louis Frenkel
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class  ReferenceIterator from PCDM inherits Transient from Standard

uses MetaData from CDM,  
    SequenceOfReference from PCDM,  
    Document from CDM, Application from CDM,
    MessageDriver from  CDM
is
    Create (theMessageDriver : MessageDriver from  CDM)
    returns ReferenceIterator from PCDM;
    ---Purpose:  Warning! The constructor does not initialization.


    LoadReferences(me: mutable; aDocument: Document from CDM; aMetaData: MetaData from CDM; anApplication: Application from CDM; UseStorageConfiguration: Boolean from Standard);
    

    Init(me: mutable;aMetaData: MetaData from CDM)
    is virtual;
  
    More(me) returns Boolean from Standard
    is virtual private;

    Next(me: mutable)
    is virtual private;
    
    MetaData(me;UseStorageConfiguration: Boolean from Standard ) 
    returns MetaData from CDM
    is virtual private;


    ReferenceIdentifier(me)  returns Integer from Standard
    is virtual private;

    DocumentVersion(me) returns Integer from Standard
    ---Purpose: returns the version of the document in the reference
    is virtual private;
    
fields
    myReferences: SequenceOfReference from PCDM;
    myIterator: Integer from Standard; 
    myMessageDriver : MessageDriver from CDM; 
   
end ReferenceIterator from PCDM;
