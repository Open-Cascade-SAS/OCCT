-- Created on: 1992-08-26
-- Created by: Remi GILET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MakeScale2d

from gce

    ---Purpose: This class implements an elementary construction algorithm for
    -- a scaling transformation in 2D space. The result is a gp_Trsf2d transformation.
    -- A MakeScale2d object provides a framework for:
    -- -   defining the construction of the transformation,
    -- -   implementing the construction algorithm, and
    -- -   consulting the result.

uses Pnt2d  from gp,
     Trsf2d from gp,
     Real   from Standard
     
is

Create(Point : Pnt2d from gp      ;
       Scale : Real  from Standard) returns MakeScale2d;
    --- Purpose:
    -- Constructs a scaling transformation with:
    -- -   Point as the center of the transformation, and
    -- -   Scale as the scale factor.
        
Value(me) returns Trsf2d from gp
    is static;
    ---C++: return const&
    ---Purpose: Returns the constructed transformation.

Operator(me) returns Trsf2d from gp
    is static;
    ---C++: return const&
    ---C++: alias "Standard_EXPORT operator gp_Trsf2d() const;"

fields

    TheScale2d : Trsf2d from gp;

end MakeScale2d;

