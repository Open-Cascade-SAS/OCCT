-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Update:
--              20-01-2009 : ABD Integration support of system fonts (using FTGL and FreeType)

package OSD

 ---History:
 --   Version   Date        Purpose
 --   1.1   24/06/92    Operating System Dependent tools
 --   1.2
 --   2.0
 --   3.0
 --   Windows NT 30/09/96 ( EUG )
 ---Purpose: Set of Operating Sytem Dependent Tools
 --         (O)perating (S)ystem (D)ependent

uses

    Standard ,
    Quantity ,
    TCollection

is

 exception OSDError inherits Failure from Standard  ;

 imported Function;
   ---Purpose: This is in fact a pointer to a function.
   --          This is not an "enumeration" but a trick to solve an omission
   --          from CDL.
   --- C++: alias "typedef int (* OSD_Function)(...);"

 enumeration OEMType is Unavailable,SUN,DEC,SGI,NEC,MAC,PC,HP,IBM,VAX,LIN,AIX;
   ---Purpose: This is set of possible machine types
   --          used in OSD_Host::MachineType

 enumeration SysType is Unknown,Default,UnixBSD, UnixSystemV, VMS, OS2,
                        OSF, MacOs, Taligent, WindowsNT, LinuxREDHAT,Aix;
   ---Purpose: Thisd is a set of possible system types.
   --          'Default' means SysType of machine operating this process.
   --          This can be used with the Path class.
   --          All UNIX-like are grouped under "UnixBSD" or "UnixSystemV".
   --          Such systems are Solaris, NexTOS ...
   --          A category of systems accept MSDOS-like path such as
   --          WindowsNT and OS2.

 enumeration FromWhere is FromBeginning, FromHere, FromEnd;
   ---Purpose: Used by OSD_File in the method Seek.

 enumeration LockType is NoLock, ReadLock, WriteLock, ExclusiveLock;
   ---Purpose: locks for files.
   --          NoLock is the default value when opening a file.
   --
   --          ReadLock allows only one reading of the file at a time.
   --
   --          WriteLock prevents others writing into a file(excepted the user
   --          who puts the lock)but allows everybody to read.
   --
   --          ExclusiveLock prevents reading and writing except for the
   --          current user of the file.
   --          So ExclusiveLock means only one user on the file and this
   --          user is the one who puts the lock.

 enumeration SingleProtection is None,R,W,RW,X,RX,WX,RWX,D,RD,WD,RWD,XD,RXD,WXD,RWXD;
   ---Purpose: Access rights for files.
   --          R means Read, W means Write, X means eXecute and D means Delete.
   --          On UNIX, the right to Delete is combined with Write access.
   --          So if "W"rite is not set and "D"elete is, "W"rite will be set
   --          and if "W" is set, "D" will be too.

 enumeration OpenMode is ReadOnly, WriteOnly, ReadWrite;
   ---Purpose: Specifies the file open mode.

 enumeration LoadMode is RTLD_LAZY, RTLD_NOW;
   ---Purpose: This enumeration is used to load shareable libraries.

 enumeration KindFile is FILE, DIRECTORY, LINK, SOCKET, UNKNOWN;
   ---Purpose: Specifies the type of files.

 private enumeration WhoAmI is  WDirectory, WDirectoryIterator,
             WEnvironment, WFile, WFileNode, WFileIterator,
             WPath, WProcess, WProtection, WHost, WDisk,
             WChronometer, WTimer, WPackage, WPrinter,
             WEnvironmentIterator;
   ---Purpose: Allows great accuracy for error management.
   --          This is private.


         class Error;
             ---Purpose: Accurate management of OSD specific errors.

         class Protection;
             ---Purpose: Gets and sets protection attributes of 'system , user ,
             --          group, and world'.

         class Path;
             ---Purpose: Manages independent system path translation.

         deferred class FileNode;
             ---Purpose: A set of file/directory manipulation tools.

         class Disk;
             ---Purpose: A set of disk oriented tools.

         class File;
             ---Purpose: A set of file oriented tools.

         class FileIterator;
             ---Purpose: Searches for child files in current directory.

         class Directory;
             ---Purpose: A set of directory oriented tools

         class DirectoryIterator;
             ---Purpose: Searches sub-directories in current directory.

         class Chronometer;
             ---Purpose: Measures time elapsed for performance program tests.
             --          Measures CPU time consumed by a method call.

         class Timer;
             ---Purpose: Measures the effective time elapsed for a method call.

         class Printer;
             ---Purpose: Selects a printer (used by File).

         class Host;
             ---Purpose: Carries information about a host.
             --          System version ,host name, nodename ...

         class Environment;
             ---Purpose: Manages environment variables.

         class EnvironmentIterator;
             ---Purpose: Get all environment variables.

         class Process;
             ---Purpose: Process specific oriented tools

--         class Mutex is alias Mutex from Standard;
             ---Purpose: Mutex object to synchronize threads within one process

         class SharedLibrary;
             ---Purpose: Provides tools to load a shared library
             --          and retrieve the address of an entry point.

     imported MemInfo;
     imported PThread;
     imported ThreadFunction;
         class Thread;
             ---Purpose: A tool to manage threads

    -----------------------------------------------
    --  UNIX specific exceptions and enumeration --
    -----------------------------------------------

    exception Signal  inherits Failure from  Standard;
    exception SIGHUP  inherits Signal;
    exception SIGINT  inherits Signal;
    exception SIGQUIT inherits Signal;
    exception SIGILL  inherits Signal;
    exception SIGKILL inherits Signal;
    exception SIGBUS  inherits Signal;
    exception SIGSEGV inherits Signal;
    exception SIGSYS  inherits Signal;

    ----------------------------------------
    -- Exceptions ( Windows NT specific ) --
    ----------------------------------------

    exception Exception inherits Failure   from  Standard;

    exception Exception_ACCESS_VIOLATION         inherits Exception;
    exception Exception_ARRAY_BOUNDS_EXCEEDED    inherits Exception;
    exception Exception_FLT_DENORMAL_OPERAND     inherits Exception;
    exception Exception_FLT_DIVIDE_BY_ZERO       inherits Exception;
    exception Exception_FLT_INEXACT_RESULT       inherits Exception;
    exception Exception_FLT_INVALID_OPERATION    inherits Exception;
    exception Exception_FLT_OVERFLOW             inherits Exception;
    exception Exception_FLT_STACK_CHECK          inherits Exception;
    exception Exception_FLT_UNDERFLOW            inherits Exception;
    exception Exception_ILLEGAL_INSTRUCTION      inherits Exception;
    exception Exception_IN_PAGE_ERROR            inherits Exception;
    exception Exception_INT_DIVIDE_BY_ZERO       inherits Exception;
    exception Exception_INT_OVERFLOW             inherits Exception;
    exception Exception_INVALID_DISPOSITION      inherits Exception;
    exception Exception_NONCONTINUABLE_EXCEPTION inherits Exception;
    exception Exception_PRIV_INSTRUCTION         inherits Exception;
    exception Exception_STACK_OVERFLOW           inherits Exception;
    exception Exception_STATUS_NO_MEMORY         inherits Exception; -- generating by 'HeapAlloc'
    exception Exception_CTRL_BREAK               inherits Exception; -- generating by 'Ctrl-C' keystroke

    SetSignal(theFloatingSignal: Boolean = Standard_True);
    ---Purpose:
    -- Sets signal and exception handlers.
    -- <b>Windows-specific notes<\b>
    -- Compiled with MS VC++ sets 3 main handlers:
    -- @li Signal handlers (via ::signal() functions) that translate system signals
    --     (SIGSEGV, SIGFPE, SIGILL) into C++ exceptions (classes inheriting
    --     Standard_Failure). They only be called if user calls ::raise() function
    --     with one of supported signal type set.
    -- @li Exception handler OSD::WntHandler() (via ::SetUnhandledExceptionFilter())
    --     that will be used when user's code is compiled with /EHs option.
    -- @li Structured exception (SE) translator (via _set_se_translator()) that
    --     translates SE exceptions (aka asynchronous exceptions) into the
    --     C++ exceptions inheriting Standard_Failure. This translator will be
    --     used when user's code is compiled with /EHa option.
    -- .
    -- This approach ensures that regardless of the option the user chooses to
    -- compile his code with (/EHs or /EHa), signals (or SE exceptions) will be
    -- translated into Open CASCADE C++ exceptions.
    -- .
    -- If @a theFloatingSignal is TRUE then floating point exceptions will be
    -- generated in accordance with the mask
    -- <tt>_EM_INVALID | _EM_DENORMAL | _EM_ZERODIVIDE | _EM_OVERFLOW<\tt> that is
    -- used to call ::_controlfp() system function. If @a theFloatingSignal is FALSE
    -- corresponding operations (e.g. division by zero) will gracefully complete
    -- without an exception.
    -- .
    -- <b>Unix-specific notes<\b>
    -- OSD::SetSignal() sets handlers (via ::sigaction()) for multiple signals
    -- (SIGFPE, SIGSEGV, etc). Currently the number of handled signals is much
    -- greater than for Windows, in the future this may change to provide better
    -- consistency with Windows.
    -- .
    -- @a theFloatingSignal is recognized on Sun Solaris, Linux, and SGI Irix to
    -- generate floating-point exception according to the mask
    -- <tt>FE_INVALID | FE_DIVBYZERO | FE_OVERFLOW</tt> (in Linux conventions).<br>
    -- When compiled with OBJS macro defined, already set signal handlers (e.g.
    -- by Data Base Managers) are not redefined.
    -- .
    -- <b>Common notes<\b>
    -- If OSD::SetSignal() method is used in at least one thread, it must also be
    -- called in any other thread where Open CASCADE will be used, to ensure
    -- consistency of behavior. Its @a aFloatingSignal argument must be consistent
    -- across threads.
    -- .
    -- Keep in mind that whether the C++ exception will really be thrown (i.e.
    -- ::throw() will be called) is regulated by the NO_CXX_EXCEPTIONS and
    -- OCC_CONVERT_SIGNALS macros used during compilation of Open CASCADE and
    -- user's code. Refer to Foundation Classes User's Guide for further details.
    --

    AvailableMemory returns Integer from Standard;
    ---Purpose: Returns available memory in Kilobytes.
    ---Level: Advanced

    SecSleep(aDelay: Integer from Standard);
    ---Purpose: Commands the process to sleep for a number of seconds.
    ---Level: Public

    MilliSecSleep(aDelay: Integer from Standard);
    ---Purpose: Commands the process to sleep for a number of milliseconds
    ---Level: Public

    RealToCString(aReal: Real; aString:out PCharacter)
        returns Boolean ;
    ---Purpose:
    --  Converts aReal into aCstring in exponential format with a period as
    --  decimal point, no thousand separator and no grouping of digits.
    --  The conversion is independant from the current locale
    ---Level: Public

    CStringToReal(aString: CString; aReal: out Real) returns Boolean ;
    ---Purpose:
    --  Converts aCstring representing a real with a period as
    --  decimal point, no thousand separator and no grouping of digits
    --  into aReal .
    --  The conversion is independant from the current locale.
    ---Level: Public

    IsDivisible(aDividend, aDivisor: Real from Standard)
    returns Boolean from Standard;
    ---Purpose: Tests if the quotient theDividend/theDivisor
    --          does not overflow
    ---Level: Public

    GetExponent(aReal: Real from Standard)
    returns Integer from Standard;
    ---Purpose: Returns the exponent in base 2 of a floating-point number.
    ---Level: Public

    GetMantissa(aReal: Real from Standard)
    returns Real from Standard;
    ---Purpose: Returns the mantissa of a floating-point number.
    ---Level: Public

    -------------------------
    -- Windows NT specific --
    -------------------------

    ControlBreak raises  Exception_CTRL_BREAK;
    ---Purpose: since Windows NT does not support 'SIGINT' signal like UNIX,
    --          then this method checks whether Ctrl-Break keystroke was or
    --          not. If yes then raises Exception_CTRL_BREAK.

end OSD;
