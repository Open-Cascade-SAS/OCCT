-- File:	StepShape_EdgeBasedWireframeModel.cdl
-- Created:	Fri Dec 28 16:02:01 2001 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class EdgeBasedWireframeModel from StepShape
inherits GeometricRepresentationItem from StepGeom

    ---Purpose: Representation of STEP entity EdgeBasedWireframeModel

uses
    HAsciiString from TCollection,
    HArray1OfConnectedEdgeSet from StepShape

is
    Create returns EdgeBasedWireframeModel from StepShape;
	---Purpose: Empty constructor

    Init (me: mutable; aRepresentationItem_Name: HAsciiString from TCollection;
                       aEbwmBoundary: HArray1OfConnectedEdgeSet from StepShape);
	---Purpose: Initialize all fields (own and inherited)

    EbwmBoundary (me) returns HArray1OfConnectedEdgeSet from StepShape;
	---Purpose: Returns field EbwmBoundary
    SetEbwmBoundary (me: mutable; EbwmBoundary: HArray1OfConnectedEdgeSet from StepShape);
	---Purpose: Set field EbwmBoundary

fields
    theEbwmBoundary: HArray1OfConnectedEdgeSet from StepShape;

end EdgeBasedWireframeModel;
