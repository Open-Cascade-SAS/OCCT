-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package TColStd 

                             
uses TCollection

is

    imported PackedMapOfInteger; 
    imported MapIteratorOfPackedMapOfInteger;


--                  Instantiations de TCollection                         --
--                  *****************************                         --
------------------------------------------------------------------------
 
    class HPackedMapOfInteger; 
 
    imported Array1OfInteger;
    imported Array1OfReal;
    imported Array1OfCharacter;
    imported Array1OfBoolean;
    imported Array1OfAsciiString;
    imported Array1OfExtendedString;
    imported Array1OfTransient;
    imported Array1OfByte;


    imported transient class HArray1OfInteger;
    imported transient class HArray1OfReal;
    imported transient class HArray1OfCharacter;
    imported transient class HArray1OfBoolean;
    imported transient class HArray1OfAsciiString;
    imported transient class HArray1OfExtendedString;
    imported transient class HArray1OfTransient;
    imported transient class HArray1OfByte;


    imported Array2OfInteger;
    imported Array2OfReal;
    imported Array2OfCharacter;
    imported Array2OfBoolean;
    imported Array2OfTransient;


    imported transient class HArray2OfInteger;
    imported transient class HArray2OfReal;
    imported transient class HArray2OfCharacter;
    imported transient class HArray2OfBoolean;
    imported transient class HArray2OfTransient;

imported SequenceOfInteger;
imported SequenceOfReal; 
imported SequenceOfAsciiString;
imported SequenceOfHAsciiString;
imported SequenceOfExtendedString;
imported SequenceOfHExtendedString;
imported SequenceOfTransient;
imported SequenceOfAddress;
imported SequenceOfBoolean;


imported transient class HSequenceOfInteger;
imported transient class HSequenceOfReal;
imported transient class HSequenceOfAsciiString;
imported transient class HSequenceOfHAsciiString;
imported transient class HSequenceOfExtendedString;
imported transient class HSequenceOfHExtendedString;
imported transient class HSequenceOfTransient;

--                    
--       Instantiations List (Integer,Real,Transient)
--       ********************************************
--       
imported ListOfInteger;
imported ListIteratorOfListOfInteger;
imported ListOfReal;
imported ListIteratorOfListOfReal;
imported ListOfTransient;
imported ListIteratorOfListOfTransient;
imported ListOfAsciiString;
imported ListIteratorOfListOfAsciiString;

--                    
--       Instantiations MapHasher (Integer,Real, Transient, Persistent)
--       **************************************************************
--       
imported MapIntegerHasher;
imported MapRealHasher;
imported MapTransientHasher;


--       Instantiations Map (Integer, Real, Transient, Persistent)
--       *********************************************************
--       
imported MapOfInteger;
imported MapIteratorOfMapOfInteger;
imported MapOfReal;
imported MapIteratorOfMapOfReal;
imported MapOfTransient;
imported MapIteratorOfMapOfTransient;
imported MapOfAsciiString;
imported MapIteratorOfMapOfAsciiString;

--                    
--       Instantiations IndexedMap (Integer, Real, Transient, Persistent)
--       ****************************************************************
--       
imported IndexedMapOfInteger;
imported IndexedMapOfReal;
imported IndexedMapOfTransient;

imported IndexedDataMapOfTransientTransient; 

--                    
--       Instantiations DataMap
--       **********************
--       
imported DataMapOfIntegerReal;
imported DataMapIteratorOfDataMapOfIntegerReal;

imported DataMapOfIntegerInteger;

imported DataMapIteratorOfDataMapOfIntegerInteger;

imported DataMapOfIntegerListOfInteger;

imported DataMapIteratorOfDataMapOfIntegerListOfInteger;

imported DataMapOfTransientTransient;

imported DataMapIteratorOfDataMapOfTransientTransient;

imported DataMapOfAsciiStringInteger;

imported DataMapIteratorOfDataMapOfAsciiStringInteger;

imported DataMapOfIntegerTransient;

imported DataMapIteratorOfDataMapOfIntegerTransient;

imported DataMapOfStringInteger;

imported DataMapIteratorOfDataMapOfStringInteger;

--
--  Arrays of lists...
--  ******************
--

imported Array1OfListOfInteger;

imported transient class HArray1OfListOfInteger;

end TColStd;

