-- Created on: 1991-07-24
-- Created by: Michel CHAUVAT
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

private generic class FuncExtPC from Extrema 
(Curve    as any;
 Tool     as any;
 POnC     as any;
 Pnt      as any;
 Vec      as any)
						     
    inherits FunctionWithDerivative from math
    --- Purpose: Function to find extrema of the distance between a
    --- point and a curve.

uses    SequenceOfReal    from TColStd,
	SequenceOfInteger from TColStd
	
raises  OutOfRange   from Standard,
        TypeMismatch from Standard

private class SeqPC instantiates Sequence from TCollection(POnC);	


is

    Create returns FuncExtPC;

    Create (P: Pnt; C: Curve) returns FuncExtPC;
    	---Purpose: 

    Initialize(me: in out; C: Curve)
    	---Purpose: sets the field mycurve of the function.
    is static;
    
    SetPoint(me: in out; P: Pnt)
    	---Purpose: sets the field P of the function.
    is static;


    -- In all next methods, an exception is raised if the fields 
    -- were not initialized.

    Value (me: in out; U: Real; F: out Real) returns Boolean;
    	---Purpose: Calculation of F(U).

    Derivative (me: in out; U: Real; DF: out Real) returns Boolean;
    	---Purpose: Calculation of F'(U).

    Values (me: in out; U: Real; F,DF: out Real) returns Boolean;
    	---Purpose: Calculation of F(U) and F'(U).

    GetStateNumber (me: in out) returns Integer
    	---Purpose: Save the found extremum.
    	is redefined;

    NbExt (me) returns Integer
    	---Purpose: Return the nunber of found extrema.
    raises TypeMismatch from Standard;

    SquareDistance (me; N: Integer) returns Real
    	---Purpose: Returns the Nth distance.
    	raises  OutOfRange from Standard,
                TypeMismatch from Standard;
	    	-- if N < 1 or N > NbExt(me).

    IsMin (me; N: Integer) returns Boolean
    	---Purpose: Shows if the Nth distance is a minimum.
    	raises  OutOfRange from Standard,
                TypeMismatch from Standard;
	    	-- if N < 1 or N > NbExt(me).

    Point (me; N: Integer) returns POnC
        ---C++: return const &
    	---Purpose: Returns the Nth extremum.
    	raises  OutOfRange from Standard,
                TypeMismatch from Standard;
	    	-- if N < 1 or N > NbExt(me).

    SubIntervalInitialize(me: in out; theUfirst, theUlast: Real from Standard);
    	---Purpose: Determines boundaries of subinterval for find of root.
    
    SearchOfTolerance(me: in out) returns Real from Standard;
    	---Purpose: Computes a Tol value. If 1st derivative of curve
    	--          |D1|<Tol, it is considered D1=0.      
    

fields
    myP    : Pnt;
    myC    : Address from Standard;

    myU    : Real;          -- current
    myPc   : Pnt;           -- current point 
    myD1f  : Real;          -- value of derivative of the function

    mySqDist: SequenceOfReal    from TColStd;
    myIsMin: SequenceOfInteger from TColStd;
    myPoint: SeqPC;
    myPinit: Boolean;
    myCinit: Boolean;
    myD1Init: Boolean;
    
    myTol: Real from Standard;  -- toolerance for derivate

--Supremum of search 1st non-zero derivative    
    myMaxDerivOrder: Integer from Standard;
    
--boundaries of subinterval for find of root
    myUinfium, myUsupremum: Real from Standard;
    

end FuncExtPC;
