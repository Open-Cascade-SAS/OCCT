-- File:        SiUnitAndTimeUnit.cdl
-- Created:     Mon Dec  4 12:02:36 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWSiUnitAndTimeUnit from RWStepBasic

	---Purpose : Read & Write Module for SiUnitAndTimeUnit

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     SiUnitAndTimeUnit from StepBasic

is

	Create returns RWSiUnitAndTimeUnit;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable SiUnitAndTimeUnit from StepBasic);

	WriteStep (me; SW : in out StepWriter; ent : SiUnitAndTimeUnit from StepBasic);

end RWSiUnitAndTimeUnit;
