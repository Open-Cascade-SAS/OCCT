-- Created on: 1993-01-14
-- Created by: Philippe DAUTRY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class Builder from BRepSweep 

	---Purpose: implements the abstract Builder with the BRep Builder

uses
    Builder from BRep,
        
    Shape	from TopoDS,
    Shell	from TopoDS,
    Face	from TopoDS,
    Wire	from TopoDS,
    Edge	from TopoDS,
    Vertex	from TopoDS,
    
    Orientation from TopAbs
    
is

    Create(aBuilder : Builder from BRep) returns Builder from BRepSweep;
	---Purpose: Creates a Builder.
	
    Builder(me) returns Builder from BRep
	---C++: inline
	---C++: return const &
    is static;
	
        -- implements the Builder methods

    MakeCompound (me; aCompound : out Shape from TopoDS)
    	---Purpose: Returns an empty Compound.
    is static;

    MakeCompSolid (me; aCompSolid : out Shape from TopoDS)
    	---Purpose: Returns an empty CompSolid.
    is static;

    MakeSolid (me; aSolid : out Shape from TopoDS)
    	---Purpose: Returns an empty Solid.
    is static;

    MakeShell (me; aShell : out Shape from TopoDS)
    	---Purpose: Returns an empty Shell.
    is static;

    MakeWire (me; aWire : out Shape from TopoDS)
    	---Purpose: Returns an empty Wire.
    is static;

    
    Add(me; aShape1 : in out Shape from TopoDS; 
	    aShape2 : in     Shape from TopoDS;
    	    Orient  : in     Orientation from TopAbs)
    	---Purpose: Adds the Shape 1 in the Shape 2, set to
    	--          <Orient> orientation.
    is static;
    
    Add(me; aShape1 : in out Shape from TopoDS; 
	    aShape2 : in     Shape from TopoDS)
    	---Purpose: Adds the Shape 1 in the Shape 2.
    is static;

fields

    myBuilder : Builder from BRep;

end Builder;

