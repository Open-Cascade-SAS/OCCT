-- Created on: 2007-01-25
-- Created by: Sergey KOCHETKOV
-- Copyright (c) 2007-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SensitiveMesh from MeshVS inherits SensitiveEntity from Select3D

	---Purpose: This class provides custom mesh sensitive entity used in advanced mesh selection.  
    	---It provides detection of mesh entities accordingly to activated selection mode 

uses
  EntityOwner from SelectBasics,
  Array1OfPnt2d from TColgp, 
  Box from Bnd, 
  Box2d from Bnd, 
  Location from TopLoc, 
  Lin from gp, 
  ListOfBox2d from SelectBasics,
  PickArgs from SelectBasics,
  Projector from Select3D      
is

  Create ( theOwner    : EntityOwner from SelectBasics; 
           theMode     : Integer = 0 )
    returns mutable SensitiveMesh from MeshVS; 
      
  GetMode( me ) returns Integer from Standard;     
     
  GetConnected( me: mutable;  aLocation  :  Location from TopLoc )
    returns SensitiveEntity from Select3D is redefined; 

  Matches (me : mutable;
           thePickArgs : PickArgs from SelectBasics;
           theMatchDMin, theMatchDepth : out Real from Standard)
    returns Boolean is redefined;

  Matches  ( me: mutable;   XMin, YMin, XMax, YMax  : Real;
             	    	    aTol                    : Real ) returns Boolean  
    is redefined;

  Matches  ( me: mutable;   Polyline  :  Array1OfPnt2d from TColgp;
                            aBox      :  Box2d;  
    	    	    	    aTol      :  Real ) returns Boolean  
    is redefined; 
      
  Project ( me:mutable; aProjector : Projector from Select3D ) is redefined static;
     
  Areas   ( me: mutable ; boxes : in out ListOfBox2d from SelectBasics ) is redefined static;  
   
  ProjectOneCorner( me: mutable; aProjector : Projector from Select3D; 
    	    	    	    	 X,Y,Z      : Real from Standard ) is private;     
 
fields 
   
  myMode  : Integer from Standard;          
  mybox   : Box    from Bnd; 
  mybox2d : Box2d  from Bnd;   
 
end SensitiveMesh;
