-- Created on: 1995-05-30
-- Created by: Christian CAILLET
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

generic class JaggedArray  from Interface
    (TheKey as TShared)
    inherits TShared

    ---Purpose : This class allows to define an HArray1 Of HArray1 ...
    --           which is not possible with the actual system of
    --           genericity supported by CasCade

uses Array1OfTransient

is

    Create (low, up : Integer) returns mutable JaggedArray;

    Lower  (me) returns Integer;
    Upper  (me) returns Integer;
    Length (me) returns Integer;

    SetValue (me : mutable; num : Integer; val : any TheKey);

    Value (me; num : Integer) returns any TheKey;
    -- C++ : return const & (NO , DownCast required)

--    ChangeValue (me : mutable; num : Integer) returns any TheKey;
    -- C++ : return & (NO , DownCast required !)

fields

    thelist : Array1OfTransient;

end JaggedArray;
