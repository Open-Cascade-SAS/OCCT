-- Created on: 1994-08-31
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class VertexInfo from Draft

	---Purpose: 

uses Pnt                       from gp,
     Edge                      from TopoDS,
     ListOfShape               from TopTools,
     ListOfReal                from TColStd,
     ListIteratorOfListOfShape from TopTools

raises DomainError  from Standard,
       NoMoreObject from Standard

is

    Create
    
    	returns VertexInfo from Draft;
	
	
    Add(me: in out; E: Edge from TopoDS)
    
    	is static;


    Geometry(me)
    
    	returns Pnt from gp
	is static;
	---C++: return const&


    Parameter(me: in out; E: Edge from TopoDS)
    
    	returns Real from Standard
	raises DomainError from Standard
	is static;


    InitEdgeIterator(me: in out)

    	is static;

    
    Edge(me)
    	returns Edge from TopoDS
	is static;
	---C++: return const&


    NextEdge(me: in out)
    
    	raises NoMoreObject from Standard
    	is static;


    MoreEdge(me)
    
    	returns Boolean from Standard
	is static;



    ChangeGeometry(me: in out)
    
    	returns Pnt from gp
	is static;
	---C++: return &


    ChangeParameter(me: in out; E: Edge from TopoDS)
    
    	returns Real from Standard
	is static;
	---C++: return &


fields

    myGeom    : Pnt  from gp;
    myEdges   : ListOfShape from TopTools;
    myParams  : ListOfReal  from TColStd;
    myItEd    : ListIteratorOfListOfShape from TopTools;

end VertexInfo;
