-- Created on: 1992-09-04
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




package IntStart

    	---Purpose: This package provides generic algorithms to
    	--          find specific points (points on boundaries
    	--          and points inside a surface) used as starting
    	--          points for marching algorithms.

        ---Level: Internal
        --
        -- All the methods of the classes of this package are Internal.
	--

uses Standard, MMgt, TCollection, StdFail, TopAbs, GeomAbs, gp, IntSurf, math

is

    deferred generic class ArcTool;

    deferred generic class SOBTool;

    deferred generic class TopolTool;

    deferred generic class SOBFunction;

    generic class Segment;
    
    generic class PathPoint;

    generic class SearchOnBoundaries, ThePathPoint, SequenceOfPathPoint, 
                                      TheSegment, SequenceOfSegment;

    deferred generic class PSurfaceTool;

    deferred generic class SITool;

    deferred class SITopolTool;

    deferred generic class SIFunction;

    generic class SearchInside;


end IntStart;



