-- Created on: 1993-01-27
-- Created by: Philippe DAUTRY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



deferred generic class Iterator from Sweep (TheShape as any)

	---Purpose: This  is a  signature class describing   iteration
	--          services   required      by the Swept   Primitives
	--          algorithms from  a Directing or a Generating Line.
	--          This  tool is  used   to  iterate   on the  direct
	--          sub-shapes  of a  Shape. 
	--          

uses

    Orientation from TopAbs

raises

    NoMoreObject from Standard,
    NoSuchObject from Standard

is

    Init(me : in out; aShape: TheShape)
	---Purpose: Resest the Iterator on sub-shapes of <aShape>.
    is deferred;
    
    More(me) returns Boolean
	---Purpose: Returns True if there is a current sub-shape.
	--          
	-- -C++: inline
    is deferred;
    
    Next(me : in out)
	---Purpose: Moves to the next sub-shape.
    raises
    	NoMoreObject from Standard
    is deferred;
    
    Value(me) returns TheShape
	---Purpose: Returns the current sub-shape.
    raises
    	NoSuchObject from Standard
	-- -C++: return const &
	-- -C++: inline
    is deferred;
    
    Orientation(me) returns Orientation from TopAbs
	---Purpose: Returns the orientation of the current sub-shape.
    raises
    	NoSuchObject from Standard
	---C++: return const &
	---C++: inline
    is deferred;
    
end Iterator;
