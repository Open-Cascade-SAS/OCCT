-- Created on: 1998-11-10
-- Created by: Igor FEOKTISTOV
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class ElementsOfRefMatrix from FEmTool inherits  FunctionSet  from  math

	---Purpose: this  class  describes  the  functions  needed  for   
    	--          calculating  matrix  elements  of  RefMatrix  for  linear   
	--          criteriums  (Tension,  Flexsion  and  Jerk).
	--          Each  function  from  set  gives  value  Pi(u)'*Pj(u)'  or 
	--          Pi(u)''*Pj(u)''  or  Pi(u)'''*Pj(u)'''  for  each  i  and  j,  
    	--          where  Pi(u)  is  i-th  basis  function  of  expansion  and 
	--          (')  means  derivative.
uses 
    Vector  from  math, 
    Base  from  PLib

raises 
    ConstructionError  from  Standard

is 
    Create(TheBase  :  Base  from  PLib;  DerOrder  :  Integer  from  Standard)
    
     	--  DerOrder  is  order  of  derivative  (1,  2,  3)  
	 
    returns ElementsOfRefMatrix  from  FEmTool 
    raises  ConstructionError  from  Standard; 
    --  if  DerOrder  is  not  valid
     
    NbVariables(me)
    	---Purpose: returns the number of variables of the function. 
	--  It  is  supposed  that  NbVariables  =  1.

    returns Integer;

    
    
    NbEquations(me)
    	---Purpose: returns the number of equations of the function.

    returns Integer;
    
    
    Value(me: in out; X: Vector; F: out Vector)
    	---Purpose: computes the values <F> of the functions for the 
    	--          variable <X>.
    	--          returns True if the computation was done successfully, 
    	--          False otherwise. 
	--          F  contains  results  only  for  i<=j  in  following  order: 
	--          P0*P0,  P0*P1,  P0*P2...  P1*P1,  P1*P2,...  (upper  triangle of 
	--          matrix  {PiPj})

    returns Boolean;

fields 
    myBase  :  Base  from  PLib; 
    myDerOrder  :  Integer; 
    myNbEquations  :  Integer;

end ElementsOfRefMatrix;
