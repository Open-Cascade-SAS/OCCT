-- Created on: 2000-11-24
-- Created by: Michael KLOKOV
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class RoughShapeIntersector from BOPTools

   	---Purpose: The class RoughShapeIntersector describes the algorithm of
    	--         intersection of bounding boxes of 
    	--         shapes stored in ShapesDataStructure.
	--         It stores statuses of intersection in 2 dimension array.
    
uses
    Array1OfListOfInteger from TColStd,
    ListOfInteger         from TColStd, 
    HArray2OfIntersectionStatus from BOPTools,
    IntersectionStatus          from BOPTools, 
    HArray1OfBox from Bnd,
    PShapesDataStructure from BooleanOperations
is

    Create(PDS: PShapesDataStructure from BooleanOperations)  
    	returns RoughShapeIntersector from BOPTools;
	---Purpose:
	-- Initializes algorithm by shapes data structure
	--
    
    Perform(me: in out);
    	---Purpose: 
    	-- Perform computations.
	--
	--  Warning: 
    	-- Using this function, after the destructor of
    	-- the object pointed by PDS (see constructor)
    	-- was invoked, lead to crash.
	--
    
    TableOfStatus(me)
    	returns HArray2OfIntersectionStatus from BOPTools;
	---C++: return const &
	---Purpose:
	--  Returns 2 dimension array of status flags.
    	-- First indices of the array corresponds to indices of 
    	-- subshapes of Object of myPDS.
    	-- Second indices of array corresponds to indices of 
    	-- subshapes of Tool of myPDS.
	--

    IsDone(me) returns Boolean from Standard;
    	---Purpose:
	-- Returns False if some errors occured during
	-- computations or method Perform
	-- was not invoked before, 
    	-- otherwise returns True.
	--
    
    --    private methods
    Prepare(me: in out)  
    	is private;

    PropagateForSuccessors1(me: in out; AncestorsIndex1: Integer from Standard;
    	    	    	    	    	AncestorsIndex2: Integer from Standard;
    	    	    	    	    	theStatus      : IntersectionStatus from BOPTools)
    	is private;

    PropagateForSuccessors2(me: in out; AncestorsIndex1: Integer from Standard;
    	    	    	    	    	AncestorsIndex2: Integer from Standard;
    	    	    	    	    	theStatus      : IntersectionStatus from BOPTools)
    	is private;

fields   
    myPDS: PShapesDataStructure from BooleanOperations;
    myBoundingBoxes: HArray1OfBox from Bnd;
    
    myTableOfStatus: HArray2OfIntersectionStatus from BOPTools;
    ---Purpose: First indices of array corresponds to indices of subshapes of Object of myPDS.
    --          Second indices of array corresponds to indices of subshapes of Tool of myPDS.
    
    myIsDone: Boolean from Standard;
       
end RoughShapeIntersector from BOPTools;

