-- Created on: 1991-04-15
-- Created by: Philippe DAUTRY
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


generic class QualifiedCurv from GccEnt (TheCurve as any)

	---Purpose: Creates a qualified 2d line.

uses Position from GccEnt

is

Create(Curve     : TheCurve                ;
       Qualifier : Position from GccEnt ) 
returns QualifiedCurv from GccEnt;
-- is private;

Qualified(me) returns TheCurve
is static;

Qualifier(me) returns Position from GccEnt
is static;

IsUnqualified(me) returns Boolean from Standard
is static;
    	---Purpose: Returns true if the solution is unqualified and false in the 
    	--          other cases.

IsEnclosing(me) returns Boolean from Standard
is static;
    	---Purpose: Returns true if the solution is Enclosing the Curv and false in 
    	--          the other cases.

IsEnclosed(me) returns Boolean from Standard
is static;
    	---Purpose: Returns true if the solution is Enclosed in the Curv and false in 
    	--          the other cases.

IsOutside(me) returns Boolean from Standard
is static;
    	---Purpose: Returns true if the solution is Outside the Curv and false in 
    	--          the other cases.

fields

TheQualifier : Position from GccEnt;
TheQualified : TheCurve;

-- friends

-- Unqualified(Obj : Curv2d) from GccEnt,
-- Enclosing  (Obj : Curv2d) from GccEnt,
-- Enclosed   (Obj : Curv2d) from GccEnt,
-- Outside    (Obj : Curv2d) from GccEnt

end QualifiedCurv;


