-- Created on: 1993-01-09
-- Created by: CKY / Contract Toubro-Larsen ( Kiran )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Point from IGESGeom  inherits IGESEntity

        ---Purpose: defines IGESPoint, Type <116> Form <0>
        --          in package IGESGeom

uses

        SubfigureDef from IGESBasic,
        Pnt          from gp,
        XYZ          from gp
is

        Create returns mutable Point;

        -- Specific Methods pertaining to the class

        Init (me : mutable; aPoint : XYZ; aSymbol : SubfigureDef);
        ---Purpose : This method is used to set the fields of the class Point
        --       - aPoint  : Coordinates of point
        --       - aSymbol : SubfigureDefinition entity specifying the
        --                   display symbol if there exists one, or zero

        Value (me) returns Pnt;
        ---Purpose : returns co-ordinates of the point

        TransformedValue (me) returns Pnt;
        ---Purpose : returns co-ordinates of the point after applying Transf. Matrix

        HasDisplaySymbol (me) returns Boolean;
        ---Purpose : returns True if symbol exists

        DisplaySymbol (me) returns SubfigureDef;
        ---Purpose : returns display symbol entity if it exists

fields

--
-- Class    : IGESGeom_Point
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class Point.
--
-- Reminder : A Point instance is defined by :
--            The coordinates of the point and display symbol if any

        thePoint  : XYZ;
        theSymbol : SubfigureDef;

end Point;
