-- Created on: 1993-04-07
-- Created by: Christian CAILLET
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MultipleBinder  from Transfer  inherits Binder

    ---Purpose : Allows direct binding between a starting Object and the Result
    --           of its transfer, when it can be made of several Transient
    --           Objects. Compared to a Transcriptor, it has no Transfer Action
    --           
    --           Result is a list of Transient Results. Unique Result is not
    --           available : SetResult is redefined to start the list on the
    --           first call, and refuse the other times.
    --           
    --           rr
    --           
    --           Remark : MultipleBinder itself is intended to be created and
    --           filled by TransferProcess itself (method Bind). In particular,
    --           conflicts between Unique (Standard) result and Multiple result
    --           are avoided through management made by TransferProcess.
    --           
    --           Also, a Transcriptor (with an effective Transfer Method) which
    --           can produce a Multiple Result, may be defined as a sub-class
    --           of MultipleBinder by redefining method Transfer.

uses CString, Transient, Type, HSequenceOfTransient from TColStd

raises TransferFailure, OutOfRange

is

    Create returns MultipleBinder;
    ---Purpose : normal standard constructor, creates an empty MultipleBinder

    IsMultiple (me) returns Boolean  is redefined;
    ---Purpose : Returns True if a starting object is bound with SEVERAL
    --           results : Here, returns allways True

    ResultType (me) returns Type;
    ---Purpose : Returns the Type permitted for Results, i.e. here Transient

    ResultTypeName (me) returns CString;
    ---Purpose : Returns the Name of the Type which characterizes the Result
    --           Here, returns "(list)"


    AddResult (me : mutable; res : Transient);
    ---Purpose : Adds a new Item to the Multiple Result

    NbResults (me) returns Integer;
    ---Purpose : Returns the actual count of recorded (Transient) results

    ResultValue (me; num : Integer) returns Transient
    ---Purpose : Returns the value of the recorded result n0 <num>
    	raises OutOfRange;
    --           Error if <num> is out of range

    MultipleResult (me) returns  HSequenceOfTransient from TColStd;
    ---Purpose : Returns the Multiple Result, if it is defined (at least one
    --           Item). Else, returns a Null Handle

    SetMultipleResult (me : mutable;
    	    	       mulres : HSequenceOfTransient from TColStd)
    	raises TransferFailure;
    ---Purpose : Defines a Binding with a Multiple Result, given as a Sequence
    --           Error if a Unique Result has yet been defined

fields

    themulres : HSequenceOfTransient from TColStd;

end MultipleBinder;
