-- Created on: 1995-03-21
-- Created by: Laurent BOURESCHE
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Regul from ChFiDS 

	---Purpose: Storage of  a curve  and its 2 faces or surfaces of  support.

is

    Create returns Regul from ChFiDS;
    
    SetCurve(me : in out; IC : Integer from Standard)
    is static;
    
    SetS1(me     : in out; 
    	  IS1    : Integer from Standard;
	  IsFace : Boolean from Standard = Standard_True)
    is static;
	  
    SetS2(me     : in out; 
    	  IS2    : Integer from Standard;
	  IsFace : Boolean from Standard = Standard_True)
    is static;
	  
    IsSurface1(me) returns Boolean from Standard is static;

    IsSurface2(me) returns Boolean from Standard is static;
    
    Curve(me) returns Integer from Standard is static;

    S1(me) returns Integer from Standard is static;

    S2(me) returns Integer from Standard is static;

fields

    icurv : Integer from Standard;
    is1   : Integer from Standard;
    is2   : Integer from Standard;

end Regul;
