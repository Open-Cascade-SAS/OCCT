-- Created on: 1995-12-01
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class DrawableC2D from TestTopOpeDraw inherits Curve2d from DrawTrSurf

uses  

    Interpretor from Draw,
    Curve from Geom2d,
    Color from Draw,
    Display from Draw,
    Text2D from Draw,
    CString from Standard,
    Pnt2d from gp

is

    Create (C : Curve from Geom2d; CColor : Color from Draw)
    returns mutable DrawableC2D from TestTopOpeDraw;

    Create (C : Curve from Geom2d; CColor : Color from Draw;
    	    Text : CString; TextColor : Color from Draw)
    returns mutable DrawableC2D from TestTopOpeDraw;

    Create (C : Curve from Geom2d; CColor : Color from Draw;
    	    Text : CString; TextColor : Color from Draw;
    	    Discret : Integer;
    	    DispOrigin : Boolean = Standard_True;
            DispCurvRadius : Boolean = Standard_False;
	    RadiusMax : Real = 1.0e3;
	    RatioOfRadius : Real = 0.1)
    returns mutable DrawableC2D from TestTopOpeDraw;

    Pnt2d(me) returns Pnt2d from gp is virtual;
    
    ChangePnt2d(me : mutable; P : Pnt2d);
    
    ChangeCurve(me : mutable; C : Curve from Geom2d);
    
    ChangeText(me : mutable; T : CString from Standard);
    
    Name(me : mutable; N : CString) is redefined;
    
    Whatis(me; I : in out Interpretor from Draw) is redefined;
    ---Purpose: For variable whatis command.

    DrawOn(me; dis : in out Display from Draw) is redefined;
    
fields

    myText2D : Text2D from Draw is protected;
    myText : CString from Standard is protected;
    myTextColor : Color from Draw;

end DrawableC2D;
