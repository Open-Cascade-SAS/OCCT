-- Created on: 1993-07-12
-- Created by: Yves FRICAUD
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



deferred class SketchExplorer from MAT2d

	---Purpose: SketchExplorer  is  an iterator on  a  sketch.   A
	--          sketch is a set of contours, each contour is a set
	--          of curves from Geom2d.

uses

    Curve           from Geom2d
is
    
    NumberOfContours(me)
	--- Purpose : Returns the number of contours in the figure.
    returns Integer;
       
    Init(me : in out ; ContourIndex : Integer );
	--- Purpose : Initializes the curves explorer on the contour
	--            of range <ContourIndex>.           
   
    More(me) returns Boolean from Standard;
       	--- Purpose: Returns False if  there is no  more curves on the
       	--           current contour.
    
    Next(me : in out);
	--- Purpose  : Moves to the next curve of the current contour.
    
    Value(me) returns Curve from Geom2d; 
        --- Purpose : Returns the current curve on the current contour.
    

end SketchExplorer;




