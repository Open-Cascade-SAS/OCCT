-- File:	AppParCurves_MLineTool.cdl
-- Created:	Wed Jan 20 16:22:17 1993
-- Author:	Laurent PAINNOT
--		<lpa@sdsun1>
---Copyright:	 Matra Datavision 1993



deferred generic class MLineTool from AppParCurves (MLine  as any)

    ---Purpose: Template which defines all the services relative to
    --          a MultiLine for approximation algorithms.


uses Pnt           from gp,
     Pnt2d         from gp,
     Vec           from gp,
     Vec2d         from gp,
     Array1OfPnt   from TColgp,
     Array1OfPnt2d from TColgp,
     Array1OfVec   from TColgp,
     Array1OfVec2d from TColgp

is
    
    
    FirstPoint(myclass; ML: MLine) returns Integer;
    	---Purpose: Returns the first index of multipoints of the MLine.


    LastPoint(myclass; ML: MLine) returns Integer;
    	---Purpose: Returns the last index of multipoints of the MLine.



    NbP2d(myclass; ML: MLine) returns Integer;
    	---Purpose: Returns the number of 2d points of a MLine.


    NbP3d(myclass; ML: MLine) returns Integer;
    	---Purpose: Returns the number of 3d points of a MLine.



    Value(myclass; ML: MLine; MPointIndex: Integer; tabPt: out Array1OfPnt);
    	---Purpose: returns the 3d points of the multipoint <MPointIndex>
    	--          when only 3d points exist.


    Value(myclass; ML: MLine; MPointIndex: Integer; 
          tabPt2d: out Array1OfPnt2d);
    	---Purpose: returns the 2d points of the multipoint <MPointIndex>
    	--          when only 2d points exist.


    Value(myclass; ML: MLine; MPointIndex: Integer; 
          tabPt: out Array1OfPnt; tabPt2d: out Array1OfPnt2d);
    	---Purpose: returns the 3d and 2d points of the multipoint 
    	--          <MPointIndex>.


    Tangency(myclass; ML: MLine; MPointIndex: Integer; tabV: out Array1OfVec)
    returns Boolean;
    	---Purpose: returns the 3d points of the multipoint <MPointIndex>
    	--          when only 3d points exist.


    Tangency(myclass; ML: MLine; MPointIndex: Integer; 
          tabV2d: out Array1OfVec2d)
    returns Boolean;
    	---Purpose: returns the 2d tangency points of the multipoint 
    	--          <MPointIndex> only when 2d points exist.


    Tangency(myclass; ML: MLine; MPointIndex: Integer; 
             tabV: out Array1OfVec; tabV2d: out Array1OfVec2d)
    returns Boolean;
    	---Purpose: returns the 3d and 2d points of the multipoint 
    	--          <MPointIndex>.





end MLineTool;    
