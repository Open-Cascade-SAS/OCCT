-- Created on: 1998-04-09
-- Created by: Andre LIEUTIER
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class NLPlate from NLPlate
---Purpose: 
--
--       

uses 
     XY from gp,
     XYZ from gp, 
     StackOfPlate  from  NLPlate,
     HGPPConstraint  from  NLPlate,
     SequenceOfHGPPConstraint from  NLPlate, 
     Shape   from GeomAbs,
     Surface  from  Geom
is

    Create(InitialSurface  :  Surface  from  Geom) returns NLPlate;
-- 
-- Geometric Constraints
-- 
    Load (me : in out;  GConst : HGPPConstraint);

    Solve(me : in out; ord : Integer = 2;  InitialConsraintOrder  :  Integer=1);

    Solve2(me : in out; ord : Integer = 2;  InitialConsraintOrder  :  Integer=1);

    IncrementalSolve(me : in out; ord : Integer = 2;  InitialConsraintOrder  :  Integer=1; 
    	NbIncrements  :  Integer  =  4;  UVSliding  :  Boolean  =  Standard_False);

    IsDone(me)
        ---Purpose: returns True if all has been correctly done.
    returns Boolean;

    destroy(me : in out);
     ---C++: alias ~
 
    
    Init(me: in out );
    	---Purpose: reset the Plate in the initial state
    	--           ( same as after Create((Surface))
    
    Evaluate(me ; point2d : XY from gp )  
    returns XYZ from gp ; 
    
    EvaluateDerivative(me; point2d: XY  from gp;  
                       iu,iv  : Integer)  
    returns XYZ from gp ; 
         
    Continuity(me)  returns  Integer;

        -- private methods :
    Iterate(me : in out;  
        ConstraintOrder,  ResolutionOrder  :Integer; 
    	IncrementalLoading  : Real  =  1.0) returns Boolean
    is  private;  
     
    ConstraintsSliding(me : in out;  NbIterations  :  Integer  =  3);
    
    MaxActiveConstraintOrder(me) returns Integer;
    
    

fields 
    myInitialSurface  :  Surface  from  Geom;
    myHGPPConstraints : SequenceOfHGPPConstraint; 
    mySOP  :  StackOfPlate;
    OK : Boolean;
end;


