-- Created by: DAUTRY Philippe
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

--      	--------

---Version:	0.0
--Version	Date		Purpose
--		0.0	Feb  5 1997	Creation


package TDF 

	---Purpose: This package provides data framework for binding
	--          features and data structures.
	--          
	--          The feature structure is a tree used to bind
	--          semantic informations about each feature together.
	--          
	--          The only one concrete   attribute defined in  this
	--           package is the TagSource attribute.This attribute
	--          is used for  random creation of child labels under
	--          a given label. Tags are randomly delivered.
  
    	---Category: GUID - AttributeID
    	--           2a96b611-ec8b-11d0-bee7-080009dc3333	TDataStd_TagSource


uses

    Standard,
    MMgt,
    TColStd,
    TCollection

is


    ---Category: DF Structure Classes
    --           ==============================================================

    class Data;

    class Label;

    imported HAllocator;
    imported LabelNode;
    
    pointer LabelNodePtr to LabelNode from TDF;

    deferred class Attribute;

    class TagSource;

    class Reference;



    ---Category: DF Copy algorithms
    --           ==============================================================
    
    class ClosureMode;

    class ClosureTool;

    class CopyTool;

    class CopyLabel; 

    class ComparisonTool;

    ---Category: DF Transaction & Delta
    --           ==============================================================

    class Transaction;

    class Delta;

    deferred class AttributeDelta;

    class DeltaOnAddition;

    class DeltaOnForget;

    class DeltaOnResume;

    deferred class DeltaOnRemoval;

    deferred class DeltaOnModification;

    class DefaultDeltaOnRemoval;

    class DefaultDeltaOnModification;


    ---Category: DF Basic Tools
    --           ==============================================================

    class ChildIterator;

    class ChildIDIterator;

    imported AttributeIterator;

    ---Category: DF Specific Tools
    --           ==============================================================

    class DataSet;

    class RelocationTable;

    class Tool;

    class LabelMapHasher;

    class IDFilter;


    ---Category: DF Classes Instantiations
    --           ==============================================================

    -- Lists
    -- -----

    imported IDList;

    imported ListIteratorOfIDList;

    imported AttributeList;

    imported ListIteratorOfAttributeList;

    imported LabelList;

    imported ListIteratorOfLabelList;

    imported AttributeDeltaList;

    imported ListIteratorOfAttributeDeltaList;

    imported DeltaList;

    imported ListIteratorOfDeltaList;


    -- Sequences
    -- ---------

    imported AttributeSequence;

    imported LabelSequence;

    -- Arrays
    -- ------

    imported AttributeArray1;

    imported transient class HAttributeArray1;



    -- Maps
    -- ----

    imported IDMap;

    imported MapIteratorOfIDMap;

    imported AttributeMap;

    imported MapIteratorOfAttributeMap;

    imported AttributeDataMap;

    imported DataMapIteratorOfAttributeDataMap;

    imported AttributeDoubleMap;

    imported DoubleMapIteratorOfAttributeDoubleMap;

    imported AttributeIndexedMap;


    imported LabelMap;


    imported MapIteratorOfLabelMap;

    imported LabelDataMap;

    imported DataMapIteratorOfLabelDataMap;

    imported LabelDoubleMap;

    imported DoubleMapIteratorOfLabelDoubleMap;

    imported LabelIndexedMap;

    imported LabelIntegerMap;

    imported DataMapIteratorOfLabelIntegerMap;

    imported GUIDProgIDMap;

    imported DoubleMapIteratorOfGUIDProgIDMap;

    ---Category: Package methods
    --           ==============================================================

    LowestID returns GUID from Standard;
	---Purpose: Returns ID "00000000-0000-0000-0000-000000000000",
	--          sometimes used as null ID.
	--          
	---C++: return const &

    UppestID returns GUID from Standard;
	---Purpose: Returns ID "ffffffff-ffff-ffff-ffff-ffffffffffff".
	--          
	---C++: return const &


    AddLinkGUIDToProgID( ID : GUID from Standard; ProgID : ExtendedString from TCollection );
      ---Purpose: Sets link between GUID and ProgID in hidden DataMap
      
    GUIDFromProgID( ProgID : ExtendedString from TCollection; ID : in out GUID from Standard )
    returns Boolean from Standard;
	---Purpose: Returns True if there is GUID for given <ProgID> then GUID is returned in <ID>
	
    
    ProgIDFromGUID( ID : GUID from Standard; ProgID : in out ExtendedString from TCollection ) 	
    returns Boolean from Standard;
	---Purpose: Returns True if there is ProgID for given <ID> then ProgID is returned in <ProgID>
    
   
end TDF;
