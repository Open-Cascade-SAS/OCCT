-- Created on: 1996-07-08
-- Created by: Christian CAILLET
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Reader  from STEPControl inherits Reader from XSControl

	---Purpose : Reads STEP files, checks them and translates their contents
    	-- into Open CASCADE models. The STEP data can be that of
    	-- a whole model or that of a specific list of entities in the model.
    	-- As in XSControl_Reader, you specify the list using a selection.
    	-- For the translation of iges files it is possible to use next sequence:
     	-- To change translation parameters 
    	-- class Interface_Static should be used before beginning of
    	-- translation  (see STEP Parameters and General Parameters) 
    	--     Creation of reader - STEPControl_Reader reader;
    	--  To load s file in a model use method reader.ReadFile("filename.stp")
    	-- To print load results reader.PrintCheckLoad(failsonly,mode)
    	-- where mode is equal to the value of enumeration IFSelect_PrintCount 
    	--   For definition number of candidates :
    	-- Standard_Integer nbroots = reader. NbRootsForTransfer();
    	-- To transfer entities from a model the following methods can be used:
    	-- for the whole model - reader.TransferRoots(); 
    	-- to transfer a list of entities: reader.TransferList(list);
    	-- to transfer one entity Handle(Standard_Transient)
    	-- ent = reader.RootForTransfer(num);
    	-- reader.TransferEntity(ent), or 
    	-- reader.TransferOneRoot(num), or
    	-- reader.TransferOne(num), or 
    	-- reader.TransferRoot(num)
    	--   To obtain the result the following method can be used:
    	-- reader.NbShapes() and reader.Shape(num); or reader.OneShape(); 
    	-- To print the results of transfer use method:
    	-- reader.PrintCheckTransfer(failwarn,mode);
    	-- where printfail is equal to the value of enumeration
    	-- IFSelect_PrintFail, mode see above; or reader.PrintStatsTransfer();
    	-- Gets correspondence between a STEP entity and a result
    	-- shape obtained from it.
    	-- Handle(XSControl_WorkSession)
    	-- WS = reader.WS();
    	-- if ( WS->TransferReader()->HasResult(ent) )
    	-- TopoDS_Shape shape = WS->TransferReader()->ShapeResult(ent);

uses

    CString, OStream, Transient, SequenceOfTransient from TColStd,
    StepModel from StepData, WorkSession from XSControl,
    ReturnStatus from IFSelect, PrintCount from IFSelect,
    Shape from TopoDS, SequenceOfShape from TopTools,
    SequenceOfAsciiString from TColStd,
    Array1OfAsciiString from TColStd,
    Array1OfReal from TColStd,
    SequenceOfAsciiString from TColStd,
    RepresentationContext from StepRepr
is

    Create returns Reader;
    ---Purpose : Creates a reader object with an empty STEP model.

    Create (WS : mutable WorkSession from XSControl;
    	    	 scratch : Boolean = Standard_True) returns Reader;
    ---Purpose : Creates a Reader for STEP from an already existing Session
    --           Clears the session if it was not yet set for STEP

    StepModel (me) returns StepModel;
    ---Purpose : Returns the model as a StepModel.
    --           It can then be consulted (header, product)

    TransferRoot (me : in out; num : Integer = 1) returns Boolean;
    ---Purpose : Transfers a root given its rank in the list of candidate roots
    --           Default is the first one
    --           Returns True if a shape has resulted, false else
    --           Same as inherited TransferOneRoot, kept for compatibility

    NbRootsForTransfer (me : in out) returns Integer is redefined;
    ---Purpose : Determines the list of root entities from Model which are candidate for
    --           a transfer to a Shape (type of entities is PRODUCT)
    
    FileUnits(me : in out; theUnitLengthNames : in out SequenceOfAsciiString from TColStd;
    	    	  theUnitAngleNames : in out SequenceOfAsciiString from TColStd;
    	    	  theUnitSolidAngleNames : in out SequenceOfAsciiString from TColStd );
     ---Purpose : Returns sequence of all unit names for shape representations 
     --           found in file
     
    findUnits(me : in out ; theReprContext : RepresentationContext from StepRepr;
     	theNameUnits : in out Array1OfAsciiString from TColStd;
     	theFactorUnits : in out Array1OfReal from TColStd) returns Boolean is private;
     ---Purpose : Returns  units for length , angle and solidangle for shape representations 
    
    
end Reader;
