-- File:        SweptAreaSolid.cdl
-- Created:     Mon Dec  4 12:02:32 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWSweptAreaSolid from RWStepShape

	---Purpose : Read & Write Module for SweptAreaSolid

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     SweptAreaSolid from StepShape,
     EntityIterator from Interface

is

	Create returns RWSweptAreaSolid;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable SweptAreaSolid from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : SweptAreaSolid from StepShape);

	Share(me; ent : SweptAreaSolid from StepShape; iter : in out EntityIterator);

end RWSweptAreaSolid;
