-- Created on: 1994-09-23
-- Created by: Yves FRICAUD
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class CutCurve from MAT2d 

	---Purpose: Cuts a curve at the extremas of curvature
	--          and at the inflections. Constructs a trimmed
	--          Curve for each interval.

uses
    Curve           from Geom2d,
    TrimmedCurve    from Geom2d,
    SequenceOfCurve from TColGeom2d,
    Side            from MAT
    
raises 
    OutOfRange from Standard
    
is
    Create;
    
    Create  (C : Curve from Geom2d) returns CutCurve from MAT2d;
    
    Perform (me : in out; C : Curve from Geom2d) 	    
	---Purpose: Cuts a curve at the extremas of curvature
	--          and at the inflections.
    is static;
    
    Perform (me : in out; C : Curve from Geom2d; aSide : Side from MAT)
    	---Purpose: Cuts a curve at the inflections, and at the extremas
    	--          of curvature where the concavity is on <aSide>. 
    is static;
    
    PerformInf (me : in out; C : Curve from Geom2d)    	
    	---Purpose: Cuts a curve at the inflections.
    is static;
    
    UnModified (me) returns Boolean from Standard
    	---Purpose: Returns True if the curve is not cut.
    is static;
    

    NbCurves (me) returns Integer from Standard
    	---Purpose: Returns the number of curves.
    	--          it's allways greatest than 2.    
    	--          
    	raises
    	    OutOfRange from Standard
	    ---Purpose: raises if the Curve is UnModified;        
    is static;
    

    Value (me ; Index : Integer from Standard) returns TrimmedCurve from Geom2d
	---Purpose: Returns the Indexth curve.    
        raises
    	    OutOfRange from Standard
	    ---Purpose: raises if Index not in the range [1,NbCurves()]
    is static;

    
fields
    theCurves : SequenceOfCurve from TColGeom2d;
    
end CutCurve;
