-- Created on: 1991-05-23
-- Created by: Didier PIFFAULT
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package Intf 

	---Purpose: Interference computation  between polygons, lines  and
	--          polyhedra with only  triangular  facets. These objects
	--          are polygonal  representations of complex   curves and
	--          triangulated representations of complex surfaces.


uses Standard, TCollection, TColStd, gp, Bnd, IntAna2d


is

--  Enumeration :

    enumeration PIType is EXTERNAL, FACE, EDGE, VERTEX;
    ---Purpose: Describes the different intersection  point types for this
    --          application.


--  Classes input data :

    deferred class Polygon2d;

    class Array1OfLin instantiates Array1 from TCollection
     	    	    (Lin from gp);
    ---Purpose: Describes  a set of Straight Lines  to  intersect with the
    --          Polyhedron.



--	Classes output data :

    class SectionPoint;

    class SeqOfSectionPoint instantiates Sequence from TCollection
    	    	    	    	    	    (SectionPoint);


    class SectionLine;

    class SeqOfSectionLine instantiates Sequence from TCollection
    	    	    	    	    	    (SectionLine);


    class TangentZone;

    class SeqOfTangentZone instantiates Sequence from TCollection
    	    	    	    	    	    (TangentZone);


    deferred class Interference;

-- Algorithms :

    class Tool;


    class InterferencePolygon2d;
    ---Purpose: Computes   the  interference between   two polygons in  2d.
    --          Result : points of intersections and zones of tangence.

    generic class InterferencePolygonPolyhedron;
    ---Purpose: Computes the interference  between a polygon or  a straight
    --          line and a polyhedron.   Points of intersection  and zones
    --          of tangence.


    --- Package Methods :
    --  

    PlaneEquation  (P1            : in Pnt from gp;
		    P2            : in Pnt from gp;
		    P3            : in Pnt from gp;
		    NormalVector  : out XYZ from gp;
		    PolarDistance : out Real from Standard);
    ---Purpose: Give the plane equation of the triangle <P1> <P2> <P3>.


    Contain	   (P1            : in Pnt from gp;
		    P2            : in Pnt from gp;
		    P3            : in Pnt from gp;
		    ThePnt	  : in Pnt from gp)
		    returns Boolean;
    ---Purpose: Compute if the triangle <P1> <P2> <P3> contain <ThePnt>.


end Intf;
