-- Created on: 1993-09-14
-- Created by: Jean-Louis FRENKEL
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Text from Prs3d inherits Root from Prs3d

    	--- Purpose: A framework to define the display of texts.
uses
    Presentation from Prs3d,
    Pnt from gp,
    Drawer from Prs3d,
    TextAspect from Prs3d,
    ExtendedString from TCollection
    
is
    Draw(myclass; aPresentation: Presentation from Prs3d;
    	          aDrawer: Drawer from Prs3d;
		  aText: ExtendedString from TCollection;
                  AttachmentPoint: Pnt from gp);
    	---Purpose: Defines the display of the text aText at the point AttachmentPoint.
    	-- The drawer aDrawer specifies the display attributes which texts will have.
    	-- The presentation object aPresentation stores the
    	-- information defined in this framework.
    	-- static void Draw (const Handle(Prs3d_Presentation)&
    	-- aPresentation, const Handle(Prs3d_TextAspect)&
    	-- anAspect, const TCollection_ExtendedString& aText,
    	-- const gp_Pnt& AttachmentPoint);    

    Draw(myclass; aPresentation: Presentation from Prs3d;
    	          anAspect: TextAspect from Prs3d;
		  aText: ExtendedString from TCollection;
                  AttachmentPoint: Pnt from gp);
    
    	---Purpose: Defines the display of the text aText at the point
    	-- AttachmentPoint.
    	-- The text aspect object anAspect specifies the display
    	-- attributes which texts will have.
	-- The presentation object aPresentation stores the
    	-- information defined in this framework.
    	-- This syntax could be used if you had not already
    	-- defined text display attributes in a drawer or if you
    	-- wanted to exceptionally overide the definition
    	-- provided in your drawer.    
		  
end Text from Prs3d;
