-- Created by: Peter KURNEV
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Pave from BOPDS  

	---Purpose: 
    	-- The class BOPDS_Pave is to store  
    	-- information about vertex on an edge 
--uses
--raises

is 
    Create 
    	returns Pave from BOPDS; 
    ---C++: alias "Standard_EXPORT virtual ~BOPDS_Pave();"   
    ---C++: inline  
    	---Purpose:  
    	--- Empty contructor  
    	---  
     
    SetIndex(me:out;  
    	    theIndex: Integer from Standard); 
    ---C++: inline    
    	---Purpose:   
	--- Modifier   
	--- Sets the index of vertex <theIndex>
	
    Index(me)  
    	returns Integer from Standard; 
    ---C++: inline  
     	---Purpose: 
    	--- Selector   
	--- Returns the index of vertex 
    SetParameter(me:out;  
    	    theParameter: Real from Standard); 
    ---C++: inline      
     	---Purpose:   
	--- Modifier   
	--- Sets the parameter of vertex <theParameter> 
	
    Parameter(me)  
    	returns Real from Standard; 
    ---C++: inline     	
    	---Purpose: 
    	--- Selector   
	--- Returns the parameter of vertex
    Contents(me; 
    	    theIndex:out Integer from Standard; 
	    theParameter:out Real from Standard); 
    ---C++: inline 
       	---Purpose: 
    	--- Selector  
    	--- Returns the index of vertex <theIndex>  
	--- Returns the parameter of vertex <theParameter> 
	
    IsLess(me; 
    	    theOther:  Pave from BOPDS) 
    	returns Boolean from Standard;  
    ---C++: alias operator <	 
    ---C++: inline  
    	---Purpose: 
    	--- Query  
    	--- Returns true if thr parameter od this is less   
    	--  than the parameter of  <theOther> 
    
    IsEqual(me; 
    	    theOther:  Pave from BOPDS) 
    	returns Boolean from Standard;  
    ---C++: alias operator == 
    ---C++: inline  
     	---Purpose: 
    	--- Query  
    	--- Returns true if thr parameter od this is equal   
    	--  to the parameter of  <theOther> 
	 
    Dump(me); 

fields 
    myIndex    : Integer from Standard is protected;     
    myParameter: Real from Standard is protected;     

end Pave;
