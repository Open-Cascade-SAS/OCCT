-- File:        SurfaceStyleUsage.cdl
-- Created:     Fri Dec  1 11:11:28 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class SurfaceStyleUsage from StepVisual 

inherits TShared from MMgt

uses

	SurfaceSide from StepVisual, 
	SurfaceSideStyle from StepVisual
is

	Create returns mutable SurfaceStyleUsage;
	---Purpose: Returns a SurfaceStyleUsage

	Init (me : mutable;
	      aSide : SurfaceSide from StepVisual;
	      aStyle : mutable SurfaceSideStyle from StepVisual) is virtual;

	-- Specific Methods for Field Data Access --

	SetSide(me : mutable; aSide : SurfaceSide);
	Side (me) returns SurfaceSide;
	SetStyle(me : mutable; aStyle : mutable SurfaceSideStyle);
	Style (me) returns mutable SurfaceSideStyle;

fields

	side : SurfaceSide from StepVisual; -- an Enumeration
	style : SurfaceSideStyle from StepVisual;

end SurfaceStyleUsage;
