-- Created on: 1993-07-08
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class BoxSort from TopOpeBRepTool

uses

    Box from Bnd,
    BoundSortBox from Bnd,
    HArray1OfBox from Bnd,
    HArray1OfInteger from TColStd,
    ListOfInteger from TColStd,
    ListIteratorOfListOfInteger from TColStd,
    ShapeEnum from TopAbs,
    Shape from TopoDS,
    IndexedMapOfShape from TopTools,
    Box from Bnd,
    HBoxTool from TopOpeBRepTool
    
is

    Create returns BoxSort;
    Create(T:HBoxTool) returns BoxSort;
    SetHBoxTool(me:in out;T:HBoxTool);
    HBoxTool(me) returns HBoxTool;---C++: return const &
    Clear(me:in out);
    AddBoxes(me:in out;S:Shape;TS:ShapeEnum;TA:ShapeEnum=TopAbs_SHAPE);
    MakeHAB(me:in out;S:Shape;TS:ShapeEnum;TA:ShapeEnum=TopAbs_SHAPE);
    HAB(me) returns HArray1OfBox from Bnd;---C++:return const &
    MakeHABCOB(myclass;HAB:HArray1OfBox from Bnd;COB:out Box from Bnd);
    HABShape(me; I:Integer) returns Shape;---C++: return const &
    MakeCOB(me:in out;S:Shape;TS:ShapeEnum;TA:ShapeEnum=TopAbs_SHAPE);
    AddBoxesMakeCOB(me:in out;S:Shape;TS:ShapeEnum;TA:ShapeEnum=TopAbs_SHAPE);
    Compare(me:out;S:Shape) returns ListIteratorOfListOfInteger;---C++:return const&
    TouchedShape(me;I:ListIteratorOfListOfInteger) returns Shape;---C++:return const&
    Box(me;S:Shape) returns Box from Bnd;---C++:return const & 
    
--modified by NIZNHY-PKV Mon Dec 16 10:24:42 2002  f
    Destroy(me: out); 
    ---C++:  alias  "Standard_EXPORT ~TopOpeBRepTool_BoxSort() {Destroy();}"
--modified by NIZNHY-PKV Mon Dec 16 10:25:22 2002  t

fields

    myCOB:Box from Bnd;
    myBSB:BoundSortBox from Bnd;
    myIterator:ListIteratorOfListOfInteger from TColStd;
    myLastCompareShape:Shape from TopoDS;
    myLastCompareShapeBox:Box from Bnd;
    myHBT:HBoxTool from TopOpeBRepTool;
    myHAB:HArray1OfBox from Bnd;
    myHAI:HArray1OfInteger from TColStd;    

end BoxSort;
