-- File:	BRepPrimAPI_MakeOneAxis.cdl
-- Created:	Thu Jul 22 15:13:07 1993
-- Author:	Remi LEQUETTE
--		<rle@nonox>
---Copyright:	 Matra Datavision 1993


deferred class MakeOneAxis from BRepPrimAPI inherits MakeShape from BRepBuilderAPI

	---Purpose: The abstract class MakeOneAxis is the root class of
    	-- algorithms used to construct rotational primitives.

uses
    Address from Standard,
    Face    from TopoDS,
    Shell   from TopoDS,
    Solid   from TopoDS

raises
    NotDone     from StdFail

is
    OneAxis(me : in out) returns Address from Standard
	---Purpose: The inherited commands should provide the algorithm.
	--          Returned as a pointer.
	---Level: Public
    is deferred;
    
    Build(me : in out)
	---Purpose: Stores the solid in myShape.
	---Level: Public
    is redefined;

    Face(me : in out) 
	---Purpose: Returns the lateral face of the rotational primitive.
	--          
	---C++: return const &
	---C++: alias "Standard_EXPORT operator TopoDS_Face();" 
	---Level: Public
    returns Face from TopoDS
    is static;

    Shell(me : in out) 
	---Purpose: Returns the constructed rotational primitive as a shell.
    	---C++: return const &
	---C++: alias "Standard_EXPORT operator TopoDS_Shell();" 
    returns Shell from TopoDS
    is static;

    Solid(me : in out) 
	---Purpose: Returns the constructed rotational primitive as a solid.
	---C++: return const &
	---C++: alias "Standard_EXPORT operator TopoDS_Solid();" 
    returns Solid from TopoDS 
    is static;


end MakeOneAxis;
