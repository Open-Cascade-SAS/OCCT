-- Created on: 1995-01-25
-- Created by: Jean-Louis Frenkel
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Modified by  Rob (18/12/96) -> information about modes to update.
--              Rob (04/07/97) ->   TypeOfPresentation3d () Method 
--                                  changed to Public Method.
--                             -> Option Projector Dependant/Independant
--                                may be set at any time , not only in
--                                the constructor or the presentable.
--                               ->Insert Locations Methods...
--              Rob (16/12/97) -> Get the list of modes to be updated
--                             -> Flags all the Prs to be updated...                 

deferred class PresentableObject from PrsMgr inherits TShared from MMgt


    	---Purpose: A framework to supply the Graphic3d
    	-- structure of the object to be presented. On the first
    	-- display request, this structure is created by calling the
    	-- appropriate algorithm and retaining this frameworkfor
    	-- further display.
    	-- This abstract framework is inherited in Application
    	-- Interactive Services (AIS), notably in:
    	-- -   AIS_InteractiveObject
    	-- -   AIS_ConnectedInteractive
    	-- -   AIS_MultipleConnectedInteractive
    	-- -   AIS_Shape
    	--   Consequently, 3D presentation should be handled by
    	-- the relevant daughter classes and their member
    	-- functions in AIS. This is particularly true in the
    	-- creation of new interactive objects.

uses
    Presentation           from PrsMgr,
    Presentation           from Prs3d,
    Presentations          from PrsMgr,
    PresentationManager    from PrsMgr,
    PresentationManager3d  from PrsMgr,
    TypeOfPresentation3d   from PrsMgr,
    ListOfPresentableObjects from PrsMgr,
    PresentableObjectPointer from PrsMgr,
    DataStructureManager   from Graphic3d,
    Projector              from Prs3d,
    Transformation         from Geom,
    ListOfInteger          from TColStd,
    Location               from TopLoc, 
    ClipPlane              from Graphic3d,
    SequenceOfHClipPlane   from Graphic3d,
    TransModeFlags         from Graphic3d, 
    Pnt                    from gp,
    Trsf                   from gp, 
    CTransPersStruct       from  Graphic3d,
    ZLayerId from Graphic3d

raises
    NotImplemented from Standard
is


    Initialize(aTypeOfPresentation3d: TypeOfPresentation3d from PrsMgr = PrsMgr_TOP_AllView);
      ---C++: alias "Standard_EXPORT virtual ~PrsMgr_PresentableObject();"
    
---Category: deferred methods.
--           
    
    Compute(me:mutable;
                aPresentationManager: PresentationManager3d from PrsMgr;
                aPresentation: Presentation from Prs3d;
                aMode: Integer from Standard = 0)
    	---Purpose: Calculates the 3D view aPresentation and its
    	-- updates. The latter are managed by aPresentationManager.
    	-- aPresentableObject has the display mode aMode;
    	-- this has the default value of 0, that is, the wireframe display mode.
    raises NotImplemented from Standard
    is virtual protected;
    
    Compute(me            : mutable;
            aProjector    : Projector from Prs3d;
            aPresentation  : Presentation from Prs3d)
    	---Purpose: Calculates the 3D view aPresentation and its
    	-- updates. The latter are managed by
    	-- aPresentationManager. Each of the views in the
    	-- viewer and every modification such as rotation, for
    	-- example, entails recalculation.
    	-- It must be redefined to implement hidden line removal
    	-- for the object. The user never calls this method
    	-- himself. This is done via the InteractiveContext object
    	-- and is dependent on the point of view from which the
    	-- object is displayed.
    raises NotImplemented from Standard
    is virtual protected;

    Compute(me            : mutable;
            aProjector    : Projector from Prs3d;
            aTrsf         : Transformation from Geom;
            aPresentation : Presentation from Prs3d)
    is virtual protected;
    	---Purpose: Calculates the 3D view aPresentation and its
    	-- updates. The latter are managed by
    	-- aPresentationManager. A point of view is provided
    	-- by the projector aProjector, and the geometric
    	-- transformation which has transformed associated
    	-- presentable objects is specified by aTrsf.
    	-- This function is to be used in case where a hidden
    	-- line removal display cannot be calculated
    	-- automatically. This occurs   when associated
    	-- presentable objects have been transformed
    	-- geometrically, but not translated.
    	-- Warning
    	-- The transformation aTrsf must be applied to the
    	-- object before computation.

    Update(me: mutable;AllModes: Boolean=Standard_False)
    	---Purpose: recomputes all presentations of the object.
    	---Level: Public 
    is protected;

    Update(me: mutable; aMode: Integer from Standard; ClearOther: Boolean from Standard)
    	---Purpose: Recomputes the presentation in the given mode.
    	--          If ClearOther is true, other presentation will be cleared.
    is protected;
    
    Fill(me: mutable; 
                aPresentationManager: PresentationManager from PrsMgr;
                aPresentation: Presentation from PrsMgr;
                aMode: Integer from Standard = 0)
    -- 22-03-04 OCC4895 SAN High-level interface for controlling polygon offsets
    is virtual protected;
    	--- Purpose: High-level interface for controlling polygon offsets
        
        -- 22-03-04 OCC4895 SAN High-level interface for controlling polygon offsets

    
    -- Presentations(me: mutable) returns Presentations from PrsMgr
    -- is static private;
    
    Presentations(me : mutable) returns Presentations from PrsMgr
    is static;
    	---C++: return &
            
   TypeOfPresentation3d(me) returns TypeOfPresentation3d from PrsMgr
   is static;
    	---Purpose: Returns information on whether the object accepts display in HLR mode or not.
    
   --   ABD 29/10/04  Transform Persistence of Presentation( pan, zoom, rotate ) 
   SetTransformPersistence(  me     :  mutable; 
   			     aFlag  :  TransModeFlags  from  Graphic3d; 
    	    	    	     APoint :  Pnt from gp )
   is virtual; 
   ---Level:    Public 
   ---Purpose:  Sets up Transform Persistence Mode for this object.
   -- This function used to lock in object position, rotation and / or zooming relative to camera position.
   -- Object will be drawn in the origin setted by APoint parameter (except Graphic3d_TMF_TriedronPers flag
   -- - see description later). aFlag should be:
   -- -   Graphic3d_TMF_None - no persistence attributes (reset);
   -- -   Graphic3d_TMF_PanPers - object doesn't move;
   -- -   Graphic3d_TMF_ZoomPers - object doesn't resize;
   -- -   Graphic3d_TMF_RotatePers - object doesn't rotate;
   -- -   Graphic3d_TMF_FullPers - pan, zoom and rotate transform persistence;
   -- -   Graphic3d_TMF_TriedronPers - object behaves like trihedron;
   -- -   combination (Graphic3d_TMF_PanPers | Graphic3d_TMF_ZoomPers);
   -- -   combination (Graphic3d_TMF_PanPers | Graphic3d_TMF_RotatePers);
   -- -   combination (Graphic3d_TMF_ZoomPers | Graphic3d_TMF_RotatePers).
   -- If Graphic3d_TMF_TriedronPers or Graphic3d_TMF_2d persistence mode selected APoint coordinates X and Y means:
   -- -   X = 0.0, Y = 0.0 - center of view window;
   -- -   X > 0.0, Y > 0.0 - right upper corner of view window;
   -- -   X > 0.0, Y < 0.0 - right lower corner of view window;
   -- -   X < 0.0, Y > 0.0 - left  upper corner of view window;
   -- -   X < 0.0, Y < 0.0 - left  lower corner of view window.
   -- And Z coordinate defines the gap from border of view window (except center position).
   ---Category: Graphic attributes management  
   
   SetTransformPersistence(  me     :  mutable; 
   			     aFlag  :  TransModeFlags  from  Graphic3d ) 
   is  static; 
   ---Level:    Public 
   ---Purpose:  Calls previous method  with  point  (0,0,0)
   ---Category: Graphic attributes management 
   
    
   GetTransformPersistenceMode( me )  returns  TransModeFlags  from  Graphic3d  is  static;
    
   ---Level:    Public 
   ---Purpose:  Gets  Transform  Persistence Mode  for  this  object 
   ---Category: Graphic attributes management

   GetTransformPersistencePoint( me )  returns  Pnt  from  gp  is  static;
    
   ---Level:    Public 
   ---Purpose:  Gets  point  of  transform  persistence for  this  object 
   ---Category: Graphic attributes management
    
   --   ABD 29/10/04  Transform Persistence of Presentation( pan, zoom, rotate )
    
   SetTypeOfPresentation(me:mutable; aType: TypeOfPresentation3d from PrsMgr);    

   SetToUpdate    (me:mutable;aMode:Integer from Standard);
   ---Purpose: flags the Prs of mode <AMode> to be Updated.
   --          the Update will be done when needed.
   
   SetToUpdate(me:mutable); 
   ---Purpose: flags all the Presentations to be Updated.
    
   ToBeUpdated(me;ListOfMode : out ListOfInteger from TColStd);
   ---Purpose: gives the list of modes which are flagged "to be updated".
    
   SetLocalTransformation(me:mutable; theTransformation:Trsf from gp) is virtual;
   ---Purpose: Sets local transformation to theTransformation.

   SetCombinedParentTransform(me:mutable; theTransformation:Trsf from gp) is virtual protected;
   ---Purpose: Sets myCombinedParentTransform to theTransformation. Thus object receives transformation
   -- from parent node and able to derive its own.
    
   HasTransformation(me) returns Boolean from Standard;
   ---Purpose: Returns true if object has a transformation that is different from the identity.
   
   LocalTransformation(me) returns any Trsf from gp;
   ---C++: inline
   ---C++: return const&

   Transformation(me) returns any Trsf from gp;
   ---C++: inline
   ---C++: return const&

   InversedTransformation(me) returns any Trsf from gp;
   ---C++: inline
   ---C++: return const&
   
   ResetTransformation(me:mutable)  is virtual;
   ---Purpose: resets local transformation to identity.

   UpdateTransformation(me:mutable) is virtual;
    
   UpdateTransformation(me:mutable;P : Presentation from Prs3d) is virtual;

   SetZLayer ( me         : mutable;
               theLayerId : ZLayerId from Graphic3d )
     is virtual;
   ---Purpose: Set Z layer ID and update all presentations of the presentable object.
   -- The layers mechanism allows drawing objects in higher layers in overlay of objects in lower layers.

   ZLayer ( me )
     returns ZLayerId from Graphic3d is static;
   ---Purpose: Get ID of Z layer.

   AddClipPlane (me : mutable; thePlane : ClipPlane from Graphic3d) is virtual;
   ---Purpose: Adds clip plane for graphical clipping for all display mode
   -- presentations. The composition of clip planes truncates the rendering
   -- space to convex volume. Please be aware that number of supported
   -- clip plane is limited. The planes which exceed the limit are ignored.
   -- Besides of this, some planes can be already set in view where the object
   -- is shown: the number of these planes should be substracted from limit
   -- to predict the maximum possible number of object clipping planes.
   -- @param thePlane [in] the clip plane to be appended to map of clip planes.

   RemoveClipPlane (me : mutable; thePlane : ClipPlane from Graphic3d) is virtual;
   ---Purpose: Removes previously added clip plane.
   -- @param thePlane [in] the clip plane to be removed from map of clip planes.

   SetClipPlanes (me : mutable; thePlanes : SequenceOfHClipPlane from Graphic3d) is virtual;
   ---Purpose: Set clip planes for graphical clipping for all display mode presentations.
   -- The composition of clip planes truncates the rendering space to convex
   -- volume. Please be aware that number of supported clip plane is limited.
   -- The planes which exceed the limit are ignored. Besides of this, some
   -- planes can be already set in view where the object is shown: the number 
   -- of these planes should be substracted from limit to predict the maximum
   -- possible number of object clipping planes.

   GetClipPlanes (me) returns SequenceOfHClipPlane from Graphic3d;
   ---C++: inline
   ---C++: return const&
   ---Purpose: Get clip planes.
   -- @return set of previously added clip planes for all display mode presentations.

  SetMutable ( me           : mutable;
               theIsMutable : Boolean from Standard ) is virtual;
  ---Purpose: Sets if the object has mutable nature (content or location will be changed regularly).
  -- This method should be called before object displaying to take effect.

  IsMutable (me) returns Boolean from Standard;
  ---C++: return const
  ---Purpose: Returns true if object has mutable nature (content or location are be changed regularly).
  -- Mutable object will be managed in different way than static onces (another optimizations).

  AddChild ( me           : mutable;
             theObject    : PresentableObject from PrsMgr ) is virtual;
    --- Purpose: Makes theObject child of current object in scene hierarchy. 

  RemoveChild ( me           : mutable;
                theObject    : PresentableObject from PrsMgr ) is virtual;
    --- Purpose: Removes theObject from children of current object in scene hierarchy. 

  Children (me) returns ListOfPresentableObjects from PrsMgr is static;
    ---C++: return const&
    --- Purpose: Returns children of the current object.

  HasOwnPresentations (me) returns Boolean from Standard is static;
    ---C++: return const
    --- Purpose: Returns true if object should have own presentations.

  Parent (me) returns PresentableObjectPointer from PrsMgr is static;
    ---C++: return const
    --- Purpose: Returns parent of current object in scene hierarchy.

   UpdateClipping (me : mutable) is virtual protected;
   ---Purpose: General virtual method for internal update of presentation state
   -- when some modifications on list of clip planes occurs. Base 
   -- implementation propagate clip planes to every presentation.

fields
    myPresentations: Presentations from PrsMgr is protected;
    myTypeOfPresentation3d: TypeOfPresentation3d from PrsMgr is protected;
    myClipPlanes : SequenceOfHClipPlane from Graphic3d is protected;
    myTransformPersistence  :  CTransPersStruct  from  Graphic3d;
    myIsMutable : Boolean from Standard is protected;
    myZLayer    : ZLayerId from Graphic3d is protected;

    myHasOwnPresentations : Boolean from Standard is protected; -- shows if object should have own presentations.

    myParent : PresentableObjectPointer from PrsMgr; -- Reference to parent object in scene hierarchy.
 
    myLocalTransformation : Trsf from gp;     -- Own transformation of presentable object.
    myTransformation : Trsf from gp;          -- Combined transformation of presentable object.
    myInvTransformation : Trsf from gp;       -- Inverted combined transformation of presentable object.
    myCombinedParentTransform : Trsf from gp; -- Combined transformation of presentable object excepting local transformation.

    myChildren : ListOfPresentableObjects from PrsMgr; -- Child objects in scene hierarchy.

friends
    class Presentation        from PrsMgr,
    class PresentationManager from PrsMgr,
    Compute from Presentation from PrsMgr(me : mutable; aProjector   : DataStructureManager from Graphic3d),
    Compute from Presentation from PrsMgr(me : mutable; aProjector   : DataStructureManager from Graphic3d;
                                                        aGivenStruct :  Structure from Graphic3d),
    Compute from Presentation from PrsMgr(me : mutable; aProjector   : DataStructureManager from Graphic3d;
                                                        TheTrsf   : Transformation from Geom),
    Compute from Presentation from PrsMgr(me : mutable; aProjector   : DataStructureManager from Graphic3d;
                                                        TheTrsf      : Transformation from Geom;
                                                        aGivenStruct : Structure from Graphic3d)
end PresentableObject from PrsMgr;
