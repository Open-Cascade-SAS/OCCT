-- Created on: 1995-10-23
-- Created by: Mister rmi
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class GCurve from PBRep inherits CurveRepresentation from PBRep

	---Purpose: Root   class    for    the    geometric     curves
	--          representation. Contains a range.

uses

    Location from PTopLoc,
    Pnt      from gp

is

    Initialize(L : Location from PTopLoc;
    	       First , Last : Real from Standard);

    First(me) returns Real
    is static;

    Last(me) returns Real
    is static;

    First(me : mutable; F : Real)
    is static;

    Last(me : mutable; L : Real)
    is static;

    IsGCurve(me) returns Boolean from Standard
    	---Purpose: returns TRUE
    is redefined;

fields

    myFirst    : Real;
    myLast     : Real;

end GCurve;
