-- Created on: 1994-08-24
-- Created by: Gilles DEBARBOUILLE
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class VariableGroup from Dynamic

inherits

    Variable from Dynamic
    
	---Purpose: This   inherited  class   from   variable is   for
	--          specifing  that the variable  does not accept only
	--          one   value    but a  collection   of  homogeneous
	--          values. This class is for describing the signature
	--          of the method definition. When an instance of this
	--          kind   of   method    is     done,    it   is    a
	--          CompositVariableInstance which is used.


is

    Create returns mutable VariableGroup from Dynamic;
    
    ---Level: Advanced 
    
    ---Purpose: Creates and Returns a new instance of this class.
    

end VariableGroup;
