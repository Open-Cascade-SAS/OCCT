-- Created on: 1999-09-08
-- Created by: Andrey BETENEV
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Unit from StepBasic inherits SelectType from StepData

    ---Purpose: Implements a select type unit (NamedUnit or DerivedUnit)

uses
    NamedUnit from StepBasic,
    DerivedUnit from StepBasic

is
    Create returns Unit;
    	---Purpose: Creates empty object
	
    CaseNum (me; ent : Transient) returns Integer;
	---Purpose : Recognizes a type of Unit Entity
        --        1 -> NamedUnit
        --        2 -> DerivedUnit

    NamedUnit (me) returns any NamedUnit from StepBasic;
        ---Purpose : returns Value as a NamedUnit (Null if another type)

    DerivedUnit (me) returns any DerivedUnit from StepBasic;
        ---Purpose : returns Value as a DerivedUnit (Null if another type)

end Unit;
