-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class AutoDesignGeneralOrgItem from StepAP214 inherits SelectType from StepData

	-- <AutoDesignGeneralOrgItem> is an EXPRESS Select Type construct translation.
	-- it gathers : Product, ProductDefinition, ProductDefinitionFormation, Representation

uses
     AutoDesignDocumentReference from StepAP214,
     ExternallyDefinedRepresentation from StepRepr,
     Product from StepBasic,
     ProductDefinition from StepBasic,
     ProductDefinitionFormation from StepBasic,
     ProductDefinitionRelationship from StepBasic,
     ProductDefinitionWithAssociatedDocuments from StepBasic,
     Representation from StepRepr
is

	Create returns AutoDesignGeneralOrgItem;
	---Purpose : Returns a AutoDesignGeneralOrgItem SelectType

	CaseNum (me; ent : Transient) returns Integer;
	---Purpose: Recognizes a AutoDesignGeneralOrgItem Kind Entity that is :
	-- 1     Product from StepBasic,
	-- 2     ProductDefinition from StepBasic,
	-- 3     ProductDefinitionFormation from StepBasic,
	-- 4     ProductDefinitionRelationship from StepBasic,
	-- 5     ProductDefinitionWithAssociatedDocuments from StepBasic,
	-- 6     Representation from StepRepr
	-- 7     ExternallyDefinedRepresentation from StepRepr,
	-- 8     AutoDesignDocumentReference from StepAP214,
	--        0 else

	Product (me) returns any Product;
	---Purpose : returns Value as a Product (Null if another type)

	ProductDefinition (me) returns any ProductDefinition;
	---Purpose : returns Value as a ProductDefinition (Null if another type)

	ProductDefinitionFormation (me) returns any ProductDefinitionFormation;
	---Purpose : returns Value as a ProductDefinitionFormation (Null if another type)

	ProductDefinitionRelationship (me) returns any ProductDefinitionRelationship;
	---Purpose : returns Value as a ProductDefinitionRelationship (Null if another type)

	ProductDefinitionWithAssociatedDocuments (me) returns any ProductDefinitionWithAssociatedDocuments;
	---Purpose : returns Value as a ProductDefinitionWithAssociatedDocuments (Null if another type)

	Representation (me) returns any Representation;
	---Purpose : returns Value as a Representation (Null if another type)

	ExternallyDefinedRepresentation (me) returns any ExternallyDefinedRepresentation;
	---Purpose : returns Value as a Representation (Null if another type)

    	AutoDesignDocumentReference (me) returns AutoDesignDocumentReference;

end AutoDesignGeneralOrgItem;
