-- Created on: 1992-04-13
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Quadric from IntSurf 

	---Purpose: 


uses Ax3         from gp,
     Pnt         from gp,
     Vec         from gp,
     Dir         from gp,
     Lin         from gp,
     Pln         from gp,
     Cylinder    from gp,
     Sphere      from gp,
     Cone        from gp,
     SurfaceType from GeomAbs     

is

    Create
    
        returns Quadric from IntSurf;


    Create(P: Pln from gp)
    
    	returns Quadric from IntSurf;


    Create(C: Cylinder from gp)
    
    	returns Quadric from IntSurf;


    Create(S: Sphere from gp)
    
    	returns Quadric from IntSurf;


    Create(C: Cone from gp)
    
    	returns Quadric from IntSurf;


    SetValue(me: in out; P: Pln from gp)
    
    	is static;


    SetValue(me: in out; C: Cylinder from gp)
    
    	is static;


    SetValue(me: in out; S: Sphere from gp)
    
    	is static;


    SetValue(me: in out; C: Cone from gp)
    
    	is static;


    Distance(me; P: Pnt from gp)
    
    	returns Real from Standard

        is static;


    Gradient(me; P: Pnt from gp)

    	returns Vec from gp
	
	is static;


    ValAndGrad(me; P: Pnt from gp; Dist: out Real from Standard;
               Grad: out Vec from gp)
    
      	is static;


    TypeQuadric(me)
    
    	returns SurfaceType from GeomAbs
	---C++: inline
	
	is static;


    Plane(me)
    
    	returns Pln from gp
	---C++: inline
	
	is static;


    Sphere(me)
    
    	returns Sphere from gp
	---C++: inline
	
	is static;


    Cylinder(me)
    
    	returns Cylinder from gp
	---C++: inline
	
	is static;


    Cone(me)
    
    	returns Cone from gp
	---C++: inline
	
	is static;



    Value(me; U,V: Real)
    
    	returns Pnt from gp
	
	is static;


    D1(me; U,V: Real; P: out Pnt; D1U,D1V: out Vec from gp)
    
	is static;


    DN(me; U,V: Real; Nu,Nv: Integer)
    
    	returns Vec from gp
	
	is static;


    Normale(me; U,V: Real)
    
    	returns Vec from gp
	
	is static;


    Parameters(me; P: Pnt from gp; U,V: out Real)
    
    	is static;


    Normale(me; P: Pnt from gp)
    
    	returns Vec from gp
	
	is static;


fields

    ax3      : Ax3         from gp;
    lin      : Lin         from gp;
    typ      : SurfaceType from GeomAbs;
    prm1     : Real        from Standard;
    prm2     : Real        from Standard;
    prm3     : Real        from Standard;
    prm4     : Real        from Standard;
    ax3direc : Boolean     from Standard;

end Quadric;
