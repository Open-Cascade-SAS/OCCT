-- Created on: 1994-11-25
-- Created by: Frederic MAUPAS
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Builder from TopoDSToStep
    inherits Root from TopoDSToStep

    ---Purpose: This builder Class provides services to build
    --          a ProSTEP Shape model from a Cas.Cad BRep.                 

uses

    FinderProcess                 from Transfer,
    Shape                         from TopoDS,
    Tool                          from TopoDSToStep,
    BuilderError                  from TopoDSToStep,
    TopologicalRepresentationItem from StepShape

raises NotDone from StdFail 
    
is 

--  -----------------------------------------------------------
--  Constructor
--  -----------------------------------------------------------

    Create returns Builder from TopoDSToStep;
    
    Create(S           : Shape from TopoDS;
           T           : in out Tool from TopoDSToStep;
           FP          : FinderProcess from Transfer)
    	returns Builder from TopoDSToStep;
    
    Init(me          : in out;
         S           : Shape from TopoDS;
         T           : in out Tool from TopoDSToStep;
         FP          : FinderProcess from Transfer);
    
--  -----------------------------------------------------------    
--  Get the Result
--  -----------------------------------------------------------

    Error(me) returns BuilderError from TopoDSToStep;
    
    Value (me) returns TopologicalRepresentationItem from StepShape
    	raises NotDone
    	is static;
    	---C++: return const &

fields

    myResult : TopologicalRepresentationItem from StepShape;
    
    myError  : BuilderError                  from TopoDSToStep;

end Builder;
