-- Created on: 1993-08-06
-- Created by: Martine LANGLOIS
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PointPair from StepToTopoDS 

	---Purpose: Stores a pair of Points from step

uses
    CartesianPoint from StepGeom

is
    Create(P1, P2 : CartesianPoint from StepGeom)
    returns PointPair from StepToTopoDS;
    

fields
    myP1 : CartesianPoint from StepGeom;
    myP2 : CartesianPoint from StepGeom;

friends
    class PointPairHasher from StepToTopoDS

end PointPair;
