-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PersonalAddress from StepBasic 

inherits Address from StepBasic 

uses

	HArray1OfPerson from StepBasic, 
	HAsciiString from TCollection, 
	Person from StepBasic
is

	Create returns PersonalAddress;
	---Purpose: Returns a PersonalAddress


	Init (me : mutable;
	      hasAinternalLocation : Boolean from Standard;
	      aInternalLocation : HAsciiString from TCollection;
	      hasAstreetNumber : Boolean from Standard;
	      aStreetNumber : HAsciiString from TCollection;
	      hasAstreet : Boolean from Standard;
	      aStreet : HAsciiString from TCollection;
	      hasApostalBox : Boolean from Standard;
	      aPostalBox : HAsciiString from TCollection;
	      hasAtown : Boolean from Standard;
	      aTown : HAsciiString from TCollection;
	      hasAregion : Boolean from Standard;
	      aRegion : HAsciiString from TCollection;
	      hasApostalCode : Boolean from Standard;
	      aPostalCode : HAsciiString from TCollection;
	      hasAcountry : Boolean from Standard;
	      aCountry : HAsciiString from TCollection;
	      hasAfacsimileNumber : Boolean from Standard;
	      aFacsimileNumber : HAsciiString from TCollection;
	      hasAtelephoneNumber : Boolean from Standard;
	      aTelephoneNumber : HAsciiString from TCollection;
	      hasAelectronicMailAddress : Boolean from Standard;
	      aElectronicMailAddress : HAsciiString from TCollection;
	      hasAtelexNumber : Boolean from Standard;
	      aTelexNumber : HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      hasAinternalLocation : Boolean from Standard;
	      aInternalLocation : HAsciiString from TCollection;
	      hasAstreetNumber : Boolean from Standard;
	      aStreetNumber : HAsciiString from TCollection;
	      hasAstreet : Boolean from Standard;
	      aStreet : HAsciiString from TCollection;
	      hasApostalBox : Boolean from Standard;
	      aPostalBox : HAsciiString from TCollection;
	      hasAtown : Boolean from Standard;
	      aTown : HAsciiString from TCollection;
	      hasAregion : Boolean from Standard;
	      aRegion : HAsciiString from TCollection;
	      hasApostalCode : Boolean from Standard;
	      aPostalCode : HAsciiString from TCollection;
	      hasAcountry : Boolean from Standard;
	      aCountry : HAsciiString from TCollection;
	      hasAfacsimileNumber : Boolean from Standard;
	      aFacsimileNumber : HAsciiString from TCollection;
	      hasAtelephoneNumber : Boolean from Standard;
	      aTelephoneNumber : HAsciiString from TCollection;
	      hasAelectronicMailAddress : Boolean from Standard;
	      aElectronicMailAddress : HAsciiString from TCollection;
	      hasAtelexNumber : Boolean from Standard;
	      aTelexNumber : HAsciiString from TCollection;
	      aPeople : HArray1OfPerson from StepBasic;
	      aDescription : HAsciiString from TCollection) is virtual;

	-- Specific Methods for Field Data Access --

	SetPeople(me : mutable; aPeople : HArray1OfPerson);
	People (me) returns HArray1OfPerson;
	PeopleValue (me; num : Integer) returns Person;
	NbPeople (me) returns Integer;
	SetDescription(me : mutable; aDescription : HAsciiString);
	Description (me) returns HAsciiString;

fields

	people : HArray1OfPerson from StepBasic;
	description : HAsciiString from TCollection;

end PersonalAddress;
