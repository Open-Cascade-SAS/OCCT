-- Created on: 1993-06-08
-- Created by: Laurent BOURESCHE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Iterator from BRepSweep

	---Purpose: This class provides iteration services required by
	--          the Generating Line (TopoDS Shape) of a BRepSweep.
	--          This   tool is  used  to   iterate  on the  direct
	--          sub-shapes of a Shape.
	--          

uses

    Iterator from TopoDS,
    Shape from TopoDS,
    Orientation from TopAbs

raises

    NoMoreObject from Standard,
    NoSuchObject from Standard

is

    Create;

    Init(me : in out; aShape: Shape from TopoDS)
	---Purpose: Resest the Iterator on sub-shapes of <aShape>.
    is static;
    
    More(me) returns Boolean
	---Purpose: Returns True if there is a current sub-shape.
	--          
	---C++: inline
    is static;
    
    Next(me : in out)
	---Purpose: Moves to the next sub-shape.
    raises
    	NoMoreObject from Standard
    is static;
    
    Value(me) returns Shape from TopoDS
	---Purpose: Returns the current sub-shape.
    raises
    	NoSuchObject from Standard
	---C++: return const &
	---C++: inline
    is static;
    
    Orientation(me) returns Orientation from TopAbs
	---Purpose: Returns the orientation of the current sub-shape.
    raises
    	NoSuchObject from Standard
	---C++: inline
    is static;

fields

    myIterator : Iterator from TopoDS;

end Iterator from BRepSweep;
