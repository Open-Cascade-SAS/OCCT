-- Created on: 1997-08-26
-- Created by: SMO
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package MPrsStd 

	---Purpose: Storage    and  Retrieval  drivers   for graphic
	--          attributes.   Transient  attributes are defined in
	--          package TPrsStd and persistent one are defined in
	--          package PPrsStd

uses TDF,
     PDF,
     MDF, 
     CDM

is

    	    ---Category: StorageDriver

	class AISPresentationStorageDriver;
	class PositionStorageDriver;


        ---Category: RetrievalDriver

        class AISPresentationRetrievalDriver;
        class AISPresentationRetrievalDriver_1;	
	class PositionRetrievalDriver;
	
    AddStorageDrivers(aDriverTable : ASDriverHSequence from MDF;theMessageDriver : MessageDriver from CDM);
	---Purpose: Adds the attribute storage drivers to <aDriverTable>.
    	---Category: StorageDriversTable


    AddRetrievalDrivers(aDriverTable : ARDriverHSequence from MDF;theMessageDriver : MessageDriver from CDM);
	---Purpose: Adds the attribute retrieval drivers to <aDriverTable>.
    	---Category: RetrievalDriversTable


end MPrsStd;



