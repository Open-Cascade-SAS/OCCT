-- File:        MechanicalDesignGeometricPresentationRepresentation.cdl
-- Created:     Mon Dec  4 12:02:28 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWMechanicalDesignGeometricPresentationRepresentation from RWStepVisual

	---Purpose : Read & Write Module for MechanicalDesignGeometricPresentationRepresentation

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     MechanicalDesignGeometricPresentationRepresentation from StepVisual,
     EntityIterator from Interface

is

	Create returns RWMechanicalDesignGeometricPresentationRepresentation;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable MechanicalDesignGeometricPresentationRepresentation from StepVisual);

	WriteStep (me; SW : in out StepWriter; ent : MechanicalDesignGeometricPresentationRepresentation from StepVisual);

	Share(me; ent : MechanicalDesignGeometricPresentationRepresentation from StepVisual; iter : in out EntityIterator);

end RWMechanicalDesignGeometricPresentationRepresentation;
