-- Created on: 1997-03-03
-- Created by: Jean-Pierre COMBE
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SymmetricRelation from AIS inherits Relation from AIS

	---Purpose: A framework to display constraints of symmetricity
    	-- between two or more datum Interactive Objects.
    	-- A plane serves as the axis of symmetry between the
    	-- shapes of which the datums are parts.

uses Shape                 from TopoDS,
     Presentation          from Prs3d,
     PresentationManager3d from PrsMgr,
     Selection             from SelectMgr,
     Dir                   from gp,
     Pnt                   from gp,
     Projector             from Prs3d,
     Transformation        from Geom,
     ExtendedString        from TCollection,
     Plane                 from Geom

is
    Create(aSymmTool   : Shape from TopoDS;
    	   FirstShape  : Shape from TopoDS;
    	   SecondShape : Shape from TopoDS;
	   aPlane      : Plane from Geom)
    returns SymmetricRelation from AIS;
    	--- Purpose: Constructs an object to display constraints of symmetricity.
    	-- This object is defined by a tool aSymmTool, a first
    	-- shape FirstShape, a second shape SecondShape, and a plane aPlane.
    	-- aPlane serves as the axis of symmetry.
    	-- aSymmTool is the shape composed of FirstShape
    	-- SecondShape and aPlane. It may be queried and
    	-- edited using the functions GetTool and SetTool.
    	-- The two shapes are typically two edges, two vertices or two points.   

    IsMovable(me) returns Boolean from Standard 
    	---Purpose: Returns true if the symmetric constraint display is movable.
    	---C++: inline       
      
    is redefined;        
    
    SetTool(me:mutable; aSymmetricTool : Shape from TopoDS);
        ---Purpose: Sets the tool aSymmetricTool composed of a first
    	-- shape, a second shape, and a plane.
    	-- This tool is initially created at construction time.
        ---C++: inline

    GetTool(me)
    	---Purpose: Returns the tool composed of a first shape, a second
    	-- shape, and a plane. This tool is created at construction time.
 	---C++: inline
   	---C++: return const &
    returns Shape from TopoDS;
    
-- Methods from PresentableObject

    Compute(me            : mutable;
  	    aPresentationManager: PresentationManager3d from PrsMgr;
    	    aPresentation : Presentation from Prs3d;
    	    aMode         : Integer from Standard= 0) 
    is redefined static private;
    
    Compute(me:mutable;
    	        aProjector: Projector from Prs3d;
                aPresentation: Presentation from Prs3d)
    is redefined static private;     

    Compute(me            : mutable;
    	    aProjector    : Projector from Prs3d;
    	    aTrsf         : Transformation from Geom;
	    aPresentation : Presentation from Prs3d)
    is redefined;
    	---Purpose: computes the presentation according to a point of view
    	--          given by <aProjector>. 
    	--          To be Used when the associated degenerated Presentations 
    	--          have been transformed by <aTrsf> which is not a Pure
    	--          Translation. The HLR Prs can't be deducted automatically
    	--          WARNING :<aTrsf> must be applied
    	--           to the object to display before computation  !!!

--     SymmetricRelation Methods from SelectableObject

    ComputeSelection(me         : mutable;
    	    	     aSelection : Selection from SelectMgr;
    	    	     aMode      : Integer from Standard)is private;

--
--     Computation private methods
--

    ComputeTwoFacesSymmetric(me: mutable; aprs : Presentation from Prs3d)
    is private;
    
    ComputeTwoEdgesSymmetric(me: mutable; aprs : Presentation from Prs3d)
    is private;
    
    ComputeTwoVerticesSymmetric(me: mutable; aprs : Presentation from Prs3d)
    is private;
    
    
fields

    myTool          : Shape from TopoDS;
    myFAttach       : Pnt   from gp;
    mySAttach       : Pnt   from gp;
    myFDirAttach    : Dir   from gp;
    myAxisDirAttach : Dir   from gp;
    
end SymmetricRelation;
