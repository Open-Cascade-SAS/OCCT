-- Created on: 1999-02-15
-- Created by: Andrey BETENEV
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class SurfaceCurveAndBoundedCurve from StepGeom 
    inherits SurfaceCurve from StepGeom

	---Purpose: complex type: bounded_curve + surface_curve
	--          needed for curve_bounded_surfaces (S4132)

uses
    
    BoundedCurve from StepGeom

is

    Create returns mutable SurfaceCurveAndBoundedCurve;
	---Purpose: creates empty object

    BoundedCurve (me: mutable) returns mutable BoundedCurve from StepGeom;
        ---Purpose: returns field BoundedCurve
	---C++: return &

fields

    myBoundedCurve : BoundedCurve from StepGeom;

end SurfaceCurveAndBoundedCurve;
