-- Created on: 2003-06-02
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 2003-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package StepDimTol


    ---Purpose :Collects definition of STEP GD&T entities TR12J
    	

uses    TCollection,
     	StepRepr, 
    	StepShape,
    	StepVisual,
	StepBasic,
    	TColStd, 
    	StepData, 
    	Interface, 
    	MMgt

is 

enumeration LimitCondition is 
   MaximumMaterialCondition,
   LeastMaterialCondition,
   RegardlessOfFeatureSize
end;
    
    class ShapeToleranceSelect;
    class AngularityTolerance;
    class CircularRunoutTolerance;
    class ConcentricityTolerance;
    class CylindricityTolerance;
    class CoaxialityTolerance;
    class FlatnessTolerance;
    class LineProfileTolerance;
    class ParallelismTolerance;
    class PerpendicularityTolerance;
    class PositionTolerance;
    class RoundnessTolerance;
    class StraightnessTolerance;
    class SurfaceProfileTolerance;
    class SymmetryTolerance;
    class TotalRunoutTolerance;
    
    class GeometricTolerance;
    class GeometricToleranceRelationship;
    class GeometricToleranceWithDatumReference;
    class ModifiedGeometricTolerance;
     
    class Datum;
    class DatumFeature;
    class DatumReference;
    class CommonDatum;
    class DatumTarget;
    class PlacedDatumTargetFeature;

    class GeoTolAndGeoTolWthDatRefAndModGeoTolAndPosTol;

    imported Array1OfDatumReference;
    imported transient class HArray1OfDatumReference;
    
end StepDimTol;
