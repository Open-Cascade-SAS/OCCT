-- File:        PlotMgt_PlotterParameter.cdl
-- Created:     Quebex 30 October 1998
-- Author:      DCB
---Copyright:   MatraDatavision 1998

class PlotterParameter from PlotMgt inherits TShared from MMgt

uses
  FStream                 from Aspect,
  Plotter                 from PlotMgt,
  TypeOfPlotterParameter  from PlotMgt,
  HSequenceOfAsciiString  from TColStd,
  AsciiString             from TCollection,
  File                    from OSD

is
  -------------------------
  -- Category: Constructors
  -------------------------
  Create (
    aName  : AsciiString from TCollection
  ) returns mutable PlotterParameter from PlotMgt;
  ---Purpose: Create the class instance WITH undefined TYPE

  -----------------------------------------------
  -- Category: Methods to change class definition
  -----------------------------------------------
  Save (me: mutable; aFile: in out File from OSD)
  returns Boolean from Standard;
  ---Purpose:

  SetState (me: mutable; aState: Boolean from Standard);
  ---Purpose:

  SetType (me: mutable; aType: TypeOfPlotterParameter from PlotMgt);
  ---Purpose:

  ProcessParamVal (me: mutable;
    aParamSign :     CString from Standard;
    aFlag      :     Integer from Standard;
    aValue     : out AsciiString from TCollection
  ) is private;

  CheckListValue (me: mutable
  ) returns Boolean from Standard is private;
  ---Purpose:

  Normalize (me: mutable)
  is protected;
  ---Purpose:

  ----------------------------
  -- Category: Inquire methods
  ----------------------------
  SValue (me; aValue: out AsciiString from TCollection);
  ---Purpose:

  BValue (me)
  returns Boolean from Standard;
  ---Purpose:

  IValue (me)
  returns Integer from Standard;
  ---Purpose:

  RValue (me)
  returns Real from Standard;
  ---Purpose:

  LValues (me; aList: out HSequenceOfAsciiString from TColStd);
  ---Purpose:

  MValue (me
  ) returns HSequenceOfAsciiString from TColStd;
  ---Purpose:

  Name (me)
  returns AsciiString from TCollection;
  ---Purpose:

  OldName (me)
  returns AsciiString from TCollection;
  ---Purpose:

  Description (me : mutable)
  returns HSequenceOfAsciiString from TColStd
  is protected;
  ---Purpose:
  ---C++: return &

  NeedToBeSaved (me)
  returns Boolean from Standard;
  ---Purpose:

  Dump (me);
  ---Purpose:

  PutCommandInfo (me; outStream: FStream from Aspect);
  ---Purpose: Used to put parameter's information in a cmd file
  -- used in PlotterDriver's Spool method.

  ----------------------------------------
  -- Category: Methods to modify parameter
  ----------------------------------------
  SetSValue (me: mutable; aValue: AsciiString from TCollection);
  ---Purpose:

  SetBValue (me: mutable; aValue: Boolean from Standard);
  ---Purpose:

  SetIValue (me: mutable; aValue: Integer from Standard);
  ---Purpose:

  SetRValue (me: mutable; aValue: Real from Standard);
  ---Purpose:

  SetMValue (me: mutable; aMap: HSequenceOfAsciiString from TColStd);
  ---Purpose:

fields
  myName           : AsciiString            from TCollection;
  myOldName        : AsciiString            from TCollection;
  myType           : TypeOfPlotterParameter from PlotMgt;
  myIndex          : Integer                from Standard;
  myState          : Boolean                from Standard;
  myConfigState    : Boolean                from Standard;
  myIsModified     : Boolean                from Standard;
  --------------------------------------------------------
  myFlags          : Integer                from Standard;
  myDialog         : AsciiString            from TCollection;
  myMinValue       : AsciiString            from TCollection;
  myMaxValue       : AsciiString            from TCollection;
  myValues         : AsciiString            from TCollection;
  myDefValue       : AsciiString            from TCollection;
  myMapLength      : Integer                from Standard;
  myMap            : HSequenceOfAsciiString from TColStd;

  myDescription    : HSequenceOfAsciiString from TColStd;

friends
  class Plotter from PlotMgt

end PlotterParameter from PlotMgt;
