-- Created on: 1992-06-04
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package Geom2dInt 

	---Purpose: Intersection between two Curves2 from Geom2dAdaptor

        ---Level: Public
        --
        -- All the methods of the classes are public.
        --


uses Standard, gp, TColStd, GeomAbs, Geom2d, Adaptor3d, Adaptor2d, IntCurve

is

   class Geom2dCurveTool;
    	 
   class GInter instantiates IntCurveCurveGen from IntCurve
            (Curve2d         from Adaptor2d,
             Geom2dCurveTool from Geom2dInt);

end Geom2dInt; 
 
