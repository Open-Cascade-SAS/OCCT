-- Created on: 2004-05-13
-- Created by: Sergey ZARITCHNY <szy@opencascade.com>
-- Copyright (c) 2004-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class NamingDriver from BinMNaming inherits ADriver from BinMDF

	---Purpose: Naming  Attribute Driver.

uses
    SRelocationTable from BinObjMgt,
    RRelocationTable from BinObjMgt,
    Persistent       from BinObjMgt,
    MessageDriver    from CDM,
    Attribute        from TDF


is
    Create (theMessageDriver:MessageDriver from CDM)
        returns NamingDriver from BinMNaming;

    NewEmpty (me)  returns Attribute from TDF;

    Paste(me; Source     : Persistent from BinObjMgt;
              Target     : Attribute from TDF;
              RelocTable : out RRelocationTable from BinObjMgt)
        returns Boolean from Standard;

    Paste(me; Source     : Attribute from TDF;
              Target     : in out Persistent from BinObjMgt;
              RelocTable : out SRelocationTable from BinObjMgt);
    

end NamedShapeDriver;

