-- Created on: 1993-01-11
-- Created by: CKY / Contract Toubro-Larsen ( Anand NATRAJAN )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class NodalConstraint from IGESAppli  inherits IGESEntity

        ---Purpose: defines NodalConstraint, Type <418> Form <0>
        --          in package IGESAppli
        --          Relates loads and/or constraints to specific nodes in
        --          the Finite Element Model by creating a relation between
        --          Node entities and Tabular Data Property that contains
        --          the load or constraint data

uses

        TabularData          from IGESDefs,
        Node                 from IGESAppli,
        HArray1OfTabularData from IGESDefs

raises OutOfRange

is

        Create returns NodalConstraint;

        -- Specific Methods pertaining to the class

        Init (me         : mutable;
              aType      : Integer;
              aNode      : Node;
              allTabData : HArray1OfTabularData);
        ---Purpose : This method is used to set the fields of the class
        --           NodalConstraint
        --       - aType      : Loads / Constraints
        --       - aNode      : the Node
        --       - allTabData : Tabular Data Property carrying the load
        --                      or constraint vector

        NbCases (me) returns Integer;
        ---Purpose : returns total number of cases

        Type (me) returns Integer;
        ---Purpose : returns whether Loads (1) or Constraints (2)

        NodeEntity (me) returns Node;
        ---Purpose : returns the Node

        TabularData (me; Index : Integer) returns TabularData
        raises OutOfRange;
        ---Purpose : returns Tabular Data Property carrying load or constraint vector
        -- raises exception if Index <= 0 or Index > NbCases

fields

--
-- Class    : IGESAppli_NodalConstraint
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class NodalConstraint.
--
-- Reminder : A NodalConstraint instance is defined by :
--            - indicator whether Loads or Constraints
--            - a Node
--            - Tabular Data Property carrying load or constraint vector

        theType             : Integer;
        theNode             : Node;
        theTabularDataProps : HArray1OfTabularData;

end NodalConstraint;
