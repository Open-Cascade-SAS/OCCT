-- Created on: 1993-01-27
-- Created by: Isabelle GRIGNON
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PolyArc from IntPatch

inherits Polygo from IntPatch

uses Box2d         from Bnd,
     Pnt2d         from gp,
     Array1OfPnt2d from TColgp,
     Array1OfReal  from TColStd,
     HCurve2d from Adaptor2d

raises ConstructionError from Standard

is

    Create(A: HCurve2d from Adaptor2d; NbSample: Integer from Standard; 
    	   Pfirst,Plast : Real from Standard;
           BoxOtherPolygon: Box2d from Bnd)

    	---Purpose: Creates the polygon of the arc A on the surface S.
    	--          The arc is limited by the parameters Pfirst and Plast.
    	--          None of these parameters can be infinite.

    	returns PolyArc from IntPatch
	
	raises ConstructionError from Standard;
    	--- This exception is raised if Pfirst=RealFirst or Plast=RealLast or
    	--  NbSample<=1.

    Closed(me)                   returns Boolean from Standard is redefined virtual;

    NbPoints(me)                 returns Integer;
 
    Point(me; Index : Integer)   returns Pnt2d from gp;
                                      	    	 
    Parameter(me ; Index : Integer) returns Real from Standard;
     
    SetOffset(me:in out;  OffsetX,OffsetY: Real from Standard);
       
		
fields

    brise  : Array1OfPnt2d from TColgp;
    param  : Array1OfReal  from TColStd;
    offsetx: Real          from Standard;
    offsety: Real          from Standard;
    ferme  : Boolean       from Standard;

end PolyArc;
