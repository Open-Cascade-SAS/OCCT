-- Created on: 1995-02-27
-- Created by: Christian CAILLET
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class BinderOfTransientInteger  from Transfer  inherits SimpleBinderOfTransient

    ---Purpose : This type of Binder allows to attach as result, besides a
    --           Transient Object, an Integer Value, which can be an Index
    --           in the Object if it defines a List, for instance
    --           
    --           This Binder is otherwise a kind of SimpleBinderOfTransient,
    --           i.e. its basic result (for iterators, etc) is the Transient

uses Integer

is

    Create returns mutable BinderOfTransientInteger;
    ---Purpose : Creates an empty BinderOfTransientInteger; Default value for
    --           the integer part is zero

    SetInteger (me : mutable; value : Integer);
    ---Purpose : Sets a value for the integer part

    Integer (me) returns Integer;
    ---Purpose : Returns the value set for the integer part

fields

    theintval : Integer;

end BinderOfTransientInteger;
