-- Created on: 1998-06-30
-- Created by: Christian CAILLET
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class DocumentReference  from StepBasic    inherits TShared from MMgt

uses
     Document from StepBasic,
     HAsciiString from TCollection

is

    Init0 (me : mutable;
    	   aAssignedDocument : Document;
	   aSource : HAsciiString);

    AssignedDocument (me) returns Document;
    SetAssignedDocument (me : mutable; aAssignedDocument : Document);

    Source (me) returns HAsciiString;
    SetSource (me : mutable; aSource : HAsciiString);

fields

    theAssignedDocument : Document;
    theSource : HAsciiString;

end DocumentReference;
