
-- File:	Graphic2d_Primitive.cdl
-- Created:	Tue Jun 22 16:33:45 1993
-- Author:	Jean Louis FRENKEL, Gerard GRAS.
--		<jlf@stylox>
-- Updated:	GG 19/08/98 PERFORMANCE 
--		A new method ComputeMinMax(...) could be redefined for 
--		each primitive to recompute the MinMax values at the right time.
--		GG 14/04/00 G002 Add SetPickedIndex() method
--				 Add DrawElement() and DrawVertex() methods
--		GG 05/05/00 G002 Add IsOn() method.
--				 Add Highlight(),Unhilight(),IsHighlighted()
--				 HighlightIndex() methods.
--	TCL : 12-06-00 : G002 : new method Pick( Xmin, Ymin, Xmax, Ymax,...)
--	TCL : 07-07-00 : G002 : new method HighlightIndices()
--				method HighlightIndex() was removed
--	TCL : 25-07-00 : G002 : new methods SetDisplayMode( aMode ) and DisplayMode()

--      SAV : 14/11/01 : Added a set of methods (marked SAV before declaration)
--                       to provide highlighting/selection
--                       of SetOfMarkers elements. These methods should be redefined
--                       for other SetOf<>.
--                       
--      SAV : 03/07/02 : SetElementsSelected() prototype changed to avoid regression
--                       during elements single selection.
---Copyright:	 Matra Datavision 1993

deferred class Primitive from Graphic2d inherits TShared from MMgt

	---Version:

	---Purpose: Groups all drawing elements which can be stored
	--	    in a graphic object.
	--	    Each primitive have a postion in the space model.

uses

	Buffer		   from Graphic2d,
	GOPtr		   from Graphic2d,
	Drawer		   from Graphic2d,
	GraphicObject	   from Graphic2d,
	TypeOfPrimitive	   from Graphic2d,
	Length		   from Quantity,
	PickMode	   from Graphic2d,
	HSequenceOfInteger from TColStd,
--	IFStream	   from Aspect,
	FStream		   from Aspect,
	MapOfInteger       from TColStd

is
	-------------------------
	-- Category: Constructors
	-------------------------

	Initialize (aGraphicObject: GraphicObject from Graphic2d);
	---Level: Public
	---Purpose: Creates a primitive in a graphic object <aGraphicObject>.
	---Category: Constructors

	----------------------------------------------
	-- Category: Methods to manage color attribute
	----------------------------------------------

	SetColorIndex(me: mutable; anIndex: Integer from Standard)
		is static;
	---Level: Public
	---Purpose: Defines the index, in the color map, of the primitive color.
	--  Warning: For an image, this method defines the color of the
	--	    boundary rectangle.
	---Category: Methods to manage color attribute

	ColorIndex (me)
		returns Integer from Standard
		is static;
	---Level: Public
	---Purpose: Returns the index, in the color map, of the primitive color.
	--  Warning: For an image, it is the color of the border.
	---Category: Methods to manage color attribute

	--------------------------
	-- Category: Draw and Pick
	--------------------------

	Draw (me : mutable; aDrawer: Drawer from Graphic2d)
	is deferred;
	---Level: Internal
	---Purpose: Draws the primitive <me>.

	DrawElement (me : mutable; aDrawer: Drawer from Graphic2d;
				   anElement: Integer from Standard)
	is virtual protected;
	---Level: Internal
	---Purpose: Draws the element <anElement> of the primitive <me>.

    	---SAV
	DrawPickedElements(me : mutable; aDrawer: Drawer from Graphic2d )
	is virtual protected;
	---Level: Internal
	---Purpose: Draws the all picked elements of the primitive <me>.

    	---SAV
    	DrawSelectedElements(me : mutable; aDrawer: Drawer from Graphic2d )
	is virtual protected;
	---Level: Internal
	---Purpose: Draws the all picked elements of the primitive <me>.

    	---SAV
    	SetElementsSelected(me : mutable) returns Boolean from Standard
	is virtual;
	---Level: Public
	---Purpose: Declares that previously highlighted elements will be selected ones.
	--  Warning: If a descendant redefines this method then it  must return <true>!

    	---SAV
    	HasSelectedElements(me : mutable)
	returns Boolean from Standard is virtual;
	---Level: Public

    	---SAV
    	ClearSelectedElements(me : mutable)
	is virtual;
	---Level: Public

	DrawVertex (me : mutable; aDrawer: Drawer from Graphic2d;
				  aVertex: Integer from Standard)
	is virtual protected;
	---Level: Internal
	---Purpose: Draws the vertex <aVertex> of the primitive <me>.

	Pick (me : mutable; X, Y: ShortReal from Standard;
		aPrecision: ShortReal from Standard;
		aDrawer: Drawer from Graphic2d)
	returns Boolean from Standard
	is deferred protected;
	---Level: Internal
	---Purpose: Returns Standard_True if the primitive <me> is picked,
	--	    Standard_False if not.

    	---SAV
	PickByCircle (me : mutable; X, Y, Radius : ShortReal from Standard;
		    	    aDrawer: Drawer from Graphic2d;
		    	    aPickMode: PickMode from Graphic2d = Graphic2d_PM_INCLUDE )
	returns Boolean from Standard
	is virtual protected;
	---Level: Internal
	---Purpose: Returns Standard_True if the primitive <me> is picked,
	--	    Standard_False if not.

	Pick( me: mutable; Xmin, Ymin, Xmax, Ymax: ShortReal from Standard;
		  aDrawer: Drawer from Graphic2d; 
		  aPickMode: PickMode from Graphic2d = Graphic2d_PM_INCLUDE )
	returns Boolean from Standard is virtual protected;
	---Level: Internal
	---Purpose: Returns Standard_True if the primitive <me> is:
	--		included in rectangle (<aPickMode = PM_INCLUDE>),
	--		excluded from rectangle (<aPickMode = PM_EXLUDE>),
	--		intersected by rectangle (<aPickMode = PM_INTERSECT>),
	--		defined by Xmin, Ymin, Xmax, Ymax. 
	--	    Standard_False if not.

	NumOfElemIndices( me ) returns Integer from Standard
		is virtual;
	---Level: Internal
	---Purpose: Returns number of elements of primitive

	NumOfVertIndices( me ) returns Integer from Standard
		is virtual;
	---Level: Internal
	---Purpose: Returns number of vertices of primitive

	SetPickedIndex (me : mutable; anIndex: Integer from Standard)
	is static protected;
	---Level: Public
	---Purpose: Sets the index of the picked primitive element if any.
	---Category: Methods to manage picking 

	PickedIndex (me) returns Integer from Standard is static;
	---Level: Public
	---Purpose: Returns the index of the last picked primitive element.
	--  Warning: This is available only if the Pick() method has
	--         returned Standard_True.
	---Category: Methods to manage picking 

    
    	---SAV
    	PickedIndices(me) returns MapOfInteger from TColStd is static;
	---C++: return const &

	Highlight (me: mutable;
		   anIndex: Integer from Standard = 0)
	is static;
	---Level: Public
	---Purpose: Highlights the primitive <me> or a part of the
	--	    primitive with the override color of the view.
	--	    When <anIndex> is 0 all the primitive is highlighted
	--		 >0 only the requested element is highlighted.
	--		 <0 only the requested vertex is highlighted.
	---Category: Methods to manage the highlight

	Unhighlight (me: mutable)
	is static;
	---Level: Public
	---Purpose: Suppress the highlight on the primitive <me>.
	---Category: Methods to manage the highlight

	IsHighlighted (me)
	returns Boolean from Standard
	is static;
	---Level: Public
	---Purpose: Returns Standard_True if the primitive <me>
	--          is highlighted, Standard_False if not.
	---Category: Methods to manage the highlight

	HighlightIndices(me) returns HSequenceOfInteger from TColStd;
	---Level: Public
	---Purpose: Returns the sequence of highlight indices of the primitive <me>
	---Category: Methods to manage the highlight

	SetDisplayMode( me: mutable; aMode: Integer from Standard );
	---Level    : Public;
	---Purpose  : Sets the display mode of primitive
	---Category : Methods to manage the display mode

	DisplayMode( me ) returns Integer from Standard;
	---Level    : Public;
	---Purpose  : Indicates the display mode of primitive
	---Category : Methods to manage the display mode


	----------------------------
	-- Category: Private methods
	----------------------------

	MinMax (me : mutable; Minx, Maxx, Miny, Maxy: out ShortReal from Standard)
		returns Boolean from Standard is static;
	---Level: Internal
	---Purpose: Returns TRUE and the min max values of <me>.
	--	    or FALSE when the primitive is empty.
	--	    Called by the method Graphic2d_GraphicObject::MinMax

	ComputeMinMax (me : mutable)
	returns Boolean from Standard is virtual protected;
	---Level: Internal
	---Purpose: Computes the MinMax of the primitive if possible.

	IsOn( myclass;
	  aX1, aY1, aX2, aY2,
	  aPrecision: ShortReal from Standard)
	returns Boolean from Standard is protected ;
	---Level: Internal
	---Purpose: Returns Standard_True if (<aX1>, <aY1>) is closed
	--          to the point (<aX2>, <aY2>).
	---Category: Class methods

	IsInMinMax (me : mutable; X, Y: ShortReal from Standard;
		aPrecision: ShortReal from Standard)
	returns Boolean from Standard;
	---Level: Internal
	---Purpose: Returns Standard_True if the point <X>, <Y> is in the
	--	    rectangle defined by the min max values of <me>.
	--  Warning: If <me> is in a transformed GraphicObject then
	--	    the min max values are transformed.

	Drawer(me) returns mutable Drawer from Graphic2d is protected;
	---Level: Internal
	---Purpose: Returns the attached drawer of the view of this Primitive.
	---Category: Inquiries

	PGraphicObject(me) returns GOPtr from Graphic2d is private;
	---Level: Internal
	---Purpose: Returns the graphic-object back pointer of this Primitive.
	---Category: Inquiries

	ResetIndex (me: mutable) is protected;
	---Level: Internal
	---Purpose: Resets the starting traversal index to this primitive.

	SetFamily (me : mutable; aFamily: TypeOfPrimitive from Graphic2d)
		is protected;
	---Level: Internal
	---Purpose: Sets the family of this primitive.

	Family (me) returns TypeOfPrimitive is protected;
	---Level: Internal
	---Purpose: Returns the family of this primitive

	----------------------------------------------------------------------

	Save(me; aFStream: in out FStream from Aspect) is deferred;
--	Retrieve(me; anIFStream: in out IFStream from Aspect) is deferred;

fields

	myGOPtr           : GOPtr              from Graphic2d is protected;
	myMinX            : ShortReal          from Standard  is protected;
	myMinY            : ShortReal          from Standard  is protected;
	myMaxX            : ShortReal          from Standard  is protected;
	myMaxY            : ShortReal          from Standard  is protected;
	myColorIndex      : Integer            from Standard  is protected;
	myPickedIndex     : Integer            from Standard;
	---SAV
	myPickedIndices   : MapOfInteger       from TColStd   is protected;
	myTypeOfPrimitive : TypeOfPrimitive    from Graphic2d;
	mySeqOfHighInd    : HSequenceOfInteger from TColStd;
	myNumOfElem       : Integer            from Standard  is protected;
	myNumOfVert       : Integer            from Standard  is protected;
	myDisplayMode     : Integer            from Standard  is protected;

friends

	class Buffer from Graphic2d,

	Draw from class GraphicObject from Graphic2d
		(me: mutable;
		 aDrawer: Drawer from Graphic2d;
		 Reset: Boolean from Standard),

	Draw from class GraphicObject from Graphic2d
		(me: mutable;
		 aDrawer: Drawer from Graphic2d;
		 aPrimitive: Primitive from Graphic2d),

	Pick from class GraphicObject from Graphic2d
		(me : mutable;
		 X, Y: Real from Standard;
		 aPrecision: Real from Standard;
		 aDrawer: Drawer from Graphic2d),

    	---SAV
	PickByCircle from class GraphicObject from Graphic2d
		(me : mutable;
		 X, Y: Real from Standard;
		 Radius: Real from Standard;
		 aDrawer: Drawer from Graphic2d),


	Pick from class GraphicObject from Graphic2d
		( me : mutable;
		 Xmin, Ymin, Xmax, Ymax: Real from Standard;
		 aDrawer: Drawer from Graphic2d;
		 aPickMode: PickMode from Graphic2d ),

	MinMax from class GraphicObject from Graphic2d
		(me;
		 Minx, Maxx, Miny, Maxy: out Length from Quantity),

	MarkerMinMax from class GraphicObject from Graphic2d
		(me;
		 Minx, Maxx, Miny, Maxy: out Length from Quantity),

	RemovePrimitive from class GraphicObject from Graphic2d
		(me: mutable;
		 aPrimitive: Primitive from Graphic2d),

	Draw from class TransientManager from Graphic2d
		(me: mutable;
		aPrimitive: Primitive from Graphic2d), 

	DrawElement from class TransientManager from Graphic2d
		(me: mutable;
		aPrimitive: Primitive from Graphic2d; 
		anIndex: Integer from Standard),

	DrawVertex from class TransientManager from Graphic2d
		(me: mutable;
		aPrimitive: Primitive from Graphic2d; 
		anIndex: Integer from Standard),

    	---SAV
	DrawPickedElements from class TransientManager from Graphic2d
    	    	(me : mutable;
    	    	 aPrimitive   : Primitive from Graphic2d )

end Primitive from Graphic2d;
