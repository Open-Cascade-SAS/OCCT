-- Created on: 1994-02-14
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



generic class ZerCOnSSParFunc from IntImp 
    (ThePSurface     as any;
     ThePSurfaceTool as any;   --as PSurfaceTool from IntImp(ThePSurface)
     TheCurveOnSurf  as any;
     TheCurveTool    as any     --as COnSCurveTool from IntImp(TheCurve)
    )
    
inherits FunctionSetWithDerivatives from math

      	---Purpose: this function is associated to the intersection between 
      	--          a curve on surface and a surface  .


uses Vector from math,
     Matrix from math,
     Pnt from gp

is
    Create( S1 : ThePSurface;
    	    C  : TheCurveOnSurf;
            S2 : ThePSurface )

	---Purpose: S1 is the surface on which the intersection is searched.
	--          C is a curve on the surface S2.

    	returns ZerCOnSSParFunc from IntImp;
	    

    NbVariables(me) returns Integer from Standard
    is static;
    
    NbEquations(me) returns Integer from Standard
    is static;
    
    Value(me : in out; X : in Vector from math;
    	    	       F : out Vector from math)
    returns Boolean from Standard
    is static;
    
    Derivatives(me : in out;X : in  Vector from math;
    	    	    	    D : out Matrix from math)
    returns Boolean from Standard
    is static;
    
    Values(me : in out;
    	   X  : in Vector from math;
	   F  : out Vector from math; D: out Matrix from math)
    returns Boolean from Standard
    is static;

    Point(me)
    	---C++: return const&
    	returns Pnt from gp
    	is static;
    
    Root(me) returns Real from Standard
    is static;
    
    AuxillarSurface(me)
    	---C++: return const&
    	returns ThePSurface
    	is static;

    AuxillarCurve(me)
    	---C++: return const&
    	returns TheCurveOnSurf
    	is static;
    
fields
     curve    : Address from Standard; --- TheCurveOnSurf;
     surface1 : Address from Standard; --- ThePSurface;
     surface2 : Address from Standard; --- ThePSurface;
     p	      : Pnt from gp;
     f        : Real from Standard;
     
end ZerCOnSSParFunc;
