-- Created on: 2004-05-17
-- Created by: Sergey ZARITCHNY <szy@opencascade.com>
-- Copyright (c) 2004-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package BinMPrsStd 

	---Purpose: 

uses 
    BinObjMgt, 
    TDF, 
    BinMDF,
    CDM
is
        ---Category: Storage-Retrieval drivers for graphic attributes from
        --           TPrsStd

	class AISPresentationDriver; 
	
	class PositionDriver;	
	
    AddDrivers(theDriverTable   : ADriverTable  from BinMDF;
    	       theMessageDriver : MessageDriver from CDM);
	---Purpose: Adds the attribute storage-retrieval driver to <theDriverTable>.

end BinMPrsStd;
