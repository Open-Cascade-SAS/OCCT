-- Created on: 2000-04-18
-- Created by: Andrey BETENEV
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0

class DimensionalCharacteristicRepresentation from StepShape
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity DimensionalCharacteristicRepresentation

uses
    DimensionalCharacteristic from StepShape,
    ShapeDimensionRepresentation from StepShape

is
    Create returns DimensionalCharacteristicRepresentation from StepShape;
	---Purpose: Empty constructor

    Init (me: mutable; aDimension: DimensionalCharacteristic from StepShape;
                       aRepresentation: ShapeDimensionRepresentation from StepShape);
	---Purpose: Initialize all fields (own and inherited)

    Dimension (me) returns DimensionalCharacteristic from StepShape;
	---Purpose: Returns field Dimension
    SetDimension (me: mutable; Dimension: DimensionalCharacteristic from StepShape);
	---Purpose: Set field Dimension

    Representation (me) returns ShapeDimensionRepresentation from StepShape;
	---Purpose: Returns field Representation
    SetRepresentation (me: mutable; Representation: ShapeDimensionRepresentation from StepShape);
	---Purpose: Set field Representation

fields
    theDimension: DimensionalCharacteristic from StepShape;
    theRepresentation: ShapeDimensionRepresentation from StepShape;

end DimensionalCharacteristicRepresentation;
