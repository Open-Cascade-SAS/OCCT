-- Created on: 1993-06-22
-- Created by: Jean Louis FRENKEL, Gerard GRAS
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


-- Modified: TCL G002, 07-08-00, new inquire methods FirstPoint, SecondPoint


class Segment from Graphic2d inherits Line from Graphic2d

	---Version:

	---Purpose: The primitive Segment

	---Keywords: Primitive, Segment
	---Warning:
	---References:

uses
	Drawer		from Graphic2d,
	GraphicObject	from Graphic2d,
	Length		from Quantity,
	FStream		from Aspect,
	IFStream	from Aspect

raises
	SegmentDefinitionError	from Graphic2d

is
	-------------------------------------
	-- Category: Constructors
	-------------------------------------

	Create (aGraphicObject: GraphicObject from Graphic2d;
		X1, Y1, X2, Y2: Length from Quantity)
	returns mutable Segment from Graphic2d
	---Level: Public
	---Purpose: Creates a segment in the graphic object <aGraphicObject>.
	--	    The first point is <X1>, <Y1>.
	--	    The second point is <X2>, <Y2>.
	--  Warning: Raises SegmentDefinitionError if the
	--	    first point and the second point are identical.
	raises SegmentDefinitionError from Graphic2d;

	----------------------------------------
	-- Category: Inquire methods
	----------------------------------------

	FirstPoint( me; X, Y: out Length from Quantity );  
	---Level: Public
	---Purpose: returns the coordinates of the first point of the segment
	
	SecondPoint( me; X, Y: out Length from Quantity );  
	---Level: Public
	---Purpose: returns the coordinates of the second point of the segment
	
	--------------------------------------
	-- Category: Draw and Pick
	--------------------------------------

	Draw (me : mutable; aDrawer: Drawer from Graphic2d)
	is static protected;
	---Level: Internal
	---Purpose: Draws the segment <me>.

	DrawElement( me : mutable; aDrawer: Drawer from Graphic2d;
		 anIndex: Integer from Standard)
	is redefined protected;
	---Level: Internal
	---Purpose: Draws edge <anIndex> of the segment <me>.

	DrawVertex( me : mutable; aDrawer: Drawer from Graphic2d;
		anIndex: Integer from Standard)
	is redefined protected;
	---Level: Internal
	---Purpose: Draws vertex <anIndex> of the segment <me>.

	Pick (me : mutable; X, Y: ShortReal from Standard;
		aPrecision: ShortReal from Standard;
		aDrawer: Drawer from Graphic2d)
	returns Boolean from Standard
	is static protected;
	---Level: Internal
	---Purpose: Returns Standard_True if the segment <me> is picked,
	--	    Standard_False if not.

	----------------------------------------------------------------------

	Save(me; aFStream: in out FStream from Aspect) is virtual;
	Retrieve(myclass; anIFStream: in out IFStream from Aspect;
		aGraphicObject: GraphicObject from Graphic2d);

fields

	myX1:	ShortReal from Standard;
	myY1:	ShortReal from Standard;
	myX2:	ShortReal from Standard;
	myY2:	ShortReal from Standard;

end Segment from Graphic2d;
