-- Created on: 1992-02-03
-- Created by: Christian CAILLET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package Transfer

    ---Purpose : Defines general Transfer engine, which provides tools and
    --           workframe for all kinds of file (non-direct) Interfaces.
    --           Works on the basis of data provided by package Interface
    --           (especially InterfaceModel).

uses TCollection, TColStd, MMgt, Standard, Dico, MoniTool, Interface,  Message

is

    class DataInfo;  -- used in Mapper

    deferred class Finder;
    	generic class Mapper;
	class TransientMapper  instantiates Mapper
    	    (Transient, MapTransientHasher from TColStd, DataInfo);
    class FindHasher;

    deferred class Binder;
    	class VoidBinder;
    	generic class SimpleBinder;
    	class SimpleBinderOfTransient;
	class BinderOfTransientInteger;
        class TransientListBinder;
    	class MultipleBinder;

    class ResultFromTransient;
    class ResultFromModel;

    class TransferIterator;
    generic class TransferProcess;
    generic class TransferMap;
    generic class Iterator;
    generic class Actor;

    class ProcessForTransient   instantiates TransferProcess
    	(Transient,  MapTransientHasher from TColStd,
    	 HSequenceOfTransient  from TColStd);
    ---Purpose : Manages Transfer of Transient Objects. Produces also
    --           ActorOfTransientProcess       (deferred class),
    --           IteratorOfTransientProcess    (for Results),
    --           TransferMapOfTransientProcess (internally used)
    --           Normally uses as TransientProcess, which adds some specifics

    class TransientProcess;    -- inherits TransferForTransient
    class ActorOfTransientProcess;

    class SequenceOfFinder instantiates
    	 Sequence from TCollection (Finder);
    class HSequenceOfFinder instantiates
    	HSequence from TCollection (Finder,SequenceOfFinder);

    class ProcessForFinder      instantiates TransferProcess
    	(Finder,     FindHasher,   HSequenceOfFinder);

    class FinderProcess;
    class ActorOfFinderProcess;

    class TransferOutput;
    class TransferInput;

    class DispatchControl;
    class TransferDispatch;
    class ActorDispatch;
    
    class MapContainer;

    class SequenceOfBinder instantiates
    	 Sequence from TCollection (Binder);
    class HSequenceOfBinder instantiates
    	HSequence from TCollection (Binder,SequenceOfBinder);

    enumeration StatusResult is  StatusVoid, StatusDefined, StatusUsed;
    ---Purpose : result status of transferring an entity (see Transcriptor)

    enumeration StatusExec is
    	StatusInitial, StatusRun, StatusDone, StatusError,StatusLoop;
    ---Purpose : execution status of an individual transfer (see Transcriptor)

    enumeration UndefMode is
    	UndefIgnore, UndefFailure, UndefContent, UndefUser;
    ---Purpose : used on processing Undefined Entities (see TransferOutput)

    	-- --  Exceptions  -- --

    exception TransferFailure   inherits InterfaceError  from Interface;
    exception TransferDeadLoop  inherits TransferFailure from Transfer;

end Transfer;
