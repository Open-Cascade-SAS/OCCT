-- Created on: 1996-08-30
-- Created by: Yves FRICAUD
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Inter3d from BRepOffset 

	---Purpose: Computes the intersection face face in a set of faces
	--          Store the result in a SD as AsDes.

uses
    AsDes                     from BRepAlgo,
    Image                     from BRepAlgo,
    Analyse                   from BRepOffset,	
    DataMapOfShapeOffset      from BRepOffset,
    Shape                     from TopoDS,
    Face                      from TopoDS,
    ListOfShape               from TopTools,
    --MapOfShape                from TopTools,
    IndexedMapOfShape         from TopTools,
    DataMapOfShapeShape       from TopTools,
    DataMapOfShapeListOfShape from TopTools,
    Real                      from Standard,
    State                     from TopAbs	

is
    Create(AsDes : AsDes from BRepAlgo;
           Side  : State         from TopAbs;
    	   Tol   : Real          from Standard);
    
    CompletInt (me : in out; SetOfFaces     : ListOfShape from TopTools; 
    	    	    	     InitOffsetFace : Image       from BRepAlgo  ) 
    is static;

    FaceInter (me : in out; 
    	       F1, F2         : Face  from TopoDS;
    	       InitOffsetFace : Image from BRepAlgo) 
    is static;
    
    ConnexIntByArc(me : in out; 
    	          SetOfFaces     : ListOfShape from TopTools; 
    	          ShapeInit      : Shape       from TopoDS;
    	          Analyse        : Analyse     from BRepOffset;
    	    	  InitOffsetFace : Image       from BRepAlgo)
    is static;		  
    
    ConnexIntByInt(me     : in out;  
    	    	   SI     :        Shape                from TopoDS;
    	           MapSF  :        DataMapOfShapeOffset from BRepOffset;
		   A      :        Analyse              from BRepOffset;
		   MES    : in out DataMapOfShapeShape  from TopTools;
		   Build  : in out DataMapOfShapeShape  from TopTools;
		   Failed : in out ListOfShape          from TopTools)
    is static;
     
    ContextIntByInt( me             : in  out;   
                     ContextFaces   :        IndexedMapOfShape    from TopTools; 
		     ExtentContext  :        Boolean              from Standard;	
    	             MapSF          :        DataMapOfShapeOffset from BRepOffset;
		     A              :        Analyse              from BRepOffset;
		     MES            : in out DataMapOfShapeShape  from TopTools;
		     Build          : in out DataMapOfShapeShape  from TopTools;
		     Failed         : in out ListOfShape          from TopTools) 
    is  static; 
     
    ContextIntByArc(me : in out;
    	      	    ContextFaces   :        IndexedMapOfShape from TopTools;
    	    	    ExtentContext  :        Boolean           from Standard;	
    	       	    Analyse        :        Analyse           from BRepOffset;
    	      	    InitOffsetFace :        Image             from BRepAlgo;
    	       	    InitOffsetEdge : in out Image             from BRepAlgo)
    is static;	       	
    
    AddCommonEdges(me : in out; 
    	    	   SetOfFaces : ListOfShape from TopTools)
    is static;		   
    
    SetDone(me : in out; F1,F2 : Face from TopoDS)
    is static;
    
   ---Category: Querying

    IsDone(me ; F1,F2 : Face from TopoDS) 
    returns Boolean from Standard
    is static;
    
    TouchedFaces(me : in out) returns IndexedMapOfShape from TopTools
	---C++: return &
    is static;
    
    AsDes(me) returns AsDes from BRepAlgo
    is static;
    
    NewEdges(me : in out) returns IndexedMapOfShape from TopTools
    	---C++:  return &
    is static;
    
    ---Category: Private

    Store(me : in out;F1,F2       : Face        from TopoDS;
    	              LInt1,LInt2 : ListOfShape from TopTools)
    is static private;    
    
fields

   myAsDes        : AsDes                     from BRepAlgo;
   myTouched      : IndexedMapOfShape         from TopTools;
   myDone         : DataMapOfShapeListOfShape from TopTools;
   myNewEdges     : IndexedMapOfShape         from TopTools;
   mySide         : State                     from TopAbs;
   myTol          : Real                      from Standard;
   
end Inter3d;
