-- File:	RWStepVisual_RWDraughtingModel.cdl
-- Created:	Thu Jan 13 10:08:42 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0
-- Copyright:	Matra Datavision 1999

class RWDraughtingModel from RWStepVisual

    ---Purpose: Read & Write tool for DraughtingModel

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    DraughtingModel from StepVisual

is
    Create returns RWDraughtingModel from RWStepVisual;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : DraughtingModel from StepVisual);
	---Purpose: Reads DraughtingModel

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: DraughtingModel from StepVisual);
	---Purpose: Writes DraughtingModel

    Share (me; ent : DraughtingModel from StepVisual;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWDraughtingModel;
