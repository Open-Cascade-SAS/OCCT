-- File:	LocOpe_CurveShapeIntersector.cdl
-- Created:	Mon May 29 15:54:11 1995
-- Author:	Jacques GOUSSARD
--		<jag@bravox>
---Copyright:	 Matra Datavision 1995


class CurveShapeIntersector from LocOpe

	---Purpose: This  class  provides  the intersection between an
	--          axis  or  a circle and  the  faces of a shape. The
	--          intersection   points  are   sorted in  increasing
	--          parameter along the axis.


uses SequenceOfPntFace from LocOpe,
     PntFace           from LocOpe,
     Shape             from TopoDS,
     Face              from TopoDS,
     Orientation       from TopAbs,
     Ax1               from gp,
     Circ              from gp

raises NotDone    from StdFail,
       OutOfRange from Standard

is

    Create
	---Purpose: Empty constructor.
    	returns CurveShapeIntersector from LocOpe;
	---C++: inline


    Create(Axis: Ax1 from gp; S:Shape from TopoDS)
	---Purpose: Creates  and performs the intersection     betwwen
	--          <Ax1> and <S>.
	---C++: inline
    	returns CurveShapeIntersector from LocOpe;


    Create(C: Circ from gp; S:Shape from TopoDS)
	---Purpose: Creates  and performs yte intersection     betwwen
	--          <C> and <S>.
	---C++: inline
    	returns CurveShapeIntersector from LocOpe;


    Init(me: in out;Axis: Ax1 from gp; S:Shape from TopoDS)
	---Purpose: Performs the intersection between <Ax1 and <S>.
	is static;


    Init(me: in out;C: Circ from gp; S:Shape from TopoDS)
	---Purpose: Performs the intersection between <Ax1 and <S>.
	is static;


    IsDone(me)
	---Purpose: Returns <Standard_True>  if the  intersection  has
	--          been done.
    	returns Boolean from Standard
	---C++: inline
	is static;


    NbPoints(me)
	---Purpose: Returns the number of intersection point.
    	returns Integer from Standard
	---C++: inline
	raises NotDone from StdFail
	-- The exception is raised when IsDone returns <Standard_False>.
	is static;


    Point(me; Index: Integer from Standard)
    
	---Purpose: Returns the intersection  point  of range <Index>.
	--          The points  are   sorted in increasing  order   of
	--          parameter along the axis. 

    	returns PntFace from LocOpe
	---C++: return const&
	---C++: inline
	raises NotDone    from StdFail,
	       OutOfRange from Standard
	is static;


    LocalizeAfter(me; From    : Real from Standard;
		      Or      : out Orientation from TopAbs; 
                      IndFrom : out Integer from Standard;
		      IndTo   : out Integer from Standard)
    
	---Purpose: Searches the   first intersection  point   located
	--          after the  parameter  <From>, wich  orientation is
	--          not       TopAbs_EXTERNAL.      If found,  returns
	--          <Standard_True>.  <Or> contains the orientation of
	--          the  point, <IndFrom>  and  <IndTo> represents the
	--          interval of index  in the sequence of intersection
	--          point  corresponding  to   the point. (IndFrom  <=
	--          IndTo). 
	--          
	--          Otherwise, returns <Standard_False>.
    	
    	returns Boolean from Standard
    	raises NotDone from StdFail
	is static;


    LocalizeBefore(me; From    : Real from Standard;
		       Or      : out Orientation from TopAbs; 
                       IndFrom : out Integer from Standard;
		       IndTo   : out Integer from Standard)
    
	---Purpose: Searches  the first intersection point     located
	--          before  the parameter <From>,  wich orientation is
	--          not      TopAbs_EXTERNAL.      If  found,  returns
	--          <Standard_True>.  <Or> contains the orientation of
	--          the point,  <IndFrom>  and <IndTo>  represents the
	--          interval of index  in the sequence of intersection
	--          point  corresponding   to the point   (IndFrom  <=
	--          IndTo). 
	--          
	--          Otherwise, returns <Standard_False>.
    	
    	returns Boolean from Standard
    	raises NotDone from StdFail
	is static;


    LocalizeAfter(me; FromInd : Integer from Standard;
		      Or      : out Orientation from TopAbs; 
                      IndFrom : out Integer from Standard;
		      IndTo   : out Integer from Standard)
    
	---Purpose: Searches  the first intersection point     located
	--          after the index <FromInd>  ( >= FromInd + 1), wich
	--          orientation   is   not TopAbs_EXTERNAL.   If found,
	--          returns   <Standard_True>.   <Or>  contains    the
	--          orientation of the  point, <IndFrom>  and  <IndTo>
	--          represents the interval  of index in  the sequence
	--          of  intersection  point     corresponding to   the
	--          point. (IndFrom <= IndTo).
	--          
	--          Otherwise, returns <Standard_False>.
    	
    	returns Boolean from Standard
    	raises NotDone from StdFail
	is static;


    LocalizeBefore(me; FromInd : Integer from Standard;
		       Or      : out Orientation from TopAbs; 
                       IndFrom : out Integer from Standard;
		       IndTo   : out Integer from Standard)
    
	---Purpose: Searches the  first  intersection   point  located
	--          before the index <FromInd>  ( <= FromInd -1), wich
	--          orientation is   not TopAbs_EXTERNAL.   If   found,
	--          returns   <Standard_True>.  <Or>  contains     the
	--          orientation  of the  point,  <IndFrom> and <IndTo>
	--          represents the interval  of index  in the sequence
	--          of  intersection  point corresponding to the point
	--          (IndFrom <= IndTo).
	--          
	--          Otherwise, returns <Standard_False>.
    	
    	returns Boolean from Standard
    	raises NotDone from StdFail
	is static;

fields

    myDone   : Boolean           from Standard;
    myPoints : SequenceOfPntFace from LocOpe;

end CurveShapeIntersector;
