-- File:	BSplCLib.cdl
-- Created:	Fri Aug  9 15:12:53 1991
-- Author:	Jean Claude VAUTHIER
---Copyright:	 Matra Datavision 1991, 1992
--           	 
--Modified : RLE Aug   1993  Major modifications.  
--  15-Mar-95  xab : added cache mecanism to speed up 
--  evaluation
--  25-Mar-95  xab : added Lagrange evaluator
-- mei : modified 08-Jun-95 : added method MovePoint
-- xab : modified 11-Mar-96 : added method MovePointAndTangent
-- xab : modified 18-Mar-97 : added method to reparameterise a bspline 
-- jct : modified 15-Apr-97 : added method to extend a bspline 

package BSplCLib

    ---Purpose:  BSplCLib   B-spline curve Library.
    --  
    --  The BSplCLib package is  a basic library  for BSplines. It
    --  provides three categories of functions.
    --  
    --  * Management methods to  process knots and multiplicities.
    --  
    --  * Multi-Dimensions  spline methods.  BSpline methods where
    --  poles have an arbitrary number of dimensions. They divides
    --  in two groups :
    --  
    --    - Global methods modifying the  whole set of  poles. The
    --    poles are    described   by an array   of   Reals and  a
    --    Dimension. Example : Inserting knots.
    --    
    --    - Local methods  computing  points and derivatives.  The
    --    poles  are described by a pointer  on  a local array  of
    --    Reals and a Dimension. The local array is modified.
    --  
    --  *  2D  and 3D spline   curves  methods.
    --  
    --    Methods  for 2d and 3d BSplines  curves  rational or not
    --    rational. 
    --    
    --    Those methods have the following structure :
    --    
    --     - They extract the pole informations in a working array.
    --     
    --     -  They      process the  working   array    with   the
    --     multi-dimension  methods. (for example  a  3d  rational
    --     curve is processed as a 4 dimension curve).
    --     
    --     - They get back the result in the original dimension.
    --     
    --     Note that the  bspline   surface methods found   in the
    --     package BSplSLib  uses  the same  structure and rely on
    --     BSplCLib.
    --     
    --     In the following list  of methods the  2d and 3d  curve
    --     methods   will be  described   with  the  corresponding
    --     multi-dimension method.
    --  
    --  The 3d or 2d B-spline curve is defined with :
    --  
    --  . its control points : TColgp_Array1OfPnt(2d)        Poles
    --  . its weights        : TColStd_Array1OfReal          Weights
    --  . its knots          : TColStd_Array1OfReal          Knots 
    --  . its multiplicities : TColStd_Array1OfInteger       Mults
    --  . its degree         : Standard_Integer              Degree
    --  . its periodicity    : Standard_Boolean              Periodic   
    --
    -- Warnings :
    --  The bounds of Poles and Weights should be the same.
    --  The bounds of Knots and Mults   should be the same.
    --  
    --  Weights can be a null reference (BSplCLib::NoWeights())
    --  the curve is non rational.
    --  
    --  Mults can be a null reference   (BSplCLib::NoMults())
    --  the knots are "flat" knots.
    --  
    -- KeyWords :
    --  B-spline curve, Functions, Library
    --  
    -- References :
    --  . A survey of curves and surfaces methods in CADG Wolfgang 
    --    BOHM CAGD 1 (1984)
    --  . On de Boor-like algorithms and blossoming Wolfgang BOEHM
    --    cagd 5 (1988)
    --  . Blossoming and knot insertion algorithms for B-spline curves
    --    Ronald N. GOLDMAN
    --  . Modelisation des surfaces en CAO, Henri GIAUME Peugeot SA   
    --  . Curves and Surfaces for Computer Aided Geometric Design,
    --    a practical guide Gerald Farin

uses TColStd, gp, TColgp, math


is

    imported EvaluatorFunction ;
    ---Purpose: this is a one dimensional function 
    --  typedef  void (*EvaluatorFunction)  (
    --  Standard_Integer     // Derivative Request
    --  Standard_Real    *   // StartEnd[2] 
    --  Standard_Real        // Parameter
    --  Standard_Real    &   // Result
    --  Standard_Integer &) ;// Error Code
    --  serves to multiply a given vectorial BSpline by a function 

    enumeration KnotDistribution is NonUniform, Uniform;
    ---Purpose: This enumeration describes the repartition of the
    --         knots  sequence.   If all the knots  differ  by the
    --         same positive constant from the  preceding knot the
    --         "KnotDistribution" is    <Uniform>    else   it  is
    --         <NonUniform>

    enumeration MultDistribution is NonConstant, Constant, QuasiConstant;
    ---Purpose:  This   enumeration describes the   form  of  the
    --         sequence of mutiplicities.  MultDistribution is :
    --          
    --            Constant if all the multiplicities have the same
    --            value.
    --          
    --            QuasiConstant if all the internal knots have the
    --            same multiplicity and if the first and last knot
    --            have  a different  multiplicity.  
    --            
    --            NonConstant in other cases.

    	-------------------------------------------------------------
    	-------------------------------------------------------------
    	----------					   ----------
    	----------	    Knots and Multiplicities	   ----------
    	----------					   ----------
    	-------------------------------------------------------------
    	-------------------------------------------------------------

    Hunt (XX   : in Array1OfReal from TColStd;
    	  X    : in Real;
    	  Iloc : in out Integer);
    ---Purpose:  This routine searches the position of the real
    --         value X in  the ordered set of  real  values XX.
    --         
    --         The  elements   in   the  table    XX  are   either
    --         monotonically    increasing     or    monotonically
    --         decreasing.
    --         
    --         The input   value Iloc is    used to initialize the
    --         algorithm  :  if  Iloc  is outside  of   the bounds
    --         [XX.Lower(), -- XX.Upper()] the bisection algorithm
    --         is used else  the routine searches from  a previous
    --         known position  by increasing steps  then converges
    --         by bisection.
    --         
    --         This  routine is used to  locate a  knot value in a
    --         set of knots.
    --         
    ---References : Numerical Recipes in C (William H.Press, Brian
    --            P.  Flannery,  Saul   A.  Teukolsky, William  T.
    --            Vetterling)

    FirstUKnotIndex (Degree : Integer;
    	    	     Mults  : Array1OfInteger from TColStd)
    returns Integer;
    ---Purpose: Computes the index of the knots value which gives
    --         the start point of the curve.
     

    LastUKnotIndex (Degree : Integer;
    	    	    Mults  : Array1OfInteger from TColStd)
    returns Integer;
    ---Purpose: Computes the index of the knots value which gives
    --         the end point of the curve.
     
    FlatIndex (Degree : Integer;
     	       Index  : Integer;
	       Mults  : Array1OfInteger from TColStd;
	       Periodic : Boolean)
    returns Integer;
    ---Purpose: Computes the index  of  the  flats knots  sequence
    --          corresponding  to  <Index> in  the  knots sequence
    --          which multiplicities are <Mults>.
     
    LocateParameter (Degree     : Integer; 
                     Knots      : Array1OfReal from TColStd; 
                     Mults      : Array1OfInteger from TColStd;
                     U          : Real; 
                     IsPeriodic : Boolean;
		     FromK1     : Integer;
		     ToK2       : Integer;
                     KnotIndex  : in out Integer;
                     NewU       : in out Real);
    ---Purpose:  Locates  the parametric value    U  in the knots
    --         sequence  between  the  knot K1   and the knot  K2.
    --         The value return in Index verifies.
    --  
    --          Knots(Index) <= U < Knots(Index + 1)
    --          if U <= Knots (K1) then Index = K1
    --          if U >= Knots (K2) then Index = K2 - 1
    --          
    --          If Periodic is True U  may be  modified  to fit in
    --          the range  Knots(K1), Knots(K2).  In any case  the
    --          correct value is returned in NewU.
    --  
    --  Warnings :Index is used  as input   data to initialize  the
    --          searching  function.
    --  Warning: Knots have to be "withe repetitions"
		     
    LocateParameter (Degree     : Integer; 
                     Knots      : Array1OfReal from TColStd; 
                     U          : Real; 
                     IsPeriodic : Boolean;
		     FromK1     : Integer;
		     ToK2       : Integer;
                     KnotIndex  : in out Integer;
                     NewU       : in out Real);
    ---Purpose:  Locates  the parametric value    U  in the knots
    --         sequence  between  the  knot K1   and the knot  K2.
    --         The value return in Index verifies.
    --  
    --          Knots(Index) <= U < Knots(Index + 1)
    --          if U <= Knots (K1) then Index = K1
    --          if U >= Knots (K2) then Index = K2 - 1
    --          
    --          If Periodic is True U  may be  modified  to fit in
    --          the range  Knots(K1), Knots(K2).  In any case  the
    --          correct value is returned in NewU.
    --  
    --  Warnings :Index is used  as input   data to initialize  the
    --          searching  function.
    --  Warning: Knots have to be "flat"

    LocateParameter (Knots    : Array1OfReal from TColStd; 
                     U        : Real; 
                     Periodic : Boolean;
		     K1,K2    : Integer;
                     Index    : in out Integer;
                     NewU     : in out Real;
                     Uf,Ue    : Real)
    is private;     
    ---Level: Internal	
		   
    LocateParameter (Degree   : Integer;
    	    	     Knots    : Array1OfReal    from TColStd; 
    	             Mults    : Array1OfInteger from TColStd;
                     U        : Real; 
                     Periodic : Boolean;
                     Index    : in out Integer;
                     NewU     : in out Real);
    ---Level: Internal

    MaxKnotMult (Mults  : Array1OfInteger from TColStd;
    	         K1, K2 : Integer)
    returns Integer;  
    ---Purpose: Finds the greatest multiplicity in a set of knots
    --         between  K1  and K2.   Mults  is  the  multiplicity
    --         associated with each knot value.

    MinKnotMult (Mults  : Array1OfInteger from TColStd;
    	         K1, K2 : Integer)
    returns Integer;  
    ---Purpose: Finds the lowest multiplicity in  a  set of knots
    --         between   K1  and K2.   Mults is  the  multiplicity
    --         associated with each knot value.

    NbPoles(Degree   : Integer;
    	    Periodic : Boolean;
	    Mults    : Array1OfInteger from TColStd) 
    returns Integer;
    ---Purpose: Returns the number of poles of the curve. Returns 0 if
    --          one of the multiplicities is incorrect.
    --          
    --          * Non positive.
    --          
    --          * Greater than Degree,  or  Degree+1  at the first and
    --          last knot of a non periodic curve.
    --          
    --          *  The  last periodicity  on  a periodic  curve is not
    --          equal to the first.

    KnotSequenceLength(Mults    : Array1OfInteger from TColStd;
    	    	       Degree   : Integer;
    	    	       Periodic : Boolean)
    returns Integer;
    ---Purpose: Returns the length  of the sequence  of knots with
    --          repetition.
    --          
    --          Periodic :
    --          
    --          Sum(Mults(i), i = Mults.Lower(); i <= Mults.Upper());
    --          
    --          Non Periodic :
    --          
    --          Sum(Mults(i); i = Mults.Lower(); i < Mults.Upper())
    --          + 2 * Degree

    KnotSequence (Knots    : Array1OfReal from TColStd; 
                  Mults    : Array1OfInteger from TColStd;
                  KnotSeq  : in out Array1OfReal from TColStd);
		
    KnotSequence (Knots    : Array1OfReal from TColStd; 
                  Mults    : Array1OfInteger from TColStd;
		  Degree   : Integer;
		  Periodic : Boolean;
                  KnotSeq  : in out Array1OfReal from TColStd);
    ---Purpose: Computes  the  sequence   of knots KnotSeq  with
    --         repetition  of the  knots  of multiplicity  greater
    --         than 1.
    --  
    --  Length of KnotSeq must be KnotSequenceLength(Mults,Degree,Periodic)

    KnotsLength( KnotSeq  :  Array1OfReal from TColStd; 
                 Periodic  :  Boolean  =  Standard_False) 
    returns  Integer; 
    ---Purpose: Returns the  length  of the   sequence of  knots  (and
    --          Mults)  without repetition.
           
    Knots( KnotSeq  :  Array1OfReal from TColStd; 
    	   Knots    :  out Array1OfReal from TColStd; 
	   Mults    :  out Array1OfInteger from TColStd; 
           Periodic  :  Boolean  =  Standard_False);
    ---Purpose:  Computes  the  sequence   of knots Knots  without
    --         repetition  of the  knots  of multiplicity  greater
    --         than 1.
    --  
    --       Length  of <Knots> and  <Mults> must be 
    --    KnotsLength(KnotSequence,Periodic)

    KnotForm  (Knots : Array1OfReal from TColStd;
    	       FromK1, ToK2 : Integer)
    returns KnotDistribution;
    ---Purpose: Analyses if the  knots distribution is "Uniform"
    --         or  "NonUniform" between  the  knot  FromK1 and the
    --         knot ToK2.  There is  no repetition of  knot in the
    --         knots'sequence <Knots>.

    MultForm  (Mults : Array1OfInteger from TColStd;
    	       FromK1, ToK2 : Integer)
    returns MultDistribution;
    ---Purpose:
    --  Analyses the distribution of multiplicities between
    --  the knot FromK1 and the Knot ToK2.

    Reparametrize (U1, U2 : Real;
    	    	   Knots : in out Array1OfReal from TColStd);
    ---Purpose:
    --  Reparametrizes a B-spline curve to [U1, U2].
    --  The knot values are recomputed such that Knots (Lower) = U1
    --  and Knots (Upper) = U2   but the knot form is not modified. 
    --   Warnings :
    --  In the array Knots the values must be in ascending order.
    --  U1 must not be equal to U2 to avoid division by zero.


    Reverse (Knots : in out Array1OfReal from TColStd);
    ---Purpose: Reverses  the  array   knots  to  become  the knots
    --          sequence of the reversed curve. 
	
    Reverse (Mults : in out Array1OfInteger from TColStd);
    ---Purpose: Reverses  the  array of multiplicities.
	
    Reverse (Poles    : in out Array1OfPnt  from TColgp;
    	     Last     : Integer);
    ---Purpose: Reverses the array of poles. Last is the  index of
    --          the new first pole. On  a  non periodic curve last
    --          is Poles.Upper(). On a periodic curve last is 
    --          
    --          (number of flat knots - degree - 1) 
    --          
    --          or
    --          
    --          (sum of multiplicities(but  for the last) + degree
    --          - 1)

    Reverse (Poles    : in out Array1OfPnt2d  from TColgp;
    	     Last     : Integer);
    ---Purpose: Reverses the array of poles.

    Reverse (Weights  : in out Array1OfReal  from TColStd;
    	     Last     : Integer);
    ---Purpose: Reverses the array of poles.

    IsRational(Weights : Array1OfReal from TColStd;
    	       I1,I2   : Integer;
    	       Epsilon : Real = 0.0) returns Boolean;
    ---Purpose: 
    --   Returns False if all the weights  of the  array <Weights>
    --   between   I1 an I2   are  identic.   Epsilon  is used for
    --   comparing  weights. If Epsilon  is 0. the  Epsilon of the
    --   first weight is used.

    MaxDegree  returns Integer;
    ---Purpose: returns the degree maxima for a BSplineCurve.
    ---C++: inline

    Eval(U         : Real;
    	 Degree    : Integer;
    	 Knots     : in out Real;
	 Dimension : Integer;
	 Poles     : in out Real);
    ---Purpose: Perform the Boor  algorithm  to  evaluate a point at
    --          parameter <U>, with <Degree> and <Dimension>.
    --          
    --          Poles is  an array of  Reals of size 
    --          
    --          <Dimension> *  <Degree>+1
    --          
    --          Containing  the poles.  At  the end <Poles> contains
    --          the current point.

    BoorScheme(U         : Real;
    	       Degree    : Integer;
    	       Knots     : in out Real;
	       Dimension : Integer;
	       Poles     : in out Real;
	       Depth     : Integer;
	       Length    : Integer);
    ---Purpose: Performs the  Boor Algorithm  at  parameter <U> with
    --          the given <Degree> and the  array of <Knots> on  the
    --          poles <Poles> of dimension  <Dimension>.  The schema
    --          is  computed  until  level  <Depth>  on a   basis of
    --          <Length+1> poles.
    --          
    --          * Knots is an array of reals of length :
    --          
    --            <Length> + <Degree>
    --          
    --          * Poles is an array of reals of length :
    --          
    --           (2 * <Length> + 1) * <Dimension> 
    --           
    --           The poles values  must be  set  in the array at the
    --           positions. 
    --           
    --            0..Dimension, 
    --            
    --            2 * Dimension ..  
    --            3 * Dimension
    --            
    --            4  * Dimension ..  
    --            5  * Dimension
    --            
    --            ...
    --            
    --            The results are found in the array poles depending
    --            on the Depth. (See the method GetPole).

    AntiBoorScheme(U         : Real;
    	    	   Degree    : Integer;
    	           Knots     : in out Real;
	           Dimension : Integer;
	           Poles     : in out Real;
	           Depth     : Integer;
	           Length    : Integer;
    	    	   Tolerance : Real) returns Boolean;
    ---Purpose: Compute  the content of  Pole before the BoorScheme.
    --          This method is used to remove poles. 
    --          
    --          U is the poles to  remove, Knots should contains the
    --          knots of the curve after knot removal.
    --          
    --          The first  and last poles  do not  change, the other
    --          poles are computed by averaging two possible values.
    --          The distance between  the  two   possible  poles  is
    --          computed, if it  is higher than <Tolerance> False is
    --          returned.

    Derivative(Degree    : Integer;
    	       Knots     : in out Real;
	       Dimension : Integer;
	       Length    : Integer;
	       Order     : Integer;
	       Poles     : in out Real);
    ---Purpose: Computes   the   poles of  the    BSpline  giving the
    --          derivatives of order <Order>.
    --          
    --          The formula for the first order is
    --          
    --          Pole(i) = Degree * (Pole(i+1) - Pole(i)) / 
    --                             (Knots(i+Degree+1) - Knots(i+1))
    --                             
    --          This formula  is repeated  (Degree  is decremented at
    --          each step).

    Bohm(U         : Real;
    	 Degree    : Integer;
	 N         : Integer;
    	 Knots     : in out Real;
	 Dimension : Integer;
	 Poles     : in out Real);
    ---Purpose: Performs the Bohm  Algorithm at  parameter <U>. This
    --          algorithm computes the value and all the derivatives
    --          up to order N (N <= Degree).
    --          
    --          <Poles> is the original array of poles.
    --          
    --          The   result in  <Poles>  is    the value and    the
    --          derivatives.  Poles[0] is  the value,  Poles[Degree]
    --          is the last  derivative.

    
    NoWeights returns Array1OfReal from TColStd;
    ---Purpose: Used as argument for a non rational curve.
    --          
    ---C++: return &
    ---C++: inline
    
    NoMults  returns Array1OfInteger from TColStd;
    ---Purpose: Used as argument for a flatknots evaluation.
    --          
    ---C++: return &
    ---C++: inline

    BuildKnots(Degree, Index : Integer;
    	       Periodic   : Boolean;
               Knots      : Array1OfReal    from TColStd;
    	       Mults      : Array1OfInteger from TColStd;
    	       LK         : in out Real);
    ---Purpose: Stores in LK  the usefull knots  for the BoorSchem
    --          on the span Knots(Index) - Knots(Index+1)
	  
    PoleIndex (Degree, Index : Integer;
    	       Periodic   : Boolean;
    	       Mults      : Array1OfInteger from TColStd)
    returns Integer;
    ---Purpose: Return the index of the  first Pole to  use on the
    --          span  Mults(Index)  - Mults(Index+1).  This  index
    --          must be added to Poles.Lower().
	  
    BuildEval(Degree,Index : Integer;
              Poles      : Array1OfReal    from TColStd;
    	      Weights    : Array1OfReal    from TColStd;
              LP         : in out Real);

    BuildEval(Degree,Index : Integer;
              Poles      : Array1OfPnt     from TColgp;
    	      Weights    : Array1OfReal    from TColStd;
              LP         : in out Real);

    BuildEval(Degree,Index : Integer;
              Poles      : Array1OfPnt2d   from TColgp;
    	      Weights    : Array1OfReal    from TColStd;
              LP         : in out Real);
    ---Purpose: Copy in <LP>  the poles and  weights for  the Eval
    --          scheme. starting from  Poles(Poles.Lower()+Index)

    BuildBoor(Index,Length,Dimension : Integer;
    	      Poles      : Array1OfReal    from TColStd;
              LP         : in out Real);
    ---Purpose: Copy in <LP>  poles for <Dimension>  Boor  scheme.
    --          Starting  from    <Index>     *  <Dimension>, copy
    --          <Length+1> poles.


    BoorIndex(Index, Length, Depth : Integer)
    returns Integer;
    ---Purpose: Returns the index in  the Boor result array of the
    --          poles <Index>. If  the Boor  algorithm was perform
    --          with <Length> and <Depth>.

    GetPole(Index,Length,Depth,Dimension : Integer;
   	    LocPoles : in out Real;
	    Position : in out Integer;
            Pole     : in out Array1OfReal from TColStd);
    ---Purpose: Copy  the  pole at  position  <Index>  in  the Boor
    --          scheme of   dimension <Dimension> to  <Position> in
    --          the array <Pole>. <Position> is updated.

    PrepareInsertKnots (
     Degree     : in Integer; 
     Periodic   : in Boolean;
     Knots      : in Array1OfReal    from TColStd;
     Mults      : in Array1OfInteger from TColStd;
     AddKnots   : in Array1OfReal    from TColStd;
     AddMults   : in Array1OfInteger from TColStd;
     NbPoles    : out Integer;
     NbKnots    : out Integer;
     Epsilon    : in Real;
     Add        : in Boolean = Standard_True) 
    returns Boolean;
    ---Purpose: Returns in <NbPoles, NbKnots> the  new number of poles
    --          and  knots    if  the  sequence   of  knots <AddKnots,
    --          AddMults> is inserted in the sequence <Knots, Mults>.
    --          
    --          Epsilon is used to compare knots for equality.
    --          
    --          If Add is True  the multiplicities on  equal knots are
    --          added. 
    --          
    --          If Add is False the max value of the multiplicities is
    --          kept. 
    --          
    --          Return False if :
    --            The knew knots are knot increasing.
    --            The new knots are not in the range.

    InsertKnots (
     Degree     : in Integer; 
     Periodic   : in Boolean;
     Dimension  : in Integer;
     Poles      : in Array1OfReal     from TColStd;
     Knots      : in Array1OfReal     from TColStd;
     Mults      : in Array1OfInteger  from TColStd;
     AddKnots   : in Array1OfReal     from TColStd;
     AddMults   : in Array1OfInteger  from TColStd;
     NewPoles   : out Array1OfReal    from TColStd;
     NewKnots   : out Array1OfReal    from TColStd;
     NewMults   : out Array1OfInteger from TColStd;
     Epsilon    : in Real;
     Add        : in Boolean = Standard_True);
    
    InsertKnots (
     Degree     : in Integer; 
     Periodic   : in Boolean;
     Poles      : in Array1OfPnt      from TColgp;
     Weights    : in Array1OfReal     from TColStd;
     Knots      : in Array1OfReal     from TColStd;
     Mults      : in Array1OfInteger  from TColStd;
     AddKnots   : in Array1OfReal     from TColStd;
     AddMults   : in Array1OfInteger  from TColStd;
     NewPoles   : out Array1OfPnt     from TColgp;
     NewWeights : out Array1OfReal    from TColStd;
     NewKnots   : out Array1OfReal    from TColStd;
     NewMults   : out Array1OfInteger from TColStd;
     Epsilon    : in Real;
     Add        : in Boolean = Standard_True);

    InsertKnots (
     Degree     : in Integer; 
     Periodic   : in Boolean;
     Poles      : in Array1OfPnt2d    from TColgp;
     Weights    : in Array1OfReal     from TColStd;
     Knots      : in Array1OfReal     from TColStd;
     Mults      : in Array1OfInteger  from TColStd;
     AddKnots   : in Array1OfReal     from TColStd;
     AddMults   : in Array1OfInteger  from TColStd;
     NewPoles   : out Array1OfPnt2d   from TColgp;
     NewWeights : out Array1OfReal    from TColStd;
     NewKnots   : out Array1OfReal    from TColStd;
     NewMults   : out Array1OfInteger from TColStd;
     Epsilon    : in Real;
     Add        : in Boolean = Standard_True);
    ---Purpose: Insert   a  sequence  of  knots <AddKnots> with
    --  multiplicities   <AddMults>. <AddKnots>   must  be a   non
    --  decreasing sequence and verifies :
    --  
    --  Knots(Knots.Lower()) <= AddKnots(AddKnots.Lower())
    --  Knots(Knots.Upper()) >= AddKnots(AddKnots.Upper())
    --  
    --  The NewPoles and NewWeights arrays must have a length :
    --    Poles.Length() + Sum(AddMults())
    --    
    --  When a knot  to insert is identic  to an existing knot the
    --  multiplicities   are added. 
    --  
    --  Epsilon is used to test knots for equality.
    --  
    --  When AddMult is negative or null the knot is not inserted.
    --  No multiplicity will becomes higher than the degree.
    --  
    --  The new Knots and Multiplicities  are copied in <NewKnots>
    --  and  <NewMults>. 
    --  
    --  All the New arrays should be correctly dimensioned.
    --  
    --  When all  the new knots  are existing knots, i.e. only the
    --  multiplicities  will  change it is   safe to  use the same
    --  arrays as input and output.

    InsertKnot (
     UIndex     : in Integer;
     U          : in Real; 
     UMult      : in Integer; 
     Degree     : in Integer; 
     Periodic   : in Boolean;
     Poles      : in Array1OfPnt     from TColgp;
     Weights    : in Array1OfReal    from TColStd;
     Knots      : in Array1OfReal    from TColStd;
     Mults      : in Array1OfInteger from TColStd;
     NewPoles   : out Array1OfPnt    from TColgp;
     NewWeights : out Array1OfReal   from TColStd);

    InsertKnot   (
     UIndex     : in Integer;
     U          : in Real;
     UMult      : in Integer; 
     Degree     : in Integer;
     Periodic   : in Boolean;
     Poles      : in Array1OfPnt2d   from TColgp;
     Weights    : in Array1OfReal    from TColStd;
     Knots      : in Array1OfReal    from TColStd; 
     Mults      : in Array1OfInteger from TColStd;
     NewPoles   : out Array1OfPnt2d  from TColgp;
     NewWeights : out Array1OfReal   from TColStd);
    ---Purpose: Insert a new knot U of multiplicity UMult in the
    --  knot sequence.
    --  
    --  The  location of the new Knot  should be given as an input
    --  data.  UIndex locates the new knot U  in the knot sequence
    --  and Knots (UIndex) < U < Knots (UIndex + 1).
    --  
    --  The new control points corresponding to this insertion are
    --  returned. Knots and Mults are not updated.
    
    RaiseMultiplicity (
     KnotIndex  : in Integer; 
     Mult       : in Integer;
     Degree     : in Integer;
     Periodic   : in Boolean;
     Poles      : in Array1OfPnt     from TColgp;
     Weights    : in Array1OfReal    from TColStd;
     Knots      : in Array1OfReal    from TColStd; 
     Mults      : in Array1OfInteger from TColStd; 
     NewPoles   : out Array1OfPnt    from TColgp;
     NewWeights : out Array1OfReal   from TColStd);

    RaiseMultiplicity (
     KnotIndex  : in Integer; 
     Mult       : in Integer;
     Degree     : in Integer;
     Periodic   : in Boolean;
     Poles      : in Array1OfPnt2d   from TColgp;
     Weights    : in Array1OfReal    from TColStd;
     Knots      : in Array1OfReal    from TColStd; 
     Mults      : in Array1OfInteger from TColStd; 
     NewPoles   : out Array1OfPnt2d  from TColgp;
     NewWeights : out Array1OfReal   from TColStd);
    ---Purpose: Raise the multiplicity of knot to <UMult>.
    --  
    --  The new control points  are  returned. Knots and Mults are
    --  not updated.

    RemoveKnot (
     Index      : in Integer;
     Mult       : in Integer; 
     Degree     : in Integer; 
     Periodic   : in Boolean;
     Dimension  : in Integer;
     Poles      : in Array1OfReal     from TColStd;
     Knots      : in Array1OfReal     from TColStd;
     Mults      : in Array1OfInteger  from TColStd;
     NewPoles   : out Array1OfReal    from TColStd;
     NewKnots   : out Array1OfReal    from TColStd;
     NewMults   : out Array1OfInteger from TColStd;
     Tolerance  : Real)  returns Boolean;
     
    RemoveKnot (
     Index      : in Integer;
     Mult       : in Integer; 
     Degree     : in Integer; 
     Periodic   : in Boolean;
     Poles      : in Array1OfPnt      from TColgp;
     Weights    : in Array1OfReal     from TColStd;
     Knots      : in Array1OfReal     from TColStd;
     Mults      : in Array1OfInteger  from TColStd;
     NewPoles   : out Array1OfPnt     from TColgp;
     NewWeights : out Array1OfReal    from TColStd;
     NewKnots   : out Array1OfReal    from TColStd;
     NewMults   : out Array1OfInteger from TColStd;
     Tolerance  : Real)  returns Boolean;

    RemoveKnot (
     Index      : in Integer;
     Mult       : in Integer; 
     Degree     : in Integer; 
     Periodic   : in Boolean;
     Poles      : in Array1OfPnt2d    from TColgp;
     Weights    : in Array1OfReal     from TColStd;
     Knots      : in Array1OfReal     from TColStd;
     Mults      : in Array1OfInteger  from TColStd;
     NewPoles   : out Array1OfPnt2d   from TColgp;
     NewWeights : out Array1OfReal    from TColStd;
     NewKnots   : out Array1OfReal    from TColStd;
     NewMults   : out Array1OfInteger from TColStd;
     Tolerance  : Real)  returns Boolean;
    ---Purpose: Decrement the  multiplicity  of <Knots(Index)>
    --          to <Mult>. If <Mult>   is  null the   knot  is
    --          removed. 
    --          
    --          As there are two ways to compute the new poles
    --          the midlle   will  be used  as  long    as the
    --          distance is lower than Tolerance.
    --          
    --          If a  distance is  bigger  than  tolerance the
    --          methods returns False  and  the new arrays are
    --          not modified.
    --          
    --          A low  tolerance can be  used  to test  if the
    --          knot  can be  removed  without  modifying  the
    --          curve. 
    --          
    --          A high tolerance  can be used  to "smooth" the 
    --          curve.
    
    
    IncreaseDegreeCountKnots (Degree, NewDegree : Integer;
    	    	    	      Periodic          : Boolean;
    	    	    	      Mults             : Array1OfInteger from TColStd)
    returns Integer;
    ---Purpose: Returns the   number   of  knots   of  a  curve   with
    --          multiplicities <Mults> after elevating the degree from
    --          <Degree> to <NewDegree>. See the IncreaseDegree method
    --          for more comments.

    IncreaseDegree  (Degree, 
    	    	     NewDegree   : in Integer;
		     Periodic    : in Boolean;
		     Dimension   : in Integer;
    	    	     Poles       : in Array1OfReal        from TColStd; 
    	    	     Knots       : in Array1OfReal        from TColStd; 
		     Mults       : in Array1OfInteger     from TColStd; 
		     NewPoles    : in out Array1OfReal    from TColStd;
    	    	     NewKnots    : in out Array1OfReal    from TColStd; 
		     NewMults    : in out Array1OfInteger from TColStd); 

    IncreaseDegree  (Degree, 
    	    	     NewDegree   : in Integer;
		     Periodic    : in Boolean;
    	    	     Poles       : in Array1OfPnt         from TColgp; 
		     Weights     : in Array1OfReal        from TColStd;
    	    	     Knots       : in Array1OfReal        from TColStd; 
		     Mults       : in Array1OfInteger     from TColStd; 
		     NewPoles    : in out Array1OfPnt     from TColgp; 
		     NewWeights  : in out Array1OfReal    from TColStd;
    	    	     NewKnots    : in out Array1OfReal    from TColStd; 
		    NewMults    : in out Array1OfInteger from TColStd); 

    IncreaseDegree  (Degree, 
    	    	     NewDegree   : in Integer;
		     Periodic    : in Boolean;
    	    	     Poles       : in Array1OfPnt2d       from TColgp; 
		     Weights     : in Array1OfReal        from TColStd;
    	    	     Knots       : in Array1OfReal        from TColStd; 
		     Mults       : in Array1OfInteger     from TColStd; 
		     NewPoles    : in out Array1OfPnt2d   from TColgp; 
		     NewWeights  : in out Array1OfReal    from TColStd;
    	    	     NewKnots    : in out Array1OfReal    from TColStd; 
		     NewMults    : in out Array1OfInteger from TColStd); 


    IncreaseDegree  (NewDegree   : in Integer;
    	    	     Poles       : in Array1OfPnt         from TColgp; 
		     Weights     : in Array1OfReal        from TColStd;
		     NewPoles    : in out Array1OfPnt     from TColgp; 
		     NewWeights  : in out Array1OfReal    from TColStd);
    ---Warning: To be used for Beziercurves ONLY!!!

    IncreaseDegree  (NewDegree   : in Integer;
    	    	     Poles       : in Array1OfPnt2d       from TColgp; 
		     Weights     : in Array1OfReal        from TColStd;
		     NewPoles    : in out Array1OfPnt2d   from TColgp; 
		     NewWeights  : in out Array1OfReal    from TColStd);
    ---Purpose: Increase the degree of a bspline (or bezier) curve
    --          of   dimension  <Dimension>  form <Degree>      to
    --          <NewDegree>.
    --          
    --          The number of poles in the new curve is :
    --          
    --           Poles.Length() + (NewDegree - Degree) * Number of spans
    --           
    --          Where the number of spans is :
    --          
    --           LastUKnotIndex(Mults) - FirstUKnotIndex(Mults) + 1
    --           
    --           for a non-periodic curve
    --           
    --           And Knots.Length() - 1 for a periodic curve.
    --          
    --          The multiplicities of all  knots  are increased by
    --          the degree elevation.
    --           
    --          The new knots are usually  the same knots with the
    --          exception of  a non-periodic curve with  the first
    --          and last multiplicity not  equal to Degree+1 where
    --          knots are removed  form the start  and the  bottom
    --          untils the sum of the  multiplicities is  equal to
    --          NewDegree+1  at the  knots   corresponding  to the
    --          first and last parameters of the curve.
    --          
    --          Example  :  Suppose a  curve  of degree 3 starting
    --          with following knots and multiplicities :
    --          
    --          knot : 0.  1.  2.
    --          mult : 1   2   1
    --          
    --          The  FirstUKnot is  2.     because the   sum    of
    --          multiplicities is Degree+1 : 1 + 2 + 1 = 4 = 3 + 1
    --          
    --          i.e. the first parameter  of the  curve is  2. and
    --          will still be   2.  after degree  elevation.   Let
    --          raises this curve to degree 4.  The multiplicities
    --          are increased by 2.
    --          
    --          They   become 2 3  2.   But     we need a   sum of
    --          multiplicities  of 5 at knot  2. So the first knot
    --          is removed and the new knots are :
    --          
    --          knot : 1.  2.
    --          mult : 3   2
    --          
    --          The multipicity   of the first  knot may   also be
    --          reduced if the sum is still to big.
    --          
    --          In the  most common situations (periodic  curve or
    --          curve with first and last multiplicities equals to
    --          Degree+1) the knots are knot changes.
    --          
    --          The method IncreaseDegreeCountKnots can be used to
    --          compute the new number of knots.\
    --
    ---Warning: To be used for Beziercurves ONLY!!!

    PrepareUnperiodize (Degree  : in  Integer         from Standard;
    	    	        Mults   : in  Array1OfInteger from TColStd;
    	    	        NbKnots : out Integer         from Standard; 
		        NbPoles : out Integer         from Standard);
    ---Purpose: Set in <NbKnots> and <NbPolesToAdd> the number of Knots and
    --          Poles   of  the NotPeriodic  Curve   identical  at the
    --          periodic     curve with    a  degree    <Degree>  ,  a
    --          knots-distribution with Multiplicities <Mults>.

    Unperiodize (Degree    : in  Integer         from Standard;
                 Dimension : in  Integer         from Standard;
    	         Mults     : in  Array1OfInteger from TColStd;
	         Knots     : in  Array1OfReal    from TColStd;
    	         Poles     : in  Array1OfReal    from TColStd;
    	         NewMults  : out Array1OfInteger from TColStd;
	         NewKnots  : out Array1OfReal    from TColStd;
	         NewPoles  : out Array1OfReal    from TColStd);
	       
    Unperiodize (Degree    : in  Integer         from Standard;
    	         Mults     : in  Array1OfInteger from TColStd;
	         Knots     : in  Array1OfReal    from TColStd;
    	         Poles     : in  Array1OfPnt     from TColgp;
	         Weights   : in  Array1OfReal    from TColStd;
    	         NewMults  : out Array1OfInteger from TColStd;
	         NewKnots  : out Array1OfReal    from TColStd;
	         NewPoles  : out Array1OfPnt     from TColgp;
                 NewWeights: out Array1OfReal    from TColStd);
	       
    Unperiodize (Degree    : in  Integer         from Standard;
    	         Mults     : in  Array1OfInteger from TColStd;
	         Knots     : in  Array1OfReal    from TColStd;
    	         Poles     : in  Array1OfPnt2d   from TColgp;
	         Weights   : in  Array1OfReal    from TColStd;
    	         NewMults  : out Array1OfInteger from TColStd;
	         NewKnots  : out Array1OfReal    from TColStd;
	         NewPoles  : out Array1OfPnt2d   from TColgp;
                 NewWeights: out Array1OfReal    from TColStd);
	       

    PrepareTrimming (Degree  : in  Integer         from Standard;
    	    	     Periodic: in  Boolean         from Standard;
    	    	     Knots   : in  Array1OfReal    from TColStd;
    	    	     Mults   : in  Array1OfInteger from TColStd;
		     U1      : in  Real            from Standard;
		     U2      : in  Real            from Standard;
    	    	     NbKnots : out Integer         from Standard; 
		     NbPoles : out Integer         from Standard);
    ---Purpose: Set in <NbKnots> and <NbPoles> the number of Knots and
    --          Poles of the  curve resulting  of  the trimming of the
    --          BSplinecurve definded with <degree>, <knots>, <mults>

    Trimming (Degree     : in  Integer         from Standard;
    	      Periodic   : in  Boolean         from Standard;
    	      Dimension  : in  Integer         from Standard;
              Knots      : in  Array1OfReal    from TColStd;
    	      Mults      : in  Array1OfInteger from TColStd;
	      Poles      : in  Array1OfReal    from TColStd;
	      U1         : in  Real            from Standard;
	      U2         : in  Real            from Standard;
	      NewKnots   : out Array1OfReal    from TColStd;
    	      NewMults   : out Array1OfInteger from TColStd;
	      NewPoles   : out Array1OfReal    from TColStd);


    Trimming (Degree     : in  Integer         from Standard;
    	      Periodic   : in  Boolean         from Standard;
              Knots      : in  Array1OfReal    from TColStd;
    	      Mults      : in  Array1OfInteger from TColStd;
	      Poles      : in  Array1OfPnt     from TColgp;
	      Weights    : in  Array1OfReal    from TColStd;
	      U1         : in  Real            from Standard;
	      U2         : in  Real            from Standard;
	      NewKnots   : out Array1OfReal    from TColStd;
    	      NewMults   : out Array1OfInteger from TColStd;
	      NewPoles   : out Array1OfPnt     from TColgp;
	      NewWeights : out Array1OfReal    from TColStd);


    Trimming (Degree     : in  Integer         from Standard;
    	      Periodic   : in  Boolean         from Standard;
              Knots      : in  Array1OfReal    from TColStd;
    	      Mults      : in  Array1OfInteger from TColStd;
	      Poles      : in  Array1OfPnt2d   from TColgp;
	      Weights    : in  Array1OfReal    from TColStd;
	      U1         : in  Real            from Standard;
	      U2         : in  Real            from Standard;
	      NewKnots   : out Array1OfReal    from TColStd;
    	      NewMults   : out Array1OfInteger from TColStd;
	      NewPoles   : out Array1OfPnt2d   from TColgp;
	      NewWeights : out Array1OfReal    from TColStd);





    -------------------------------------------------------------
    -------------------------------------------------------------
    ----------					   ----------
    ----------	    Curve Evaluations		   ----------
    ----------					   ----------
    -------------------------------------------------------------
    -------------------------------------------------------------
    
    D0(U        : in Real;
       Index    : in Integer; 
       Degree   : in Integer; 
       Periodic : in Boolean;
       Poles    : in Array1OfReal    from TColStd;
       Weights  : in Array1OfReal    from TColStd;
       Knots    : in Array1OfReal    from TColStd;
       Mults    : in Array1OfInteger from TColStd;
       P        : out Real);
     
    D0(U        : in Real;
       Index    : in Integer; 
       Degree   : in Integer; 
       Periodic : in Boolean;
       Poles    : in Array1OfPnt     from TColgp; 
       Weights  : in Array1OfReal    from TColStd;
       Knots    : in Array1OfReal    from TColStd;
       Mults    : in Array1OfInteger from TColStd;
       P        : out Pnt from gp);
     
    D0(U        : in Real;
       UIndex   : in Integer; 
       Degree   : in Integer; 
       Periodic : in Boolean;
       Poles    : in Array1OfPnt2d   from TColgp; 
       Weights  : in Array1OfReal    from TColStd;
       Knots    : in Array1OfReal    from TColStd;
       Mults    : in Array1OfInteger from TColStd;
       P        : out Pnt2d from gp);
     
    D0(U        : in Real;
       Poles    : in Array1OfPnt     from TColgp; 
       Weights  : in Array1OfReal    from TColStd;
       P        : out Pnt from gp);
    ---Warning: To be used for Beziercurves ONLY!!!

    D0(U        : in Real;
       Poles    : in Array1OfPnt2d   from TColgp; 
       Weights  : in Array1OfReal    from TColStd;
       P        : out Pnt2d from gp);
    ---Warning: To be used for Beziercurves ONLY!!!
     
    D1(U        : in Real;
       Index    : in Integer; 
       Degree   : in Integer; 
       Periodic : in Boolean;
       Poles    : in Array1OfReal    from TColStd; 
       Weights  : in Array1OfReal    from TColStd;
       Knots    : in Array1OfReal    from TColStd;
       Mults    : in Array1OfInteger from TColStd;
       P        : out Real;
       V        : out Real);
       
    D1(U        : in Real;
       Index    : in Integer; 
       Degree   : in Integer; 
       Periodic : in Boolean;
       Poles    : in Array1OfPnt     from TColgp; 
       Weights  : in Array1OfReal    from TColStd;
       Knots    : in Array1OfReal    from TColStd;
       Mults    : in Array1OfInteger from TColStd;
       P        : out Pnt from gp;
       V        : out Vec from gp);
       
    D1(U        : in Real;
       UIndex   : in Integer; 
       Degree   : in Integer; 
       Periodic : in Boolean;
       Poles    : in Array1OfPnt2d   from TColgp; 
       Weights  : in Array1OfReal    from TColStd;
       Knots    : in Array1OfReal    from TColStd;
       Mults    : in Array1OfInteger from TColStd;
       P        : out Pnt2d from gp;
       V        : out Vec2d from gp);
     
    D1(U        : in Real;
       Poles    : in Array1OfPnt     from TColgp; 
       Weights  : in Array1OfReal    from TColStd;
       P        : out Pnt from gp;
       V        : out Vec from gp);
    ---Warning: To be used for Beziercurves ONLY!!!

    D1(U        : in Real;
       Poles    : in Array1OfPnt2d   from TColgp; 
       Weights  : in Array1OfReal    from TColStd;
       P        : out Pnt2d from gp;
       V        : out Vec2d from gp);
    ---Warning: To be used for Beziercurves ONLY!!!

    D2(U        : in Real;
       Index    : in Integer; 
       Degree   : in Integer; 
       Periodic : in Boolean;
       Poles    : in Array1OfReal    from TColStd; 
       Weights  : in Array1OfReal    from TColStd;
       Knots    : in Array1OfReal    from TColStd;
       Mults    : in Array1OfInteger from TColStd;
       P        : out Real;
       V1,V2    : out Real);
     
    D2(U        : in Real;
       Index    : in Integer; 
       Degree   : in Integer; 
       Periodic : in Boolean;
       Poles    : in Array1OfPnt     from TColgp; 
       Weights  : in Array1OfReal    from TColStd;
       Knots    : in Array1OfReal    from TColStd;
       Mults    : in Array1OfInteger from TColStd;
       P        : out Pnt from gp;
       V1,V2    : out Vec from gp);
     
    D2(U        : in Real;
       UIndex   : in Integer; 
       Degree   : in Integer; 
       Periodic : in Boolean;
       Poles    : in Array1OfPnt2d   from TColgp; 
       Weights  : in Array1OfReal    from TColStd;
       Knots    : in Array1OfReal    from TColStd;
       Mults    : in Array1OfInteger from TColStd;
       P        : out Pnt2d from gp;
       V1,V2    : out Vec2d from gp);
     
    D2(U        : in Real;
       Poles    : in Array1OfPnt     from TColgp; 
       Weights  : in Array1OfReal    from TColStd;
       P        : out Pnt from gp;
       V1,V2    : out Vec from gp);
    ---Warning: To be used for Beziercurves ONLY!!!

    D2(U        : in Real;
       Poles    : in Array1OfPnt2d   from TColgp; 
       Weights  : in Array1OfReal    from TColStd;
       P        : out Pnt2d from gp;
       V1,V2    : out Vec2d from gp);
    ---Warning: To be used for Beziercurves ONLY!!!

    D3(U        : in Real;
       Index    : in Integer; 
       Degree   : in Integer; 
       Periodic : in Boolean;
       Poles    : in Array1OfReal    from TColStd; 
       Weights  : in Array1OfReal    from TColStd;
       Knots    : in Array1OfReal    from TColStd;
       Mults    : in Array1OfInteger from TColStd;
       P        : out Real;
       V1,V2,V3 : out Real);
     
    D3(U        : in Real;
       Index    : in Integer; 
       Degree   : in Integer; 
       Periodic : in Boolean;
       Poles    : in Array1OfPnt     from TColgp; 
       Weights  : in Array1OfReal    from TColStd;
       Knots    : in Array1OfReal    from TColStd;
       Mults    : in Array1OfInteger from TColStd;
       P        : out Pnt from gp;
       V1,V2,V3 : out Vec from gp);
     
    D3(U        : in Real;
       UIndex   : in Integer; 
       Degree   : in Integer; 
       Periodic : in Boolean;
       Poles    : in Array1OfPnt2d   from TColgp; 
       Weights  : in Array1OfReal    from TColStd;
       Knots    : in Array1OfReal    from TColStd;
       Mults    : in Array1OfInteger from TColStd;
       P        : out Pnt2d from gp;
       V1,V2,V3 : out Vec2d from gp);
       
    D3(U        : in Real;
       Poles    : in Array1OfPnt     from TColgp; 
       Weights  : in Array1OfReal    from TColStd;
       P        : out Pnt from gp;
       V1,V2,V3 : out Vec from gp);
    ---Warning: To be used for Beziercurves ONLY!!!

    D3(U        : in Real;
       Poles    : in Array1OfPnt2d   from TColgp; 
       Weights  : in Array1OfReal    from TColStd;
       P        : out Pnt2d from gp;
       V1,V2,V3 : out Vec2d from gp);
    ---Warning: To be used for Beziercurves ONLY!!!

    DN(U        : in Real;
       N        : in Integer;
       Index    : in Integer; 
       Degree   : in Integer; 
       Periodic : in Boolean;
       Poles    : in Array1OfReal    from TColStd; 
       Weights  : in Array1OfReal    from TColStd;
       Knots    : in Array1OfReal    from TColStd;
       Mults    : in Array1OfInteger from TColStd;
       VN       : out Real);
     
    DN(U        : in Real;
       N        : in Integer;
       Index    : in Integer; 
       Degree   : in Integer; 
       Periodic : in Boolean;
       Poles    : in Array1OfPnt     from TColgp; 
       Weights  : in Array1OfReal    from TColStd;
       Knots    : in Array1OfReal    from TColStd;
       Mults    : in Array1OfInteger from TColStd;
       VN       : out Vec from gp);
     
    DN(U        : in Real;
       N        : in Integer;
       UIndex   : in Integer; 
       Degree   : in Integer; 
       Periodic : in Boolean;
       Poles    : in Array1OfPnt2d   from TColgp; 
       Weights  : in Array1OfReal    from TColStd;
       Knots    : in Array1OfReal    from TColStd;
       Mults    : in Array1OfInteger from TColStd;
       V        : out Vec2d from gp);
     
    DN(U        : in Real;
       N        : in Integer;
       Poles    : in Array1OfPnt     from TColgp; 
       Weights  : in Array1OfReal    from TColStd;
       P        : out Pnt from gp;
       VN       : out Vec from gp);
    ---Warning: To be used for Beziercurves ONLY!!!

    DN(U        : in Real;
       N        : in Integer;
       Poles    : in Array1OfPnt2d   from TColgp; 
       Weights  : in Array1OfReal    from TColStd;
       P        : out Pnt2d from gp;
       VN       : out Vec2d from gp);
    ---Purpose:  The  above  functions  compute   values and
    --         derivatives in the following situations :
    --         
    --         * 3D, 2D and 1D
    --         
    --         * Rational or not Rational. 
    --         
    --         * Knots  and multiplicities or "flat knots" without
    --         multiplicities.
    --         
    --         * The  <Index>  is   the the  localization  of  the
    --         parameter in the knot sequence.  If <Index> is  out
    --         of range the correct value will be searched.
    --         
    --         
    --         VERY IMPORTANT!!!
    --         USE  BSplCLib::NoWeights()  as Weights argument for non
    --         rational curves computations.
    ---Warning: To be used for Beziercurves ONLY!!!

    EvalBsplineBasis(Side                       : in Integer ;
     	    	     DerivativeOrder            : in Integer ;
		     Order                      : in Integer ;
		     FlatKnots                  : Array1OfReal from TColStd ;
    	    	     Parameter                  : in Real    ;
		     FirstNonZeroBsplineIndex   : in out Integer ;
		     BsplineBasis               : in out Matrix from math)

    returns Integer  ; 
    ---Purpose: This  evaluates  the Bspline  Basis  at  a
    --          given  parameter  Parameter   up   to  the
    --          requested   DerivativeOrder  and store the
    --          result  in the  array BsplineBasis  in the
    --          following   fashion  
    --          BSplineBasis(1,1)   =  
    --          value of first non vanishing 
    --          Bspline function which has Index FirstNonZeroBsplineIndex 
    --            BsplineBasis(1,2)   = 
    --            value of second non vanishing 
    --          Bspline   function which  has   Index
    --          FirstNonZeroBsplineIndex + 1
    --          BsplineBasis(1,n)   = 
    --            value of second non vanishing non vanishing
    --          Bspline   function which  has   Index
    --          FirstNonZeroBsplineIndex + n (n <= Order) 
    --          BSplineBasis(2,1)   =  
    --          value of derivative of first non vanishing 
    --          Bspline function which has Index FirstNonZeroBsplineIndex 
    --            BSplineBasis(N,1)   =  
    --          value of Nth derivative of first non vanishing 
    --          Bspline function which has Index FirstNonZeroBsplineIndex
    --          if N <= DerivativeOrder + 1

    BuildBSpMatrix(Parameters   : in Array1OfReal from TColStd;
    	    	   OrderArray   : in Array1OfInteger from TColStd;
    	    	   FlatKnots    : in Array1OfReal from TColStd;
    	   	   Degree       : in Integer;
		   Matrix       : in out Matrix from math;
		   UpperBandWidth : out Integer ;
		   LowerBandWidth : out Integer) returns Integer ;
    ---Purpose: This Builds   a fully  blown   Matrix of
    --            (ni)
    --          Bi    (tj)  
    --          
    --          with i  and j within 1..Order + NumPoles
    --          The  integer ni is   the ith slot of the
    --          array OrderArray, tj is the jth slot of
    --          the array Parameters
    
    FactorBandedMatrix(Matrix            : in out Matrix from math ;
    	    	       UpperBandWidth    : in Integer ;
		       LowerBandWidth    : in Integer ;
    	    	       PivotIndexProblem : out Integer) returns Integer ; 
    ---Purpose: this  factors  the Banded Matrix in
    --         the LU form with a Banded storage of 
    --         components of the L matrix 
    --         WARNING : do not use if the Matrix is
    --         totally positive (It is the case for
    --         Bspline matrices build as above with
    --         parameters being the Schoenberg points

    SolveBandedSystem (Matrix : in Matrix from math ;
		       UpperBandWidth    : in Integer ;
		       LowerBandWidth    : in Integer ;
		       ArrayDimension    : in Integer ;
		       Array             : in out Real)
    returns Integer ;
    ---Purpose: This solves  the system Matrix.X =  B
    --         with when Matrix is factored in LU form
    --         The  Array   is    an   seen   as    an
    --         Array[1..N][1..ArrayDimension] with N =
    --         the  rank  of the  matrix  Matrix.  The
    --         result is stored   in Array  when  each
    --         coordinate is  solved that is  B is the
    --         array whose values are 
    --         B[i] = Array[i][p] for each p in 1..ArrayDimension
		    
    SolveBandedSystem (Matrix : in Matrix from math ;
    	    	       UpperBandWidth    : in Integer ;
		       LowerBandWidth    : in Integer ;
		       Array             : in out Array1OfPnt2d from TColgp)  
    returns Integer ;
    ---Purpose: This solves  the system Matrix.X =  B
    --         with when Matrix is factored in LU form
    --         The  Array   has the length of  
    --         the  rank  of the  matrix  Matrix.  The
    --         result is stored   in Array  when  each
    --         coordinate is  solved that is  B is the
    --         array whose values are 
    --         B[i] = Array[i][p] for each p in 1..ArrayDimension

    SolveBandedSystem (Matrix : in Matrix from math ;
    	    	       UpperBandWidth    : in Integer ;
		       LowerBandWidth    : in Integer ;
		       Array             : in out Array1OfPnt   from TColgp)  
    returns Integer ;
    ---Purpose: This solves  the system Matrix.X =  B
    --         with when Matrix is factored in LU form
    --         The  Array   has the length of 
    --         the  rank  of the  matrix  Matrix.  The
    --         result is stored   in Array  when  each
    --         coordinate is  solved that is  B is the
    --         array whose values are 
    --         B[i] = Array[i][p] for each p in 1..ArrayDimension

    SolveBandedSystem (Matrix : in Matrix from math ;
		       UpperBandWidth    : in Integer ;
		       LowerBandWidth    : in Integer ;
		       HomogenousFlag    : in Boolean ;
		       ArrayDimension    : Integer ; 
		       Array             : in out Real ;
                       Weights           : in out Real ) 
    returns Integer ;

    SolveBandedSystem (Matrix : in Matrix from math ;
    	    	       UpperBandWidth    : in Integer ;
		       LowerBandWidth    : in Integer ;
		       HomogenousFlag    : in Boolean ;
		       Array             : in out Array1OfPnt2d from TColgp; 
                       Weights           : in out Array1OfReal from TColStd  ) 
    returns Integer ;
    ---Purpose: This solves the  system Matrix.X =  B
    --         with when Matrix is factored in LU form
    --         The    Array   is    an   seen  as   an
    --         Array[1..N][1..ArrayDimension] with N =
    --         the  rank  of  the  matrix Matrix.  The
    --         result is  stored   in Array when  each
    --         coordinate is  solved that is B  is the
    --         array  whose   values     are   B[i]  =
    --         Array[i][p]       for     each  p    in
    --         1..ArrayDimension. If  HomogeneousFlag ==
    --         0  the  Poles  are  multiplied by   the
    --         Weights   uppon   Entry   and      once
    --         interpolation   is    carried  over the
    --         result of the  poles are divided by the
    --         result of   the   interpolation of  the
    --         weights. Otherwise if HomogenousFlag == 1
    --         the Poles and Weigths are treated homogenously 
    --         that is that those are interpolated as they
    --         are and result is returned without division
    --         by the interpolated weigths.

    SolveBandedSystem (Matrix : in Matrix from math ;
    	    	       UpperBandWidth    : in Integer ;
		       LowerBandWidth    : in Integer ;
		       HomogeneousFlag   : in Boolean ;
		       Array             : in out Array1OfPnt   from TColgp; 
                       Weights           : in out Array1OfReal from TColStd )
    returns Integer ;
    ---Purpose: This solves  the system Matrix.X =  B
    --         with when Matrix is factored in LU form
    --         The  Array   is    an   seen   as    an
    --         Array[1..N][1..ArrayDimension] with N =
    --         the  rank  of the  matrix  Matrix.  The
    --         result is stored   in Array  when  each
    --         coordinate is  solved that is  B is the
    --         array whose values are 
    --         B[i] = Array[i][p] for each p in 1..ArrayDimension
    --         If  HomogeneousFlag ==
    --         0  the  Poles  are  multiplied by   the
    --         Weights   uppon   Entry   and      once
    --         interpolation   is    carried  over the
    --         result of the  poles are divided by the
    --         result of   the   interpolation of  the
    --         weights. Otherwise if HomogenousFlag == 1
    --         the Poles and Weigths are treated homogenously 
    --         that is that those are interpolated as they
    --         are and result is returned without division
    --         by the interpolated weigths.

    MergeBSplineKnots(Tolerance         : Real from Standard  ;
    	              StartValue        : Real from Standard  ;
		      EndValue          : Real from Standard  ;
		      Degree1           : Integer from Standard ;
		      Knots1            : Array1OfReal    from TColStd ;
		      Mults1            : Array1OfInteger from TColStd ;
		      Degree2           : Integer from Standard ;
		      Knots2            : Array1OfReal    from TColStd ;
		      Mults2            : Array1OfInteger from TColStd ;
		      NumPoles          : in out Integer ;
		      NewKnots          : in out HArray1OfReal    from TColStd ;
		      NewMults          : in out HArray1OfInteger from TColStd) ;
    ---Purpose:  Merges  two knot vector by   setting the starting and
    --          ending values to StartValue and EndValue 

    FunctionReparameterise(Function            : EvaluatorFunction from BSplCLib ;          
		     BSplineDegree       : Integer ;
		     BSplineFlatKnots    : Array1OfReal from TColStd ;
    	    	     PolesDimension      : Integer ;
		     Poles               : in out Real ;
		     
    	    	     FlatKnots           : Array1OfReal from TColStd ;
		     NewDegree           : Integer ;
		     NewPoles            : in out Real ;
    	             Status              : in out Integer) ;
    ---Purpose: This function will compose  a given Vectorial BSpline F(t)
     --          defined  by its  BSplineDegree and BSplineFlatKnotsl,
     --          its Poles  array which are coded as  an array of Real
     --          of  the  form  [1..NumPoles][1..PolesDimension] with  a
     --          function     a(t) which is   assumed to   satisfy the
     --          following: 
     --
     --       1. F(a(t))  is a polynomial BSpline
     --          that can be expressed  exactly as a BSpline of degree
     --          NewDegree on the knots FlatKnots 
     --
     --       2. a(t) defines a differentiable
     --          isomorphism between the range of FlatKnots to the range
     --          of BSplineFlatKnots which is the 
     --          same as the  range of F(t)  
     --
     --  Warning: it is
     --          the caller's responsability to insure that conditions
     --          1. and  2. above are  satisfied : no check whatsoever
     --          is made in this method 
     --
     -- Status will return 0 if OK else it will return the pivot index 
     --        of the matrix that was inverted to compute the multiplied
     --        BSpline : the method used is interpolation at Schoenenberg
     --        points of F(a(t)) 	     
     
    FunctionReparameterise(
    	    	     Function            : EvaluatorFunction from BSplCLib ;          
		     BSplineDegree       : Integer ;
		     BSplineFlatKnots    : Array1OfReal from TColStd ;
		     Poles               : Array1OfReal from TColStd ;
		     
    	    	     FlatKnots           : Array1OfReal from TColStd ;
		     NewDegree           : Integer ;
		     NewPoles            : in out Array1OfReal from TColStd ;
    	             Status              : in out Integer) ;
     ---Purpose: This function will compose  a given Vectorial BSpline F(t)
     --          defined  by its  BSplineDegree and BSplineFlatKnotsl,
     --          its Poles  array which are coded as  an array of Real
     --          of  the  form  [1..NumPoles][1..PolesDimension] with  a
     --          function     a(t) which is   assumed to   satisfy the
     --          following: 
     --
     --       1. F(a(t))  is a polynomial BSpline
     --          that can be expressed  exactly as a BSpline of degree
     --          NewDegree on the knots FlatKnots 
     --
     --       2. a(t) defines a differentiable
     --          isomorphism between the range of FlatKnots to the range
     --          of BSplineFlatKnots which is the 
     --          same as the  range of F(t)  
     --
     --  Warning: it is
     --          the caller's responsability to insure that conditions
     --          1. and  2. above are  satisfied : no check whatsoever
     --          is made in this method 
     --
     -- Status will return 0 if OK else it will return the pivot index 
     --        of the matrix that was inverted to compute the multiplied
     --        BSpline : the method used is interpolation at Schoenenberg
     --        points of F(a(t)) 
     
    FunctionReparameterise( Function            : EvaluatorFunction from BSplCLib ;          
		     BSplineDegree       : Integer ;
		     BSplineFlatKnots    : Array1OfReal from TColStd ;
		     Poles               : Array1OfPnt from TColgp ;
		     
    	    	     FlatKnots           : Array1OfReal from TColStd ;
		     NewDegree           : Integer ;
		     NewPoles            : in out Array1OfPnt from TColgp ;
    	             Status              : in out Integer) ;
     ---Purpose: this will compose  a given Vectorial BSpline F(t)
     --          defined  by its  BSplineDegree and BSplineFlatKnotsl,
     --          its Poles  array which are coded as  an array of Real
     --          of  the  form  [1..NumPoles][1..PolesDimension] with  a
     --          function     a(t) which is   assumed to   satisfy the
     --          following  : 1. F(a(t))  is a polynomial BSpline
     --          that can be expressed  exactly as a BSpline of degree
     --          NewDegree on the knots FlatKnots 
     --                       2. a(t) defines a differentiable
     --          isomorphism between the range of FlatKnots to the range
     --          of BSplineFlatKnots which is the 
     --          same as the  range of F(t)  
     --  Warning: it is
     --          the caller's responsability to insure that conditions
     --          1. and  2. above are  satisfied : no check whatsoever
     --          is made in this method 
     -- Status will return 0 if OK else it will return the pivot index 
     --        of the matrix that was inverted to compute the multiplied
     --        BSpline : the method used is interpolation at Schoenenberg
     --        points of F(a(t)) 	
 
     FunctionReparameterise(
                     Function            : EvaluatorFunction from BSplCLib ;          
		     BSplineDegree       : Integer ;
		     BSplineFlatKnots    : Array1OfReal from TColStd ;
		     Poles               : Array1OfPnt2d from TColgp ;
		     
    	    	     FlatKnots           : Array1OfReal from TColStd ;
		     NewDegree           : Integer ;
		     NewPoles            : in out Array1OfPnt2d from TColgp ;
    	             Status              : in out Integer) ;     
     ---Purpose: this will compose  a given Vectorial BSpline F(t)
     --          defined  by its  BSplineDegree and BSplineFlatKnotsl,
     --          its Poles  array which are coded as  an array of Real
     --          of  the  form  [1..NumPoles][1..PolesDimension] with  a
     --          function     a(t) which is   assumed to   satisfy the
     --          following  : 1. F(a(t))  is a polynomial BSpline
     --          that can be expressed  exactly as a BSpline of degree
     --          NewDegree on the knots FlatKnots 
     --                       2. a(t) defines a differentiable
     --          isomorphism between the range of FlatKnots to the range
     --          of BSplineFlatKnots which is the 
     --          same as the  range of F(t)  
     --  Warning: it is
     --          the caller's responsability to insure that conditions
     --          1. and  2. above are  satisfied : no check whatsoever
     --          is made in this method 
     -- Status will return 0 if OK else it will return the pivot index 
     --        of the matrix that was inverted to compute the multiplied
     --        BSpline : the method used is interpolation at Schoenenberg
     --        points of F(a(t)) 	     

    FunctionMultiply(Function            : EvaluatorFunction from BSplCLib ;          
		     BSplineDegree       : Integer ;
		     BSplineFlatKnots    : Array1OfReal from TColStd ;
    	    	     PolesDimension      : Integer ;
		     Poles               : in out Real ;
    	    	     FlatKnots           : Array1OfReal from TColStd ;
		     NewDegree           : Integer ;
		     NewPoles            : in out Real ;
    	             Status              : in out Integer) ;
     ---Purpose: this will  multiply a given Vectorial BSpline F(t)
     --          defined  by its  BSplineDegree and BSplineFlatKnotsl,
     --          its Poles  array which are coded as  an array of Real
     --          of  the  form  [1..NumPoles][1..PolesDimension] by  a
     --          function     a(t) which is   assumed to   satisfy the
     --          following  : 1. a(t)  * F(t)  is a polynomial BSpline
     --          that can be expressed  exactly as a BSpline of degree
     --          NewDegree on the knots FlatKnots 2. the range of a(t)
     --           is the same as the  range of F(t)  
     --  Warning: it is
     --          the caller's responsability to insure that conditions
     --          1. and  2. above are  satisfied : no check whatsoever
     --          is made in this method 
     -- Status will return 0 if OK else it will return the pivot index 
     --        of the matrix that was inverted to compute the multiplied
     --        BSpline : the method used is interpolation at Schoenenberg
     --        points of a(t)*F(t) 

    FunctionMultiply(Function            : EvaluatorFunction from BSplCLib ;          
		     BSplineDegree       : Integer ;
		     BSplineFlatKnots    : Array1OfReal from TColStd ;
		     Poles               : Array1OfReal from TColStd ;
    	    	     FlatKnots           : Array1OfReal from TColStd ;
		     NewDegree           : Integer ;
		     NewPoles            : in out Array1OfReal from TColStd ;
    	             Status              : in out Integer) ;
     ---Purpose: this will  multiply a given Vectorial BSpline F(t)
     --          defined  by its  BSplineDegree and BSplineFlatKnotsl,
     --          its Poles  array which are coded as  an array of Real
     --          of  the  form  [1..NumPoles][1..PolesDimension] by  a
     --          function     a(t) which is   assumed to   satisfy the
     --          following  : 1. a(t)  * F(t)  is a polynomial BSpline
     --          that can be expressed  exactly as a BSpline of degree
     --          NewDegree on the knots FlatKnots 2. the range of a(t)
     --           is the same as the  range of F(t)  
     --  Warning: it is
     --          the caller's responsability to insure that conditions
     --          1. and  2. above are  satisfied : no check whatsoever
     --          is made in this method 
     -- Status will return 0 if OK else it will return the pivot index 
     --        of the matrix that was inverted to compute the multiplied
     --        BSpline : the method used is interpolation at Schoenenberg
     --        points of a(t)*F(t) 

    FunctionMultiply(Function            : EvaluatorFunction from BSplCLib ;          
		     BSplineDegree       : Integer ;
		     BSplineFlatKnots    : Array1OfReal from TColStd ;
		     Poles               : Array1OfPnt2d from TColgp ;
    	    	     FlatKnots           : Array1OfReal from TColStd ;
		     NewDegree           : Integer ;
		     NewPoles            : in out Array1OfPnt2d from TColgp ;
    	             Status              : in out Integer) ;
     ---Purpose: this will  multiply a given Vectorial BSpline F(t)
     --          defined  by its  BSplineDegree and BSplineFlatKnotsl,
     --          its Poles  array which are coded as  an array of Real
     --          of  the  form  [1..NumPoles][1..PolesDimension] by  a
     --          function     a(t) which is   assumed to   satisfy the
     --          following  : 1. a(t)  * F(t)  is a polynomial BSpline
     --          that can be expressed  exactly as a BSpline of degree
     --          NewDegree on the knots FlatKnots 2. the range of a(t)
     --           is the same as the  range of F(t)  
     --  Warning: it is
     --          the caller's responsability to insure that conditions
     --          1. and  2. above are  satisfied : no check whatsoever
     --          is made in this method 
     -- Status will return 0 if OK else it will return the pivot index 
     --        of the matrix that was inverted to compute the multiplied
     --        BSpline : the method used is interpolation at Schoenenberg
     --        points of a(t)*F(t) 

    FunctionMultiply(Function            : EvaluatorFunction from BSplCLib ;          
		     BSplineDegree       : Integer ;
		     BSplineFlatKnots    : Array1OfReal from TColStd ;
		     Poles               : Array1OfPnt from TColgp ;
    	    	     FlatKnots           : Array1OfReal from TColStd ;
		     NewDegree           : Integer ;
		     NewPoles            : in out Array1OfPnt from TColgp ;
    	             Status              : in out Integer) ;
     ---Purpose: this will  multiply a given Vectorial BSpline F(t)
     --          defined  by its  BSplineDegree and BSplineFlatKnotsl,
     --          its Poles  array which are coded as  an array of Real
     --          of  the  form  [1..NumPoles][1..PolesDimension] by  a
     --          function     a(t) which is   assumed to   satisfy the
     --          following  : 1. a(t)  * F(t)  is a polynomial BSpline
     --          that can be expressed  exactly as a BSpline of degree
     --          NewDegree on the knots FlatKnots 2. the range of a(t)
     --           is the same as the  range of F(t)  
     --  Warning: it is
     --          the caller's responsability to insure that conditions
     --          1. and  2. above are  satisfied : no check whatsoever
     --          is made in this method 
     -- Status will return 0 if OK else it will return the pivot index 
     --        of the matrix that was inverted to compute the multiplied
     --        BSpline : the method used is interpolation at Schoenenberg
     --        points of a(t)*F(t) 

    Eval(U                 : Real;
         PeriodicFlag      : Boolean ;
         DerivativeRequest : Integer ;
 	 ExtrapMode        : in out Integer ;
     	 Degree            : Integer;
         FlatKnots         : Array1OfReal from TColStd ;
	 ArrayDimension    : Integer ;
	 Poles             : in out Real ;
         Result            : in out Real) ; 
    ---Purpose: Perform the De Boor   algorithm  to  evaluate a point at
    --          parameter <U>, with <Degree> and <Dimension>.
    --          
    --          Poles is  an array of  Reals of size 
    --          
    --          <Dimension> *  <Degree>+1
    --          
    --          Containing the  poles.  At  the end <Poles> contains
    --          the current point.   Poles Contain all  the poles of
    --          the BsplineCurve, Knots  also Contains all the knots
    --          of the BsplineCurve.  ExtrapMode has two slots [0] =
    --          Degree used to extrapolate before the first knot [1]
    --          = Degre used to  extrapolate after the last knot has
    --          to be between 1 and  Degree

    Eval(U                 : Real;
         PeriodicFlag      : Boolean ;
         DerivativeRequest : Integer ;
	 ExtrapMode        : in out Integer ;
    	 Degree            : Integer;
         FlatKnots         : Array1OfReal from TColStd ;
	 ArrayDimension    : Integer ;
	 Poles             : in out Real ;
	 Weights           : in out Real ;
         PolesResult       : in out Real ;
         WeightsResult     : in out Real) ;
    ---Purpose: Perform the  De Boor algorithm  to evaluate a point at
    --          parameter   <U>,  with   <Degree>    and  <Dimension>.
    --          Evaluates by multiplying the  Poles by the Weights and
    --          gives  the homogeneous  result  in PolesResult that is
    --          the results of the evaluation of the numerator once it
    --          has     been  multiplied   by  the     weights and  in
    --          WeightsResult one has  the result of the evaluation of
    --          the denominator
    --          
    --  Warning:   <PolesResult> and <WeightsResult>  must be   dimensionned
    --          properly.

    Eval(U                 : Real;
         PeriodicFlag      : Boolean ;
	 HomogeneousFlag   : Boolean ;
	 ExtrapMode        : in out Integer ;
    	 Degree            : Integer;
         FlatKnots         : Array1OfReal from TColStd ;
	 Poles             : Array1OfPnt   from TColgp;
	 Weights           : Array1OfReal    from TColStd ;
         Point             : out Pnt from gp ;
         Weight            : in out Real) ;
    ---Purpose: Perform the evaluation of the Bspline Basis 
    --          and then multiplies by the weights
    --          this just evaluates the current point

    Eval(U                 : Real;
         PeriodicFlag      : Boolean ;
	 HomogeneousFlag   : Boolean ;
	 ExtrapMode        : in out Integer ;
    	 Degree            : Integer;
         FlatKnots         : Array1OfReal from TColStd ;
	 Poles             : Array1OfPnt2d   from TColgp;
	 Weights           : Array1OfReal    from TColStd ;
         Point             : out Pnt2d from gp ;
         Weight            : in out Real) ;
    ---Purpose: Perform the evaluation of the Bspline Basis 
    --          and then multiplies by the weights
    --          this just evaluates the current point
    --          

    TangExtendToConstraint(FlatKnots         : Array1OfReal from TColStd ;
	                   C1Coefficient     : Real ;
	                   NumPoles          : in Integer ;
	                   Poles             : in out Real ;
	                   Dimension         : Integer ;
	                   Degree            : Integer ;
	                   ConstraintPoint   : Array1OfReal from TColStd ;
	                   Continuity        : Integer ;
                           After             : Boolean ;
	                   NbPolesResult     : in out Integer ; 
			   NbKnotsRsult      : in out Integer ;
                           KnotsResult       : in out Real ;
                           PolesResult       : in out Real) ;
    ---Purpose: Extend a BSpline nD using the tangency map
    --          <C1Coefficient> is the coefficient of reparametrisation
    --          <Continuity> must be equal to 1, 2 or 3.
    --          <Degree> must be greater or equal than <Continuity> + 1.
    --          
    --  Warning:   <KnotsResult> and <PolesResult>  must be   dimensionned
    --          properly.

    CacheD0(U              : Real;
    	    Degree         : Integer;
            CacheParameter : Real;
	    SpanLenght     : Real;
	    Poles          : Array1OfPnt     from TColgp  ;
	    Weights        : Array1OfReal    from TColStd ;
            Point          : out Pnt from gp) ;
    ---Purpose: Perform the evaluation of the of the cache
    --          the parameter must be normalized between
    --          the 0 and 1 for the span.
    --          The Cache must be valid when calling this
    --          routine. Geom Package will insure that. 
    --          and then multiplies by the weights
    --          this just evaluates the current point
    --          the CacheParameter is where the Cache was
    --          constructed the SpanLength is to normalize
    --          the polynomial in the cache to avoid bad conditioning
    --          effects

    CacheD0(U              : Real;
    	    Degree          : Integer;
	    CacheParameter  : Real;
	    SpanLenght      : Real;
	    Poles           : Array1OfPnt2d   from TColgp;
	    Weights         : Array1OfReal    from TColStd ;
            Point           : out Pnt2d from gp) ;
    ---Purpose: Perform the evaluation of the Bspline Basis 
    --          and then multiplies by the weights
    --          this just evaluates the current point
    --          the parameter must be normalized between
    --          the 0 and 1 for the span.
    --          The Cache must be valid when calling this
    --          routine. Geom Package will insure that. 
    --          and then multiplies by the weights
    --          ththe CacheParameter is where the Cache was
    --          constructed the SpanLength is to normalize
    --          the polynomial in the cache to avoid bad conditioning
    --          effectsis just evaluates the current point
    
    CoefsD0(U             : Real;
	    Poles         : Array1OfPnt     from TColgp  ;
	    Weights       : Array1OfReal    from TColStd ;
            Point         : out Pnt from gp) ;
    ---Purpose: Calls CacheD0 for Bezier  Curves Arrays computed with
    --          the method PolesCoefficients. 
    --  Warning: To be used for Beziercurves ONLY!!!
    ---C++: inline
  
    CoefsD0(U             : Real;
	    Poles         : Array1OfPnt2d   from TColgp  ;
	    Weights       : Array1OfReal    from TColStd ;
            Point         : out Pnt2d from gp) ;
    ---Purpose: Calls CacheD0 for Bezier  Curves Arrays computed with
    --          the method PolesCoefficients. 
    --  Warning: To be used for Beziercurves ONLY!!!
    ---C++: inline
    
    CacheD1(U             : Real;
      	    Degree        : Integer;
            CacheParameter: Real;
	    SpanLenght    : Real;
  	    Poles         : Array1OfPnt     from TColgp  ;
	    Weights       : Array1OfReal    from TColStd ;
            Point         : out Pnt from gp ;
            Vec           : out Vec from gp) ;
    ---Purpose: Perform the evaluation of the of the cache
    --          the parameter must be normalized between
    --          the 0 and 1 for the span.
    --          The Cache must be valid when calling this
    --          routine. Geom Package will insure that. 
    --          and then multiplies by the weights
    --          this just evaluates the current point
    --          the CacheParameter is where the Cache was
    --          constructed the SpanLength is to normalize
    --          the polynomial in the cache to avoid bad conditioning
    --          effects

    CacheD1(U              : Real;
    	    Degree         : Integer;
	    CacheParameter : Real;
	    SpanLenght     : Real;
	    Poles          : Array1OfPnt2d   from TColgp;
	    Weights        : Array1OfReal    from TColStd ;
            Point          : out Pnt2d from gp ;
            Vec            : out Vec2d from gp) ;
    ---Purpose: Perform the evaluation of the Bspline Basis 
    --          and then multiplies by the weights
    --          this just evaluates the current point
    --          the parameter must be normalized between
    --          the 0 and 1 for the span.
    --          The Cache must be valid when calling this
    --          routine. Geom Package will insure that. 
    --          and then multiplies by the weights
    --          ththe CacheParameter is where the Cache was
    --          constructed the SpanLength is to normalize
    --          the polynomial in the cache to avoid bad conditioning
    --          effectsis just evaluates the current point

    CoefsD1(U             : Real;
	    Poles         : Array1OfPnt     from TColgp  ;
	    Weights       : Array1OfReal    from TColStd ;
            Point         : out Pnt from gp;
            Vec           : out Vec from gp) ;
    ---Purpose: Calls CacheD1 for Bezier  Curves Arrays computed with
    --          the method PolesCoefficients. 
    --  Warning: To be used for Beziercurves ONLY!!!
    ---C++: inline

    CoefsD1(U             : Real;
	    Poles         : Array1OfPnt2d     from TColgp  ;
	    Weights       : Array1OfReal    from TColStd ;
            Point         : out Pnt2d from gp;
            Vec           : out Vec2d from gp) ;
    ---Purpose: Calls CacheD1 for Bezier  Curves Arrays computed with
    --          the method PolesCoefficients. 
    --  Warning: To be used for Beziercurves ONLY!!!
    ---C++: inline

    CacheD2(U             : Real;
            Degree            : Integer;
            CacheParameter    : Real;
	    SpanLenght        : Real;
	    Poles             : Array1OfPnt     from TColgp  ;
	    Weights           : Array1OfReal    from TColStd ;
            Point             : out Pnt from gp ;
            Vec1,Vec2         : out Vec from gp) ;
    ---Purpose: Perform the evaluation of the of the cache
    --          the parameter must be normalized between
    --          the 0 and 1 for the span.
    --          The Cache must be valid when calling this
    --          routine. Geom Package will insure that. 
    --          and then multiplies by the weights
    --          this just evaluates the current point
    --          the CacheParameter is where the Cache was
    --          constructed the SpanLength is to normalize
    --          the polynomial in the cache to avoid bad conditioning
    --          effects

    CacheD2(U              : Real;
    	    Degree         : Integer;
	    CacheParameter : Real;
	    SpanLenght     : Real;
	    Poles          : Array1OfPnt2d   from TColgp;
	    Weights        : Array1OfReal    from TColStd ;
            Point          : out Pnt2d from gp ;
            Vec1,Vec2      : out Vec2d from gp) ;
    ---Purpose: Perform the evaluation of the Bspline Basis 
    --          and then multiplies by the weights
    --          this just evaluates the current point
    --          the parameter must be normalized between
    --          the 0 and 1 for the span.
    --          The Cache must be valid when calling this
    --          routine. Geom Package will insure that. 
    --          and then multiplies by the weights
    --          ththe CacheParameter is where the Cache was
    --          constructed the SpanLength is to normalize
    --          the polynomial in the cache to avoid bad conditioning
    --          effectsis just evaluates the current point

    CoefsD2(U             : Real;
	    Poles         : Array1OfPnt     from TColgp  ;
	    Weights       : Array1OfReal    from TColStd ;
            Point         : out Pnt from gp;
            Vec1,Vec2     : out Vec from gp) ;
    ---Purpose: Calls CacheD1 for Bezier  Curves Arrays computed with
    --          the method PolesCoefficients. 
    --  Warning: To be used for Beziercurves ONLY!!!
    ---C++: inline

    CoefsD2(U             : Real;
	    Poles         : Array1OfPnt2d     from TColgp  ;
	    Weights       : Array1OfReal    from TColStd ;
            Point         : out Pnt2d from gp;
            Vec1,Vec2     : out Vec2d from gp) ;
    ---Purpose: Calls CacheD1 for Bezier  Curves Arrays computed with
    --          the method PolesCoefficients. 
    --  Warning: To be used for Beziercurves ONLY!!!
    ---C++: inline


    CacheD3(U              : Real;
    	    Degree         : Integer;
            CacheParameter : Real;
	    SpanLenght     : Real;
	    Poles          : Array1OfPnt     from TColgp  ;
	    Weights        : Array1OfReal    from TColStd ;
            Point          : out Pnt from gp ;
            Vec1,Vec2,Vec3 : out Vec from gp) ;
    ---Purpose: Perform the evaluation of the of the cache
    --          the parameter must be normalized between
    --          the 0 and 1 for the span.
    --          The Cache must be valid when calling this
    --          routine. Geom Package will insure that. 
    --          and then multiplies by the weights
    --          this just evaluates the current point
    --          the CacheParameter is where the Cache was
    --          constructed the SpanLength is to normalize
    --          the polynomial in the cache to avoid bad conditioning
    --          effects

    CacheD3(U              : Real;
    	    Degree         : Integer;
	    CacheParameter : Real;
	    SpanLenght     : Real;
	    Poles          : Array1OfPnt2d   from TColgp;
	    Weights        : Array1OfReal    from TColStd ;
            Point          : out Pnt2d from gp ;
            Vec1,Vec2,Vec3 : out Vec2d from gp) ;
    ---Purpose: Perform the evaluation of the Bspline Basis 
    --          and then multiplies by the weights
    --          this just evaluates the current point
    --          the parameter must be normalized between
    --          the 0 and 1 for the span.
    --          The Cache must be valid when calling this
    --          routine. Geom Package will insure that. 
    --          and then multiplies by the weights
    --          ththe CacheParameter is where the Cache was
    --          constructed the SpanLength is to normalize
    --          the polynomial in the cache to avoid bad conditioning
    --          effectsis just evaluates the current point

    CoefsD3(U             : Real;
	    Poles         : Array1OfPnt     from TColgp  ;
	    Weights       : Array1OfReal    from TColStd ;
            Point         : out Pnt from gp;
            Vec1,Vec2,Vec3: out Vec from gp) ;
    ---Purpose: Calls CacheD1 for Bezier  Curves Arrays computed with
    --          the method PolesCoefficients. 
    --  Warning: To be used for Beziercurves ONLY!!!
    ---C++: inline

    CoefsD3(U             : Real;
	    Poles         : Array1OfPnt2d     from TColgp  ;
	    Weights       : Array1OfReal    from TColStd ;
            Point         : out Pnt2d from gp;
            Vec1,Vec2,Vec3: out Vec2d from gp) ;
    ---Purpose: Calls CacheD1 for Bezier  Curves Arrays computed with
    --          the method PolesCoefficients. 
    --  Warning: To be used for Beziercurves ONLY!!!
    ---C++: inline

    BuildCache(U                   : Real;
               InverseOfSpanDomain : Real;
               PeriodicFlag        : Boolean ;
	       Degree              : Integer;
               FlatKnots           : Array1OfReal  from TColStd ;
	       Poles               : Array1OfPnt   from TColgp;
	       Weights             : Array1OfReal    from TColStd ;
               CachePoles          : in out Array1OfPnt   from TColgp;
	       CacheWeights        : in out Array1OfReal    from TColStd)   ;
    ---Purpose: Perform the evaluation of the Taylor expansion
    --          of the Bspline normalized between 0 and 1.
    --          If rational computes the homogeneous Taylor expension
    --          for the numerator and stores it in CachePoles

    BuildCache(U                   : Real;
               InverseOfSpanDomain : Real;
               PeriodicFlag        : Boolean ;
	       Degree              : Integer;
               FlatKnots           : Array1OfReal    from TColStd ;
	       Poles               : Array1OfPnt2d   from TColgp;
	       Weights             : Array1OfReal    from TColStd ;
               CachePoles          : in out Array1OfPnt2d   from TColgp;
	       CacheWeights        : in out Array1OfReal    from TColStd)   ;
    ---Purpose: Perform the evaluation of the Taylor expansion
    --          of the Bspline normalized between 0 and 1.
    --          If rational computes the homogeneous Taylor expension
    --          for the numerator and stores it in CachePoles

    PolesCoefficients(Poles         : Array1OfPnt2d   from TColgp;
                      CachePoles    : in out Array1OfPnt2d   from TColgp);
    ---Warning: To be used for Beziercurves ONLY!!!
    ---C++: inline
	 
    PolesCoefficients(Poles         : Array1OfPnt2d   from TColgp;
	    	      Weights       : Array1OfReal    from TColStd ;
                      CachePoles    : in out Array1OfPnt2d   from TColgp;
	    	      CacheWeights  : in out Array1OfReal    from TColStd)   ;
    ---Warning: To be used for Beziercurves ONLY!!!
	 
    PolesCoefficients(Poles         : Array1OfPnt   from TColgp;
                      CachePoles    : in out Array1OfPnt   from TColgp);
    ---Warning: To be used for Beziercurves ONLY!!!
    ---C++: inline

    PolesCoefficients(Poles         : Array1OfPnt   from TColgp;
	    	      Weights       : Array1OfReal    from TColStd ;
                      CachePoles    : in out Array1OfPnt   from TColgp;
	    	      CacheWeights  : in out Array1OfReal    from TColStd)   ;
    ---Purpose: Encapsulation   of  BuildCache    to   perform   the
    --          evaluation  of the Taylor expansion for beziercurves
    --          at parameter 0.
    --  Warning: To be used for Beziercurves ONLY!!!

    FlatBezierKnots (Degree: Integer) returns Real;
    ---Purpose: Returns pointer to statically allocated array representing 
    --          flat knots for bezier curve of the specified degree.
    --          Raises OutOfRange if Degree > MaxDegree()
    ---C++: return const &

    BuildSchoenbergPoints(Degree    : Integer ;
			  FlatKnots :  Array1OfReal from TColStd ;
		          Parameters : in out Array1OfReal from TColStd)  ; 
    ---Purpose: builds the Schoenberg points from the flat knot
    --          used to interpolate a BSpline since the 
    --          BSpline matrix is invertible.
      
    Interpolate(Degree : Integer ;
    	        FlatKnots         : Array1OfReal    from TColStd ;
    	        Parameters        : Array1OfReal    from TColStd ;
	        ContactOrderArray : Array1OfInteger from TColStd ;
	        Poles             : in out  Array1OfPnt    from TColgp ;
	        InversionProblem  : out Integer) ;
    ---Purpose: Performs the interpolation of  the data given in
    --          the Poles  array  according  to the  requests in
    --          ContactOrderArray    that is      :           if
    --          ContactOrderArray(i) has value  d it means  that
    --          Poles(i)   containes the dth  derivative of  the
    --          function to be interpolated. The length L of the
    --          following arrays must be the same :
    --          Parameters, ContactOrderArray, Poles,
    --          The length of FlatKnots is Degree + L + 1
    --  Warning: 
    --          the method used to do that interpolation is 
    --          gauss elimination WITHOUT pivoting. Thus if the
    --          diagonal is not dominant there is no guarantee
    --          that the algorithm will work. Nevertheless for
    --          Cubic interpolation or interpolation at Scheonberg
    --          points the method will work
    --          The InversionProblem will report 0 if there was no
    --          problem else it will give the index of the faulty
    --          pivot

    Interpolate(Degree            : Integer ;
    	        FlatKnots         : Array1OfReal    from TColStd ;
    	        Parameters        : Array1OfReal    from TColStd ;
	        ContactOrderArray : Array1OfInteger from TColStd ;
	        Poles             : in out  Array1OfPnt2d    from TColgp ;
	        InversionProblem  : out Integer) ;
    ---Purpose: Performs the interpolation of  the data given in
    --          the Poles  array  according  to the  requests in
    --          ContactOrderArray    that is      :           if
    --          ContactOrderArray(i) has value  d it means  that
    --          Poles(i)   containes the dth  derivative of  the
    --          function to be interpolated. The length L of the
    --          following arrays must be the same :
    --          Parameters, ContactOrderArray, Poles,
    --          The length of FlatKnots is Degree + L + 1
    --  Warning: 
    --          the method used to do that interpolation is 
    --          gauss elimination WITHOUT pivoting. Thus if the
    --          diagonal is not dominant there is no guarantee
    --          that the algorithm will work. Nevertheless for
    --          Cubic interpolation at knots or interpolation at Scheonberg
    --          points the method will work.
    --          The InversionProblem w
    --          ll report 0 if there was no
    --          problem else it will give the index of the faulty
    --          pivot

    Interpolate(Degree : Integer ;
    	        FlatKnots         : Array1OfReal    from TColStd ;
    	        Parameters        : Array1OfReal    from TColStd ;
	        ContactOrderArray : Array1OfInteger from TColStd ;
	        Poles             : in out  Array1OfPnt    from TColgp   ; 
	        Weights           : in out  Array1OfReal    from TColStd  ;  
	        InversionProblem  : out Integer) ;
    ---Purpose: Performs the interpolation of  the data given in
    --          the Poles  array  according  to the  requests in
    --          ContactOrderArray    that is      :           if
    --          ContactOrderArray(i) has value  d it means  that
    --          Poles(i)   containes the dth  derivative of  the
    --          function to be interpolated. The length L of the
    --          following arrays must be the same :
    --          Parameters, ContactOrderArray, Poles,
    --          The length of FlatKnots is Degree + L + 1
    --  Warning: 
    --          the method used to do that interpolation is 
    --          gauss elimination WITHOUT pivoting. Thus if the
    --          diagonal is not dominant there is no guarantee
    --          that the algorithm will work. Nevertheless for
    --          Cubic interpolation at knots or interpolation at Scheonberg
    --          points the method will work.
    --          The InversionProblem will report 0 if there was no
    --          problem else it will give the index of the faulty
    --          pivot
    --          
    -- 

    Interpolate(Degree            : Integer ;
    	    	FlatKnots         : Array1OfReal    from TColStd ;
    	        Parameters        : Array1OfReal    from TColStd ;
	        ContactOrderArray : Array1OfInteger from TColStd ;
	        Poles             : in out  Array1OfPnt2d    from TColgp ; 
	        Weights           : in out  Array1OfReal from TColStd  ;
	        InversionProblem  : out Integer) ;
    ---Purpose: Performs the interpolation of  the data given in
    --          the Poles  array  according  to the  requests in
    --          ContactOrderArray    that is      :           if
    --          ContactOrderArray(i) has value  d it means  that
    --          Poles(i)   containes the dth  derivative of  the
    --          function to be interpolated. The length L of the
    --          following arrays must be the same :
    --          Parameters, ContactOrderArray, Poles,
    --          The length of FlatKnots is Degree + L + 1
    --  Warning: 
    --          the method used to do that interpolation is 
    --          gauss elimination WITHOUT pivoting. Thus if the
    --          diagonal is not dominant there is no guarantee
    --          that the algorithm will work. Nevertheless for
    --          Cubic interpolation at knots or interpolation at Scheonberg
    --          points the method will work.
    --          The InversionProblem w
    --          ll report 0 if there was no
    --          problem else it will give the i      

    Interpolate(Degree : Integer ;
    	        FlatKnots         : Array1OfReal    from TColStd ;
    	        Parameters        : Array1OfReal    from TColStd ;
	        ContactOrderArray : Array1OfInteger from TColStd ;
                ArrayDimension    : Integer ;
	        Poles             : in out Real  ;
	        InversionProblem  : out Integer) ;
    ---Purpose: Performs the interpolation of  the data given in
    --          the Poles  array  according  to the  requests in
    --          ContactOrderArray    that is      :           if
    --          ContactOrderArray(i) has value  d it means  that
    --          Poles(i)   containes the dth  derivative of  the
    --          function to be interpolated. The length L of the
    --          following arrays must be the same :
    --          Parameters, ContactOrderArray
    --          The length of FlatKnots is Degree + L + 1
    --          The  PolesArray   is    an   seen   as    an
    --          Array[1..N][1..ArrayDimension] with N = tge length
    --          of the parameters array
    --  Warning: 
    --          the method used to do that interpolation is 
    --          gauss elimination WITHOUT pivoting. Thus if the
    --          diagonal is not dominant there is no guarantee
    --          that the algorithm will work. Nevertheless for
    --          Cubic interpolation or interpolation at Scheonberg
    --          points the method will work
    --          The InversionProblem will report 0 if there was no
    --          problem else it will give the index of the faulty
    --          pivot
    --          

    Interpolate(Degree : Integer ;
    	        FlatKnots         : Array1OfReal    from TColStd ;
    	    	Parameters        : Array1OfReal    from TColStd ;
		ContactOrderArray : Array1OfInteger from TColStd ;
                ArrayDimension    : Integer ;
		Poles             : in out Real  ;
		Weights           : in out Real  ;
		InversionProblem  : out Integer) ;
		  
    MovePoint(U            : Real;          -- parameter of the point
              Displ        : Vec2d from gp; -- translation vector of the point
    	      Index1       : Integer;       -- first movable pole
	      Index2       : Integer;       -- last movable pole
              Degree       : Integer; 
              Rational     : Boolean;
              Poles        : Array1OfPnt2d   from TColgp;
              Weights      : Array1OfReal    from TColStd;
              FlatKnots    : Array1OfReal    from TColStd;
              FirstIndex   : in out Integer;       -- first pole modified
              LastIndex    : in out Integer;       -- last pole modified
              NewPoles     : in out Array1OfPnt2d  from TColgp); -- new poles
    ---Purpose: Find the new poles which allows  an old point (with a
    --          given  u as parameter) to reach a new position
    --          Index1 and Index2 indicate the range of poles we can move
    --          (1, NbPoles-1) or (2, NbPoles) -> no constraint for one side
    --                     don't enter (1,NbPoles) -> error: rigid move
    --          (2, NbPoles-1) -> the ends are enforced
    --          (3, NbPoles-2) -> the ends and the tangency are enforced
    --    if Problem in BSplineBasis calculation, no change for the curve
    --    and FirstIndex, LastIndex = 0

    MovePoint(U            : Real;          -- parameter of the point
              Displ        : Vec from gp;   -- translation vector of the point
    	      Index1       : Integer;       -- first movable pole
	      Index2       : Integer;       -- last movable pole
              Degree       : Integer; 
              Rational     : Boolean;
              Poles        : Array1OfPnt     from TColgp;
              Weights      : Array1OfReal    from TColStd;
              FlatKnots    : Array1OfReal    from TColStd;
              FirstIndex   : in out Integer;       -- first pole modified
              LastIndex   : in out Integer;       -- last pole modified
              NewPoles     : in out Array1OfPnt    from TColgp); -- new poles
    ---Purpose: Find the new poles which allows  an old point (with a
    --          given  u as parameter) to reach a new position
    --          Index1 and Index2 indicate the range of poles we can move
    --          (1, NbPoles-1) or (2, NbPoles) -> no constraint for one side
    --                     don't enter (1,NbPoles) -> error: rigid move
    --          (2, NbPoles-1) -> the ends are enforced
    --          (3, NbPoles-2) -> the ends and the tangency are enforced
    --    if Problem in BSplineBasis calculation, no change for the curve
    --    and FirstIndex, LastIndex = 0

    MovePointAndTangent(U                 : Real        ;
    	    	    	ArrayDimension    : Integer     ;
    	    	    	Delta             : in out Real ;  
			DeltaDerivative   : in out Real ;
                        Tolerance         : Real        ;
			Degree            : Integer     ; 
              	    	Rational          : Boolean     ;
			StartingCondition : Integer     ;
			EndingCondition   : Integer     ;
              	    	Poles        : in out Real      ;
              	    	Weights      : Array1OfReal           from TColStd;
              	    	FlatKnots    : Array1OfReal           from TColStd;
			NewPoles     : in out Real      ;
                        ErrorStatus  : in out Integer)  ;
    ---Purpose: This is the dimension free version of the utility
    -- U is the parameter  must be within the  first FlatKnots and the
    -- last FlatKnots  Delta is the amount the  curve has  to be moved
    -- DeltaDerivative is the  amount the derivative  has to be moved.
    -- Delta  and   DeltaDerivative   must be    array   of  dimension
    -- ArrayDimension  Degree  is the degree  of   the BSpline and the
    -- FlatKnots are the knots of the BSpline  Starting Condition if =
    -- -1 means the starting point of the curve can move 
    -- = 0 means the
    -- starting  point  of the cuve  cannot  move but  tangen  starting
    -- point of the curve cannot move
    -- = 1 means the starting point and tangents cannot move 
    -- = 2 means the starting point tangent and curvature cannot move
    -- = ...
    -- Same holds for EndingCondition
    -- Poles are the poles of the curve
    -- Weights are the weights of the curve if Rational = Standard_True
    -- NewPoles are the poles of the deformed curve 
    -- ErrorStatus will be 0 if no error happened
    --                     1 if there are not enough knots/poles
    --                          the imposed conditions
    -- The way to solve this problem is to add knots to the BSpline 
    -- If StartCondition = 1 and EndCondition = 1 then you need at least
    -- 4 + 2 = 6 poles so for example to have a C1 cubic you will need
    -- have at least 2 internal knots.

    MovePointAndTangent(U                 : Real        ;
    	    	    	Delta             : Vec from gp ;
			DeltaDerivative   : Vec from gp ;
                        Tolerance         : Real        ;
			Degree            : Integer     ; 
              	    	Rational          : Boolean     ;
			StartingCondition : Integer     ;
			EndingCondition   : Integer     ;
              	    	Poles        : Array1OfPnt  from TColgp           ;
              	    	Weights      : Array1OfReal           from TColStd;
              	    	FlatKnots    : Array1OfReal           from TColStd;
			NewPoles     : in out Array1OfPnt from TColgp      ;
                        ErrorStatus  : in out Integer)  ;
    ---Purpose: This is the dimension free version of the utility
    -- U is the parameter  must be within the  first FlatKnots and the
    -- last FlatKnots  Delta is the amount the  curve has  to be moved
    -- DeltaDerivative is the  amount the derivative  has to be moved.
    -- Delta  and   DeltaDerivative   must be    array   of  dimension
    -- ArrayDimension  Degree  is the degree  of   the BSpline and the
    -- FlatKnots are the knots of the BSpline  Starting Condition if =
    -- -1 means the starting point of the curve can move 
    -- = 0 means the
    -- starting  point  of the cuve  cannot  move but  tangen  starting
    -- point of the curve cannot move
    -- = 1 means the starting point and tangents cannot move 
    -- = 2 means the starting point tangent and curvature cannot move
    -- = ...
    -- Same holds for EndingCondition
    -- Poles are the poles of the curve
    -- Weights are the weights of the curve if Rational = Standard_True
    -- NewPoles are the poles of the deformed curve 
    -- ErrorStatus will be 0 if no error happened
    --                     1 if there are not enough knots/poles
    --                          the imposed conditions
    -- The way to solve this problem is to add knots to the BSpline 
    -- If StartCondition = 1 and EndCondition = 1 then you need at least
    -- 4 + 2 = 6 poles so for example to have a C1 cubic you will need
    -- have at least 2 internal knots.

    MovePointAndTangent(U                 : Real          ;
    	    	    	Delta             : Vec2d from gp ;
			DeltaDerivative   : Vec2d from gp ;
                        Tolerance         : Real          ;
			Degree            : Integer       ; 
              	    	Rational          : Boolean       ;
			StartingCondition : Integer       ;
			EndingCondition   : Integer       ;
              	    	Poles        : Array1OfPnt2d        from TColgp    ;
              	    	Weights      : Array1OfReal         from TColStd   ;
              	    	FlatKnots    : Array1OfReal         from TColStd   ;
			NewPoles     : in out Array1OfPnt2d from TColgp    ;
                        ErrorStatus  : in out Integer)  ;
    ---Purpose: This is the dimension free version of the utility
    -- U is the parameter  must be within the  first FlatKnots and the
    -- last FlatKnots  Delta is the amount the  curve has  to be moved
    -- DeltaDerivative is the  amount the derivative  has to be moved.
    -- Delta  and   DeltaDerivative   must be    array   of  dimension
    -- ArrayDimension  Degree  is the degree  of   the BSpline and the
    -- FlatKnots are the knots of the BSpline  Starting Condition if =
    -- -1 means the starting point of the curve can move 
    -- = 0 means the
    -- starting  point  of the cuve  cannot  move but  tangen  starting
    -- point of the curve cannot move
    -- = 1 means the starting point and tangents cannot move 
    -- = 2 means the starting point tangent and curvature cannot move
    -- = ...
    -- Same holds for EndingCondition
    -- Poles are the poles of the curve
    -- Weights are the weights of the curve if Rational = Standard_True
    -- NewPoles are the poles of the deformed curve 
    -- ErrorStatus will be 0 if no error happened
    --                     1 if there are not enough knots/poles
    --                          the imposed conditions
    -- The way to solve this problem is to add knots to the BSpline 
    -- If StartCondition = 1 and EndCondition = 1 then you need at least
    -- 4 + 2 = 6 poles so for example to have a C1 cubic you will need
    -- have at least 2 internal knots.

    Resolution(  PolesArray       : in out Real ;
    	         ArrayDimension   : Integer     ;
	         NumPoles         : Integer     ;
           	 Weights          : in Array1OfReal    from TColStd;
            	 FlatKnots        : in Array1OfReal    from TColStd;
            	 Degree           : in Integer;
    	    	 Tolerance3D      : Real     from Standard  ;
    	         UTolerance       : out Real from Standard) ;
    ---Purpose: 
    --          given a tolerance in 3D space returns a 
    --          tolerance    in U parameter space such that
    --          all u1 and u0 in the domain of the curve f(u) 
    --          | u1 - u0 | < UTolerance and 
    --          we have |f (u1) - f (u0)| < Tolerance3D

    Resolution(  Poles            : in Array1OfPnt  from TColgp  ;
           	 Weights          : in Array1OfReal from TColStd ;
		 NumPoles         : in Integer from Standard     ;
            	 FlatKnots        : in Array1OfReal from TColStd ;
            	 Degree           : in Integer from Standard     ;
    	    	 Tolerance3D      : Real     from Standard  ;
    	         UTolerance       : out Real from Standard) ;
    ---Purpose: 
    --          given a tolerance in 3D space returns a 
    --          tolerance    in U parameter space such that
    --          all u1 and u0 in the domain of the curve f(u) 
    --          | u1 - u0 | < UTolerance and 
    --          we have |f (u1) - f (u0)| < Tolerance3D

    Resolution(  Poles            : in Array1OfPnt2d from TColgp  ;
           	 Weights          : in Array1OfReal  from TColStd ;
                 NumPoles         : in Integer from Standard      ;
            	 FlatKnots        : in Array1OfReal  from TColStd ;
            	 Degree           : in Integer              ;
    	    	 Tolerance3D      : Real     from Standard  ;
    	         UTolerance       : out Real from Standard) ;
    ---Purpose: 
    --          given a tolerance in 3D space returns a 
    --          tolerance    in U parameter space such that
    --          all u1 and u0 in the domain of the curve f(u) 
    --          | u1 - u0 | < UTolerance and 
    --          we have |f (u1) - f (u0)| < Tolerance3D

end BSplCLib;

