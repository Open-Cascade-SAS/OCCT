-- Created on: 1994-10-03
-- Created by: Yves FRICAUD
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



package BRepMAT2d 

	---Purpose: 

uses
    MAT2d,
    MAT,
    TCollection,
    TColStd,
    TColGeom2d,
    Geom2d,
    gp,	
    TopoDS,
    TopTools
    
is
    class Explorer;
    	---Purpose: Construct an  explorer for  the computation of the 
    	--          bisecting locus  from a Wire, a  Face, or a set of 
    	--          curves from Geom2d.

    class BisectingLocus instantiates BisectingLocus from MAT2d 
    	    	    	    	    	  (Explorer  from BRepMAT2d);
	---Purpose: the map of bisecting locus.
					  
    class LinkTopoBilo;
    	---Purpose: Constucts links between the Wire or the Face and
    	--          the BasicElts contained in the bisecting locus.


    class SequenceOfBasicElt instantiates Sequence from TCollection
                                                         (BasicElt from MAT); 
							 
    class DataMapOfShapeSequenceOfBasicElt instantiates DataMap from TCollection 
    		    		    	      (Shape               from TopoDS, 
					       SequenceOfBasicElt  from  BRepMAT2d, 
					       ShapeMapHasher      from TopTools); 
    
    class DataMapOfBasicEltShape  instantiates
    	DataMap from TCollection (BasicElt            from MAT,
    	    	    	    	  Shape               from TopoDS,
    	    	    	    	  MapTransientHasher  from TColStd);				       

end BRepMAT2d;




