-- Created on: 1996-12-16
-- Created by: Bruno DUMORTIER
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package BiTgte 

	---Purpose: 

uses
    Adaptor3d,
    Bnd,
    GeomAbs,
    Geom2d,
    Geom,
    TopoDS,
    TopTools,
    BRepAlgo,
    BRepFill,
    BRepOffset,
    TCollection,
    TColStd,
    TColgp,
    gp

is
    enumeration ContactType is
    	FaceFace,
	FaceEdge,
	FaceVertex,
    	EdgeEdge,
	EdgeVertex,
	VertexVertex
    end ContactType;

    class Blend;

    private class CurveOnEdge;

    private class HCurveOnEdge instantiates 
    	GenHCurve from Adaptor3d(CurveOnEdge from BiTgte);

    private class CurveOnVertex;

    private class HCurveOnVertex instantiates 
    	GenHCurve from Adaptor3d(CurveOnVertex from BiTgte);

    private class DataMapOfShapeBox instantiates 
       	DataMap from TCollection(Shape          from TopoDS,
	    	    	    	 Box            from Bnd,
				 ShapeMapHasher from TopTools);

end BiTgte;
