-- Created on: 2002-12-10
-- Created by: data exchange team
-- Copyright (c) 2002-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V2.0

class CurveElementPurpose from StepElement
inherits SelectType from StepData

    ---Purpose: Representation of STEP SELECT type CurveElementPurpose

uses
    SelectMember from StepData,
    EnumeratedCurveElementPurpose from StepElement,
    HAsciiString from TCollection

is
    Create returns CurveElementPurpose from StepElement;
	---Purpose: Empty constructor

    CaseNum (me; ent: Transient) returns Integer;
	---Purpose: Recognizes a kind of CurveElementPurpose select type
	--          return 0 

    CaseMem (me; ent: SelectMember from StepData) returns Integer is redefined;
	---Purpose: Recognizes a items of select member CurveElementPurposeMember
	--          1 -> EnumeratedCurveElementPurpose
	--          2 -> ApplicationDefinedElementPurpose
	--          0 else


     NewMember(me) returns SelectMember from StepData is redefined;
	---Purpose: Returns a new select member the type CurveElementPurposeMember

    SetEnumeratedCurveElementPurpose(me: in out; aVal :EnumeratedCurveElementPurpose from StepElement);
	---Purpose: Set Value for EnumeratedCurveElementPurpose

    EnumeratedCurveElementPurpose (me) returns EnumeratedCurveElementPurpose from StepElement;
	---Purpose: Returns Value as EnumeratedCurveElementPurpose (or Null if another type)

    SetApplicationDefinedElementPurpose(me: in out; aVal :HAsciiString from TCollection);
	---Purpose: Set Value for ApplicationDefinedElementPurpose

    ApplicationDefinedElementPurpose (me) returns HAsciiString from TCollection;
	---Purpose: Returns Value as ApplicationDefinedElementPurpose (or Null if another type)

end CurveElementPurpose;
