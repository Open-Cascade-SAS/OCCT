-- Created on: 1997-02-12
-- Created by: Alexander BRIVIN
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class WWWAnchor from Vrml 

	---Purpose: defines a WWWAnchor node of VRML specifying group properties.
    	--  The  WWWAnchor  group  node  loads  a  new  scene  into  a  VRML  browser 
	--  when  one  of  its  children  is  closen.  Exactly  how  a  user  "chooses" 
	--  a  child  of  the  WWWAnchor  is  up  to  the  VRML browser. 
	--  WWWAnchor  with  an  empty  ("")  name  does  nothing  when  its   
	--  children  are  chosen. 
	--  WWWAnchor  behaves  like  a  Separator,  pushing  the  traversal  state 
	--  before  traversing  its  children  and  popping  it  afterwards.


uses
 
    AsciiString   from  TCollection,
    WWWAnchorMap  from  Vrml

is
    Create  (  aName         :  AsciiString   from  TCollection  =  "";
               aDescription  :  AsciiString   from  TCollection  =  "";
               aMap          :  WWWAnchorMap  from  Vrml  =  Vrml_MAP_NONE ) 
	 returns  WWWAnchor from Vrml;

    SetName ( me : in out;  aName : AsciiString   from  TCollection );
    Name ( me )  returns  AsciiString   from  TCollection;

    SetDescription ( me : in out;  aDescription : AsciiString   from  TCollection );
    Description ( me )  returns  AsciiString   from  TCollection;

    SetMap ( me : in out;  aMap :  WWWAnchorMap  from  Vrml );
    Map ( me )  returns  WWWAnchorMap  from  Vrml;

    Print  ( me;  anOStream: in out OStream from Standard) returns OStream from Standard;
    ---C++:  return  & 

fields
 
    myName         :  AsciiString     from  TCollection;	  -- URL name
    myDescription  :  AsciiString     from  TCollection;	  -- Useful description of scene
    myMap          :  WWWAnchorMap    from  Vrml;	          -- How to map pick to URL name

end WWWAnchor;

