-- Created on: 1993-10-14
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Cut from BRepAlgoAPI  
    inherits BooleanOperation from BRepAlgoAPI 
    
    ---Purpose:   
    -- The class Cut provides Boolean cut operation  
    -- between arguments and tools (Boolean Subtraction).

uses
    Shape from TopoDS,
    PaveFiller from BOPAlgo

is 
 
    Create 
        returns Cut from BRepAlgoAPI;   
    ---C++: alias "Standard_EXPORT virtual ~BRepAlgoAPI_Cut();"  
    --- Purpose: Empty constructor 
      
    Create (PF: PaveFiller from BOPAlgo)
        returns Cut from BRepAlgoAPI;  
    --- Purpose: Empty constructor        
    -- <PF> - PaveFiller object that is carried out 
     
    Create (S1,S2 : Shape from TopoDS)  
        returns Cut from BRepAlgoAPI;  
    ---Purpose: Constructor with two shapes  
    -- <S1>  -argument     
    -- <S2>  -tool 
    -- <anOperation> - the type of the operation
    -- Obsolete   

    Create (S1,S2 : Shape from TopoDS; 
            aDSF  : PaveFiller  from BOPAlgo; 
            bFWD  : Boolean from Standard=Standard_True)  
        returns Cut from BRepAlgoAPI;  
    ---Purpose: Constructor with two shapes  
    -- <S1>  -argument     
    -- <S2>  -tool  
    -- <anOperation> - the type of the operation 
    -- <PF> - PaveFiller object that is carried out  
    -- Obsolete    
     
end Cut;
