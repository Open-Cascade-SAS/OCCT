-- Created on: 2002-12-12
-- Created by: data exchange team
-- Copyright (c) 2002-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class Surface3dElementRepresentation from StepFEA
inherits ElementRepresentation from StepFEA

    ---Purpose: Representation of STEP entity Surface3dElementRepresentation

uses
    HAsciiString from TCollection,
    HArray1OfRepresentationItem from StepRepr,
    RepresentationContext from StepRepr,
    HArray1OfNodeRepresentation from StepFEA,
    FeaModel3d from StepFEA,
    Surface3dElementDescriptor from StepElement,
    SurfaceElementProperty from StepElement,
    ElementMaterial from StepElement

is
    Create returns Surface3dElementRepresentation from StepFEA;
	---Purpose: Empty constructor

    Init (me: mutable; aRepresentation_Name: HAsciiString from TCollection;
                       aRepresentation_Items: HArray1OfRepresentationItem from StepRepr;
                       aRepresentation_ContextOfItems: RepresentationContext from StepRepr;
                       aElementRepresentation_NodeList: HArray1OfNodeRepresentation from StepFEA;
                       aModelRef: FeaModel3d from StepFEA;
                       aElementDescriptor: Surface3dElementDescriptor from StepElement;
                       aProperty: SurfaceElementProperty from StepElement;
                       aMaterial: ElementMaterial from StepElement);
	---Purpose: Initialize all fields (own and inherited)

    ModelRef (me) returns FeaModel3d from StepFEA;
	---Purpose: Returns field ModelRef
    SetModelRef (me: mutable; ModelRef: FeaModel3d from StepFEA);
	---Purpose: Set field ModelRef

    ElementDescriptor (me) returns Surface3dElementDescriptor from StepElement;
	---Purpose: Returns field ElementDescriptor
    SetElementDescriptor (me: mutable; ElementDescriptor: Surface3dElementDescriptor from StepElement);
	---Purpose: Set field ElementDescriptor

    Property (me) returns SurfaceElementProperty from StepElement;
	---Purpose: Returns field Property
    SetProperty (me: mutable; Property: SurfaceElementProperty from StepElement);
	---Purpose: Set field Property

    Material (me) returns ElementMaterial from StepElement;
	---Purpose: Returns field Material
    SetMaterial (me: mutable; Material: ElementMaterial from StepElement);
	---Purpose: Set field Material

fields
    theModelRef: FeaModel3d from StepFEA;
    theElementDescriptor: Surface3dElementDescriptor from StepElement;
    theProperty: SurfaceElementProperty from StepElement;
    theMaterial: ElementMaterial from StepElement;

end Surface3dElementRepresentation;
