-- File:        AutoDesignPersonAndOrganizationAssignment.cdl
-- Created:     Mon Dec  4 12:02:23 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWAutoDesignPersonAndOrganizationAssignment from RWStepAP214

	---Purpose : Read & Write Module for AutoDesignPersonAndOrganizationAssignment

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     AutoDesignPersonAndOrganizationAssignment from StepAP214,
     EntityIterator from Interface

is

	Create returns RWAutoDesignPersonAndOrganizationAssignment;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable AutoDesignPersonAndOrganizationAssignment from StepAP214);

	WriteStep (me; SW : in out StepWriter; ent : AutoDesignPersonAndOrganizationAssignment from StepAP214);

	Share(me; ent : AutoDesignPersonAndOrganizationAssignment from StepAP214; iter : in out EntityIterator);

end RWAutoDesignPersonAndOrganizationAssignment;
