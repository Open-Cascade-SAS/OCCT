-- File:        Point.cdl
-- Created:     Mon Dec  4 12:02:29 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWPoint from RWStepGeom

	---Purpose : Read & Write Module for Point

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     Point from StepGeom

is

	Create returns RWPoint;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable Point from StepGeom);

	WriteStep (me; SW : in out StepWriter; ent : Point from StepGeom);

end RWPoint;
