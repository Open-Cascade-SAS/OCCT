-- Created on: 1993-03-02
-- Created by: Philippe DAUTRY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class ElementarySurface from PGeom inherits Surface from PGeom

        ---Purpose :  This class defines  the general behaviour of the
        --         following    elementary      surfaces    :   Plane,
        --         CylindricalSurface,                 ConicalSurface,
        --         SphericalSurface, ToroidalSurface.
        --  
        --  All these entities are located in 3D space with an axis
        --  placement (Location point, XAxis, YAxis, ZAxis). It is 
        --  their local coordinate system.
        --  
	---See Also : ElementarySurface from Geom.

uses Ax3     from gp

is


    Initialize;
	---Purpose: Initializes the field(s) with default value(s).
    	---Level: Internal 


    Initialize(aPosition : Ax3 from gp);
	---Purpose: Initializes the fields with these values.
    	---Level: Internal 


  Position (me: mutable; aPosition : Ax3 from gp);
       ---Purpose :  Set the field position with <aPosition>.
    	---Level: Internal 


  Position (me)  returns Ax3 from gp;
        --- Purpose : Returns the value of the field position.
    	---Level: Internal 


fields

  position               : Ax3     from gp      is protected;

end;
