-- Created on: 2002-12-12
-- Created by: data exchange team
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class ElementDescriptor from StepElement
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity ElementDescriptor

uses
    ElementOrder from StepElement,
    HAsciiString from TCollection

is
    Create returns ElementDescriptor from StepElement;
	---Purpose: Empty constructor

    Init (me: mutable; aTopologyOrder: ElementOrder from StepElement;
                       aDescription: HAsciiString from TCollection);
	---Purpose: Initialize all fields (own and inherited)

    TopologyOrder (me) returns ElementOrder from StepElement;
	---Purpose: Returns field TopologyOrder
    SetTopologyOrder (me: mutable; TopologyOrder: ElementOrder from StepElement);
	---Purpose: Set field TopologyOrder

    Description (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Description
    SetDescription (me: mutable; Description: HAsciiString from TCollection);
	---Purpose: Set field Description

fields
    theTopologyOrder: ElementOrder from StepElement;
    theDescription: HAsciiString from TCollection;

end ElementDescriptor;
