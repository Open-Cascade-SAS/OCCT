-- File:	MNaming_NanimgStorageDriver.cdl
-- Created:	Wed Sep 17 17:15:40 1997
-- Author:	Isabelle GRIGNON
--		<isg@bigbox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1997

class NamingStorageDriver from MNaming inherits ASDriver from MDF

	---Purpose: 

uses SRelocationTable from MDF,
     Attribute        from TDF,
     Attribute        from PDF, 
     MessageDriver    from CDM


is
   
    Create(theMessageDriver : MessageDriver from CDM) 
    returns mutable NamingStorageDriver from MNaming;

    VersionNumber(me) returns Integer from Standard;
	---Purpose: Returns the version number from which the driver
	--          is available: 0.

    SourceType(me) returns Type from Standard;
	---Purpose: Returns the type: Integer from TDataStd.

    NewEmpty (me) returns mutable Attribute from PDF;


    Paste(me;
    	  Source     :         Attribute from TDF;
    	  Target     : mutable Attribute from PDF;
    	  RelocTable : SRelocationTable from MDF);



end NamingStorageDriver;
