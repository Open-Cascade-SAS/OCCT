-- Created on: 1993-03-02
-- Created by: Philippe DAUTRY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SurfaceOfLinearExtrusion from PGeom inherits SweptSurface from PGeom

        ---Purpose : Generalised cylinder. This surface is obtained by
        --         sweeping a curve in a given direction.
        --         
	---See Also : SurfaceOfLinearExtrusion from Geom.

uses Dir         from gp,
     Curve       from PGeom,
     SurfaceForm from GeomAbs,
     Shape       from GeomAbs

is


  Create returns SurfaceOfLinearExtrusion from PGeom;
	---Purpose: Creates a SurfaceOfLinearExtrusion with default values.
    	---Level: Internal 


  Create (
    	    aBasisCurve : Curve from PGeom;
    	    aDirection  : Dir from gp)
     returns SurfaceOfLinearExtrusion from PGeom;
	---Purpose: Creates a SurfaceOfLinearExtrusion with these values.
    	---Level: Internal 


end;  
