-- Created on: 2008-04-10
-- Created by: Peter KURNEV <pkv@irinox>
-- Copyright (c) 2008-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


deferred class DiscretRoot from BRepMesh

inherits Transient from Standard

    ---Purpose:
    -- This is a common interface for meshing algorithms
    -- instantiated by Mesh Factory and implemented by plugins.

uses
    Shape from TopoDS

--raises

is
    Initialize
        returns DiscretRoot from BRepMesh;

    SetDeflection (           me : mutable;
                   theDeflection : Real from Standard);
    ---Purpose:
    -- Setup linear deflection.

    ---C++: alias "Standard_EXPORT virtual ~BRepMesh_DiscretRoot();"

    Deflection (me)
        returns Real from Standard;
    ---Purpose:
    -- Returns linear deflection.

    SetAngle (      me : mutable;
              theAngle : Real from Standard);
    ---Purpose:
    -- Setup angular deflection.

    Angle (me)
        returns Real from Standard;
    ---Purpose:
    -- Returns angular deflection.

    SetShape (      me : mutable;
              theShape : Shape from TopoDS);
    ---Purpose:
    -- Set the shape to triangulate.

    Shape (me)
        returns Shape from TopoDS;
    ---C++: return const &

    Perform (me : mutable)
        is deferred;
    ---Purpose:
    -- Compute triangulation for set shape.

    IsDone (me)
        returns Boolean from Standard;
    ---Purpose:
    -- Returns true if triangualtion was performed and has success.

    --
    --  Protected methods
    --
    SetDone (me : mutable)
        is protected;

    SetNotDone (me : mutable)
        is protected;

    Init (me : mutable)
        is virtual protected;

fields
    myDeflection : Real from Standard is protected;
    myAngle      : Real from Standard is protected;
    myShape      : Shape from TopoDS  is protected;
    myIsDone     : Boolean from Standard is protected;

end DiscretRoot;
