-- Created on: 1997-01-17
-- Created by: Philippe MANGIN
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class BSplineKnotSplitting from Law 

        --- Purpose :
        --  For a B-spline curve the discontinuities are localised at the
        --  knot values and between two knots values the B-spline is 
        --  infinitely continuously differentiable.
        --  At a knot of range index the continuity is equal to :
        --  Degree - Mult (Index)   where  Degree is the degree of the 
        --  basis B-spline functions and Mult the multiplicity of the knot
        --  of range Index.
        --  If for your computation you need to have B-spline curves with a 
        --  minima of continuity it can be interesting to know between which
        --  knot values, a B-spline curve arc, has a continuity of given order.
        --  This algorithm computes the indexes of the knots where you should
        --  split the curve, to obtain arcs with a constant continuity given
        --  at the construction time. The splitting values are in the range
        --  [FirstUKnotValue, LastUKnotValue] (See class B-spline curve from 
        --  package Geom).
        --  If you just want to compute the local derivatives on the curve you
        --  don't need to create the B-spline curve arcs, you can use the
        --  functions LocalD1, LocalD2, LocalD3, LocalDN of the class
        --  BSplineCurve.

        --- KeyWords : BSpline, Knot Splitting, Continuity
        --- See Also : File BSpline from package Law
        --- References : 
        --  Gerald Farin Curves and Surfaces for Computer Aided Geometric
        --  Design.


uses  Array1OfInteger      from TColStd,
      HArray1OfInteger     from TColStd,
      BSpline              from Law

raises DimensionError from Standard, 
       RangeError     from Standard
  
is

  Create (BasisLaw : BSpline from Law; ContinuityRange : Integer)
     returns BSplineKnotSplitting
        --- Purpose :
        --  Locates the knot values which correspond to the segmentation of
        --  the curve into arcs with a continuity equal to ContinuityRange.
     raises RangeError;
        --- Purpose : 
        --  Raised if ContinuityRange is not greater or equal zero.

  
  NbSplits (me)    returns Integer   is static;
        --- Purpose :
        --  Returns the number of knots corresponding to the splitting.


  Splitting (me; SplitValues : in out Array1OfInteger)
        --- Purpose : 
        --  Returns the indexes of the BSpline curve knots corresponding to 
        --  the splitting.
     raises DimensionError
        --- Purpose :
        --  Raised if the length of SplitValues is not equal to NbSPlit.
     is static;


  SplitValue (me; Index : Integer)   returns Integer 
        --- Purpose :
        --  Returns the index of the knot corresponding to the splitting
        --  of range Index.
     raises RangeError
        --- Purpose :
        --  Raised if Index < 1 or Index > NbSplits
     is static;
	      


fields  

  splitIndexes : HArray1OfInteger;

end BSplineKnotSplitting;
