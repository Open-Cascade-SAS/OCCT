-- Created on: 1992-09-28
-- Created by: Remi GILET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MakeLine from GCE2d inherits Root from GCE2d

    ---Purpose : This class implements the following algorithms used 
    --           to create a Line from Geom2d.
    --           * Create a Line parallel to another and passing 
    --             through a point.
    --           * Create a Line passing through 2 points.

uses Pnt2d from gp,
     Lin2d from gp,
     Ax2d  from gp,
     Dir2d from gp,
     Line  from Geom2d,
     Real  from Standard

raises NotDone from StdFail

is

Create (A : Ax2d from gp) returns MakeLine;
    --- Purpose :
    --  Creates a line located in 2D space with the axis placement A.
    --  The Location of A is the origin of the line. 

Create (L : Lin2d from gp) returns MakeLine;
    --- Purpose :
    --  Creates a line from a non persistent line from package gp.

Create (P : Pnt2d from gp; 
    	V : Dir2d from gp) returns MakeLine;
    --- Purpose :
    --  P is the origin and V is the direction of the line.

Create(Lin    :     Lin2d from gp;
       Point  :     Pnt2d from gp) returns MakeLine;
    ---Purpose : Make a Line from Geom2d <TheLin> parallel to another 
    --           Lin <Lin> and passing through a Pnt <Point>.

Create(Lin    :     Lin2d from gp      ;
       Dist   :     Real  from Standard) returns MakeLine;
    ---Purpose : Make a Line from Geom2d <TheLin> parallel to another 
    --           Lin <Lin> at a distance <Dist>.

Create(P1     :     Pnt2d from gp;
       P2     :     Pnt2d from gp) returns MakeLine;
    ---Purpose : Make a Line from Geom2d <TheLin> passing through 2 
    --           Pnt <P1>,<P2>.
    --           It returns false if <p1> and <P2> are confused.
    -- Warning
    -- If points P1 and P2 coincident (that is, when IsDone
    -- returns false), the Status function returns gce_ConfusedPoints.
        
Value(me) returns Line from Geom2d
    raises NotDone
    is static;
    ---C++: return const&
    ---Purpose: Returns the constructed line.
    -- Exceptions StdFail_NotDone if no line is constructed.
    ---C++: alias "operator const Handle(Geom2d_Line)& () const { return Value(); }"

fields

    TheLine : Line from Geom2d;
    --The solution from Geom2d.
    
end MakeLine;


