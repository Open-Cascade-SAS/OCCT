-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PersonOrganizationSelect from StepBasic inherits SelectType from StepData

	-- <PersonOrganizationSelect> is an EXPRESS Select Type construct translation.
	-- it gathers : Person, Organization, PersonAndOrganization

uses

	Person,
	Organization,
	PersonAndOrganization
is

	Create returns PersonOrganizationSelect;
	---Purpose : Returns a PersonOrganizationSelect SelectType

	CaseNum (me; ent : Transient) returns Integer;
	---Purpose: Recognizes a PersonOrganizationSelect Kind Entity that is :
	--        1 -> Person
	--        2 -> Organization
	--        3 -> PersonAndOrganization
	--        0 else

	Person (me) returns any Person;
	---Purpose : returns Value as a Person (Null if another type)

	Organization (me) returns any Organization;
	---Purpose : returns Value as a Organization (Null if another type)

	PersonAndOrganization (me) returns any PersonAndOrganization;
	---Purpose : returns Value as a PersonAndOrganization (Null if another type)


end PersonOrganizationSelect;

