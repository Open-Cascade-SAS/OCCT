-- File:        Torus.cdl
-- Created:     Mon Dec  4 12:02:32 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWTorus from RWStepShape

	---Purpose : Read & Write Module for Torus

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     Torus from StepShape,
     EntityIterator from Interface

is

	Create returns RWTorus;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable Torus from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : Torus from StepShape);

	Share(me; ent : Torus from StepShape; iter : in out EntityIterator);

end RWTorus;
