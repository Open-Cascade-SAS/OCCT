-- Created on: 2007-08-17
-- Created by: Sergey ZARITCHNY
-- Copyright (c) 2007-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class HDataMapOfStringByte from TDataStd inherits TShared from MMgt 

	---Purpose: Extension of TDataStd_DataMapOfStringByte class  
    	--          to be manipulated by handle.

uses
    DataMapOfStringByte from TDataStd 
    
is
    Create( NbBuckets: Integer from Standard = 1 )  
    returns mutable HDataMapOfStringByte from TDataStd;    
     
    Create( theOther:  DataMapOfStringByte from TDataStd)  
    returns mutable HDataMapOfStringByte from TDataStd;
     
    Map( me ) returns DataMapOfStringByte from TDataStd
	---C++: return const &
        ---C++: inline      
    is static;	    	
	  
    ChangeMap( me: mutable ) returns DataMapOfStringByte from TDataStd 
    	---C++: return &
        ---C++: inline 
    is static; 	    	
 
fields
    
    myMap : DataMapOfStringByte from TDataStd ;  
   
end HDataMapOfStringByte;
