-- Created by: NW,JPB,CAL
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

deferred class Window from Aspect

inherits
	TShared from MMgt

uses
        Background         from Aspect,
        GradientBackground from Aspect,
        TypeOfResize       from Aspect,
        FillMethod         from Aspect,
        GradientFillMethod from Aspect,
        Handle             from Aspect,
        Ratio              from Quantity,
        Parameter          from Quantity,
        NameOfColor        from Quantity,
        Color              from Quantity,
        AsciiString        from TCollection

raises
	WindowDefinitionError	from Aspect,
	WindowError	from Aspect

is
	Initialize;
	---Level: Public
	---Purpose: Initializes the datas of a Window.

	---------------------------------------------------
	-- Category: Methods to modify the class definition
	---------------------------------------------------

	SetBackground ( me	: mutable;
			ABack	: Background from Aspect );
	---Level: Public
	---Purpose: Modifies the window background.
	---Category: Methods to modify the class definition

    SetBackground ( me : mutable ;
                    theNameOfColor : NameOfColor from Quantity );
    ---Level: Public
    ---Purpose: Modifies the window background from a Named Color.
    ---Category: Methods to modify the class definition

    SetBackground ( me : mutable; color : Color from Quantity );
    ---Level: Public
    ---Purpose: Modifies the window background.
    ---Category: Methods to modify the class definition

    SetBackground( me: mutable;
		   ABackground: GradientBackground from Aspect);
    ---Level: Public
    ---Purpose: Modifies the window gradient background.
    ---Category: Methods to modify the class definition

    SetBackground( me: mutable;
		   theFirstColor:  Color from Quantity;
                   theSecondColor: Color from Quantity;
                   theFillMethod:  GradientFillMethod from Aspect);
    ---Level: Public
    ---Purpose: Modifies the window gradient background.
    ---Category: Methods to modify the class definition

	Map ( me )
		raises WindowError from Aspect is deferred;
	---Level: Public
	---Purpose: Opens the window <me>.
	---Category: Methods to modify the class definition

	Unmap ( me )
		raises WindowError from Aspect is deferred;
	---Level: Public
	---Purpose: Closes the window <me>.
	---Category: Methods to modify the class definition

	DoResize ( me ) returns TypeOfResize from Aspect
		raises WindowError from Aspect is deferred;
	---Level: Advanced
	---Purpose: Apply the resizing to the window <me>.
	---Category: Methods to modify the class definition

	DoMapping ( me ) returns Boolean from Standard
		raises WindowError from Aspect is deferred;
	---Level: Advanced
	---Purpose: Apply the mapping change to the window <me>.
	-- and returns TRUE if the window is mapped at screen.
	---Category: Methods to modify the class definition

        Destroy ( me : mutable )
		raises WindowError from Aspect is deferred;
	---Level: Advanced
        ---Purpose: Destroy the Window
        ---Category: Methods to modify the class definition

	----------------------------
	-- Category: Inquire methods
	----------------------------

	Background ( me ) returns Background from Aspect;
	---Level: Public
	---Purpose: Returns the window background.
	---Category: Inquire methods

	BackgroundFillMethod( me ) returns FillMethod from Aspect;
	---Level: Public
	---Purpose: Returns the current image background fill mode.

	GradientBackground ( me ) returns GradientBackground from Aspect;
	---Level: Public
	---Purpose: Returns the window gradient background.

	IsMapped ( me ) returns Boolean from Standard is deferred;
	---Level: Public
	---Purpose: Returns True if the window <me> is opened
	--	    and False if the window is closed.
	---Category: Inquire methods

        IsVirtual ( me ) returns Boolean from Standard;
        ---Level: Public
        ---Purpose: Returns True if the window <me> is virtual
        ---Category: Inquire methods

        SetVirtual ( me : mutable;
                     theVirtual : Boolean from Standard );
        ---Level: Public
        ---Purpose: Setup the virtual state
        ---Category: Inquire methods

        Ratio ( me ) returns Ratio from Quantity is deferred;
        ---Level: Public
        ---Purpose: Returns The Window RATIO equal to the physical
        --	    WIDTH/HEIGHT dimensions
        ---Category: Inquire methods

        Position ( me ;
                X1, Y1, X2, Y2 : out Integer from Standard )
        is deferred;
        ---Level: Public
        ---Purpose: Returns The Window POSITION in PIXEL
        ---Category: Inquire methods

        Size ( me ;
               Width, Height : out Integer from Standard )
        is deferred;
        ---Level: Public
        ---Purpose: Returns The Window SIZE in PIXEL
        ---Category: Inquire methods

fields
        MyBackground : Background from Aspect is protected;
        MyGradientBackground   : GradientBackground from Aspect is protected;
        MyBackgroundFillMethod : FillMethod from Aspect is protected;
        MyIsVirtual : Boolean from Standard is protected;
end Window;
