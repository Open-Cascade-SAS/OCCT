-- Created on: 1993-02-22
-- Created by: Philippe DAUTRY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class AxisPlacement from PGeom inherits Geometry from PGeom

        ---Purpose :   An  axis  placement  defines a  local cartesian
        --         coordinate  system and   can be used to  locate  an
        --         entity in 3D space.
        --  
	---See Also : AxisPlacement from Geom.

uses Ax1 from gp

is


    Initialize;
	---Purpose: Initializes the field(s) with default value(s).
    	---Level: Internal 


    Initialize(aAxis: Ax1 from gp);
	---Purpose: Initializes the field axis with <aAxis>.
    	---Level: Internal 


  Axis (me : mutable; aAxis : Ax1 from gp);
        --- Purpose : Set the field axis with <aAxis>.
    	---Level: Internal 


  Axis (me)  returns Ax1 from gp;
        --- Purpose : Returns the value of the field axis.
    	---Level: Internal 


fields

  axis : Ax1 from gp is protected;

end;
