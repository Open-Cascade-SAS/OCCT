-- Created on: 1994-01-19
-- Created by: CAL
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Modified:	GG RIC120302 add new constructor to pass Display structure
--		directly instead the connexion name.

class GraphicDevice from Graphic3d inherits GraphicDevice from Xw 

---Purpose: This class allows the definition of the Advanced
	--	    Graphic Device 
-- Warning: An Graphic Device is defined by a connexion
	--	    "host:server.screen" 


uses

	SharedLibrary	from OSD,
	GraphicDriver	from Aspect,
	Display		from Aspect,
	GraphicDriver	from Graphic3d,
	TypeOfMapping	from Xw,
	AsciiString     from TCollection

raises

	GraphicDeviceDefinitionError	from Aspect

is

	Create ( Connexion	: CString from Standard;
		 Mapping	: TypeOfMapping from Xw = Xw_TOM_COLORCUBE;
		 Ncolors	: Integer from Standard = 0;
		 UseDefault	: Boolean from Standard = Standard_True ) 
	returns mutable GraphicDevice from Graphic3d 
	---Level: Public
	---Purpose: Creates a GraphicDevice
	---Warning: Raises if the Device is badly defined
	raises GraphicDeviceDefinitionError from Aspect;

	Create ( DisplayHandle	: Display from Aspect)
	returns mutable GraphicDevice from Graphic3d 
	---Level: Public
	---Purpose: Creates a GraphicDevice from the Display structure
	---Warning: Raises if the Device is badly defined
	raises GraphicDeviceDefinitionError from Aspect;

	Destroy ( me	: mutable )
		is redefined static;
	---Level: Public
	---Purpose: Deletes the GraphicDevice <me>.
	---C++: alias ~

	GraphicDriver ( me )
		returns GraphicDriver from Aspect
		is redefined static;
	---Level: Public
	---Purpose: Returns the GraphicDriver.

	SetGraphicDriver ( me	: mutable )
		is private;
	---Level: Internal
	---Purpose: Sets the GraphicDriver.

	ShrEnvString ( me )
		returns AsciiString from TCollection
		is private;
	---Level: Internal
	---Purpose: Returns the environment string for loading shared graphics library.
	--	    The string can be defined in environment by corresponding variables,
	--      or default value will be used for loading from system library path
	--	    Environment variables : CSF_GraphicShr

fields

	MyGraphicDriver	:	GraphicDriver from Graphic3d;

end GraphicDevice from Graphic3d;
