-- Created on: 1993-07-16
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class LocationSet from TopTools 

	---Purpose: The class LocationSet stores a set of location in
	--          a relocatable state.
	--          
	--          It can be created from Locations.
	--          
	--          It can create Locations.
	--          
	--          It can be write and read from a stream.

uses
    Location             from TopLoc,
    IndexedMapOfLocation from TopLoc,
    ProgressIndicator    from Message

raises
    OutOfRange           from Standard

is
    Create returns LocationSet from TopTools;
	---Purpose: Returns an empty set of locations.
	
    Clear(me : in out)
	---Purpose: Clears the content of the set.
    is static;
	
    Add(me : in out; L : Location from TopLoc) returns Integer
	---Purpose: Incorporate a new Location in the  set and returns
	--          its index.
    is static;
    
    Location(me; I : Integer) returns Location from TopLoc
	---Purpose: Returns the location of index <I>.
	--          
	---C++: return const &
    raises
    	OutOfRange from Standard
    is static;

    Index(me; L : Location from TopLoc) returns Integer
	---Purpose: Returns the index of <L>.
    is static;
    
    Dump(me; OS : in out OStream)
	---Purpose: Dumps the content of me on the stream <OS>.
    is static;
	
    Write(me; OS : in out OStream)
	---Purpose: Writes the content of  me  on the stream <OS> in a
	--          format that can be read back by Read.
    is static;
	
    Read(me : in out; IS : in out IStream)
	---Purpose: Reads the content of me from the  stream  <IS>. me
	--          is first cleared.
	--          
    is static;
	
    SetProgress(me : in out; PR : ProgressIndicator from Message);

    GetProgress(me) returns ProgressIndicator from Message;

fields
    myMap : IndexedMapOfLocation from TopLoc;
    myProgress : ProgressIndicator from Message;

end LocationSet;


