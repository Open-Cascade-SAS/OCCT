-- Created on: 1995-10-19
-- Created by: Andre LIEUTIER
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PinpointConstraint from Plate
---Purpose : define a constraint on the Plate
--         

uses 
   XY from gp, 
   XYZ from gp

is
    Create returns PinpointConstraint;
    Create(point2d : XY ; ImposedValue : XYZ ;
           iu : Integer = 0; iv : Integer = 0) returns PinpointConstraint;

     -- Accessors :
    Pnt2d(me) returns XY from gp;
    ---C++: inline 
    ---C++: return const  &
    
    Idu(me) returns  Integer;
    ---C++: inline
    ---C++: return const &
    
    Idv(me) returns Integer;
    ---C++: inline
    ---C++: return const &
    
    Value(me) returns XYZ from gp;
    ---C++: inline
    ---C++: return const &
  
fields
    
    value : XYZ ;  
    pnt2d : XY ; 
    idu,idv : Integer;
   
end;
