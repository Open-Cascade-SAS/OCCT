-- Created by: NW,JPB,CAL
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class AspectMarker3d from Graphic3d inherits AspectMarker from Aspect

  ---Version:

  ---Purpose: Creates and updates an attribute group for
  --          marker type primitives. This group contains the type
  --          of marker, its colour, and its scale factor.
  ---Keywords: Marker, Color, Scale, Type

  ---Warning:
  ---References:

uses

  Color                 from Quantity,
  TypeOfMarker          from Aspect,
  HArray1OfByte         from TColStd,
  PixMap_Handle         from Image,
  MarkerImage_Handle    from Graphic3d,
  ShaderProgram_Handle  from Graphic3d

is

  Create
  returns AspectMarker3d from Graphic3d;
  ---Level: Public
  ---Purpose: Creates a context table for marker primitives
  --          defined with the following default values:
  --
  --          Marker type : TOM_X
  --          Colour      : YELLOW
  --          Scale factor: 1.0

  Create (theType             : TypeOfMarker from Aspect;
          theColor            : Color from Quantity;
          theScale            : Real from Standard)
  returns AspectMarker3d from Graphic3d;

  Create (theColor            : Color from Quantity;
          theWidth            : Integer from Standard;
          theHeight           : Integer from Standard;
          theTextureBitmap    : HArray1OfByte from TColStd)
  returns AspectMarker3d from Graphic3d;
  ---Level: Public
  ---Purpose: Creates a context table for marker primitives
  --          defined with the specified values.

  Create (theTextureImage     : PixMap_Handle from Image)
  returns AspectMarker3d from Graphic3d;
  ---Level: Public
  ---Purpose: Creates a context table for marker primitives
  --          defined with the specified values.

  GetTextureSize (me;
                  theWidth : out Integer from Standard;
                  theHeight: out Integer from Standard);
  ---Level: Public
  ---Purpose: Returns marker's texture size.

  GetMarkerImage (me)
  returns MarkerImage_Handle from Graphic3d;
  ---Level: Public
  ---Purpose: Returns marker's image texture.
  --- Could be null handle if marker aspect has been initialized as
  --- default type of marker.
  ---C++: return const &

  SetMarkerImage (me       : mutable;
                  theImage : MarkerImage_Handle from Graphic3d);
  ---Level: Public
  ---Purpose: Set marker's image texture.

  SetBitMap (me: mutable;
             theWidth  : Integer from Standard;
             theHeight : Integer from Standard;
             theTexture: HArray1OfByte from TColStd ) is static;

  SetShaderProgram ( me  :  mutable; 
                     theProgram  :  ShaderProgram_Handle from Graphic3d );
  ---Level: Public
  ---Purpose: Sets up OpenGL/GLSL shader program.

  ShaderProgram ( me )
  returns ShaderProgram_Handle from Graphic3d;
  ---C++: return const &

fields

--
-- Class: Graphic3d_AspectMarker3d
--
-- Purpose: Declaration of context-specific variables
--          for drawing 3d markers.
--
-- Reminder: A context for drawing 3d markers inherits:
--            - the colour
--            - the type of marker
--            - the scale factor
--           defined by AspectMarker.

myMarkerImage : MarkerImage_Handle from Graphic3d is protected;

MyShaderProgram  :  ShaderProgram_Handle  from  Graphic3d; 

end AspectMarker3d;
