-- Created by: Peter KURNEV
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.


class Context from IntTools  
    inherits TShared from MMgt


---Purpose:  
        --  The intersection Context contains geometrical  
        --  and topological toolkit (classifiers, projectors, etc). 
        --  The intersection Context is for caching the tools  
        --  to increase the performance.


uses  

    Pnt2d from gp,
    Pnt   from gp, 
    State from TopAbs,  
    Curve from Geom,   
    ProjectPointOnCurve from GeomAPI, 
    ProjectPointOnSurf  from GeomAPI,
    Vertex from TopoDS, 
    Face   from TopoDS,
    Edge   from TopoDS, 
    Solid  from TopoDS, 
    SolidClassifier from BRepClass3d, 
    FClass2d from IntTools,
    Curve    from IntTools, 
    BaseAllocator from BOPCol,
    DataMapOfShapeAddress from BOPCol, 
    DataMapOfTransientAddress from BOPCol, 
    Hatcher from Geom2dHatch, 
    SurfaceRangeLocalizeData from IntTools

--raises

is 
    Create   

    returns Context from IntTools;
    ---C++: alias "Standard_EXPORT virtual  ~IntTools_Context();"         
    Create (theAllocator: BaseAllocator from BOPCol) 

    returns Context from IntTools;
     
    FClass2d(me:mutable; 
        aF: Face from TopoDS) 
    returns FClass2d from IntTools; 
    ---C++: return & 
    ---Purpose:
    --- Returns a reference to point classifier
    --- for given face
    ---

    ProjPS (me:mutable; 
        aF: Face from TopoDS) 
    returns ProjectPointOnSurf from GeomAPI;
    ---C++: return &   
    ---Purpose:
    --- Returns a reference to point projector
    --- for given face
    ---

    ProjPC (me:mutable; 
        aE: Edge from TopoDS) 
    returns ProjectPointOnCurve from GeomAPI;
    ---C++: return &
    ---Purpose:
    --- Returns a reference to point projector
    --- for given edge
    ---

    ProjPT (me:mutable; 
        aC: Curve from Geom) 
    returns ProjectPointOnCurve from GeomAPI;
    ---C++: return &
    ---Purpose:
    --- Returns a reference to point projector
    --- for given curve
    ---

    SurfaceData(me: mutable; 
        aF: Face from TopoDS)
    returns SurfaceRangeLocalizeData from IntTools;
    ---C++: return &
    ---Purpose:
    --- Returns a reference to surface localization data
    --- for given face 
    
    SolidClassifier(me:mutable;  
        aSolid: Solid from TopoDS) 
    returns SolidClassifier from BRepClass3d; 
    ---C++: return &    
    ---Purpose:
    --- Returns a reference to solid classifier
    --- for given solid
    ---
 
    Hatcher(me: mutable;  
        aF: Face from TopoDS) 
    returns Hatcher from Geom2dHatch;
    ---C++: return &  
    ---Purpose:
    --- Returns a reference to 2D hatcher
    --- for given face
    --- 

    ComputePE  (me:mutable;  
       theP   : Pnt from gp; 
       theTolP: Real from Standard; 
       theE   : Edge   from  TopoDS; 
       theT   :out Real from Standard) 
    returns Integer from Standard;  
    ---Purpose:
    --- Computes parameter of the Point theP on
    --- the edge aE.
    --- Returns zero if the distance between point
    --- and edge is less than sum of tolerance value of edge and theTopP,
    --- otherwise and for following conditions returns
    --- negative value
    --- 1. the edge is degenerated (-1)
    --- 2. the edge does not contain 3d curve and pcurves (-2)
    --- 3. projection algorithm failed (-3)
    ---

    ComputeVE  (me:mutable;  
       aV   : Vertex from  TopoDS; 
       aE   : Edge   from  TopoDS; 
       aT   :out Real from Standard) 
    returns Integer from Standard;
    ---Purpose: 
    --- Computes parameter of the vertex aV on
    --- the edge aE.
    --- Returns zero if the distance between vertex
    --- and edge is less than sum of tolerances,
    --- otherwise and for following conditions returns
    --- negative value
    --- 1. the edge is degenerated (-1)
    --- 2. the edge does not contain 3d curve and pcurves (-2)
    --- 3. projection algorithm failed (-3)
    ---
         
    ComputeVF  (me:mutable;  
       aV  :     Vertex from  TopoDS; 
       aF  :     Face   from  TopoDS; 
       U   : out Real from Standard; 
       V   : out Real from Standard) 
    returns Integer from Standard;
    ---Purpose:
    --- Computes UV parameters of the vertex aV on face aF
    --- Returns zero if the distance between vertex and face is
    --- less than or equal the sum of tolerances and the projection 
    --- point lays inside boundaries of the face.
    --- For following conditions returns negative value
    --- 1. projection algorithm failed (-1)
    --- 2. distance is more than sum of tolerances (-2)
    --- 3. projection point out or on the boundaries of face (-3)
    --- 
    
    StatePointFace(me:mutable;    
       aF   :  Face   from  TopoDS;
       aP2D :  Pnt2d  from  gp) 
    returns State from TopAbs;  
    ---Purpose:
    --- Returns the state of the point aP2D
    --- relative to face aF
    ---
         
    IsPointInFace(me:mutable;    
       aF   :  Face   from  TopoDS;
       aP2D :  Pnt2d  from  gp) 
    returns Boolean from Standard; 
    ---Purpose:
    --- Returns true if the point aP2D is
    --- inside the boundaries of the face aF,
    --- otherwise returns false
    ---
 
    IsPointInFace(me:mutable;    
       aP3D :  Pnt   from  gp; 
       aF   :  Face  from TopoDS; 
       aTol :  Real from Standard) 
    returns Boolean from Standard; 
    ---Purpose:
    --- Returns true if the point aP2D is
    --- inside the boundaries of the face aF,
    --- otherwise returns false
    ---
    
    IsPointInOnFace(me:mutable;     
       aF   :  Face   from  TopoDS;
       aP2D :  Pnt2d  from  gp) 
    returns Boolean from Standard;
    ---Purpose:
    --- Returns true if the point aP2D is
    --- inside or on the boundaries of aF
    ---
         
    IsValidPointForFace(me:mutable;
       aP3D :  Pnt   from  gp; 
       aF   :  Face  from TopoDS; 
       aTol :  Real from Standard) 
    returns Boolean from Standard;
    ---Purpose:
    --- Returns true if the distance between point aP3D
    --- and face aF is less or equal to tolerance aTol
    --- and projection point is inside or on the boundaries
    --- of the face aF
    ---

    IsValidPointForFaces(me:mutable;
       aP3D :  Pnt   from  gp; 
       aF1  :  Face  from TopoDS; 
       aF2  :  Face  from TopoDS;
       aTol :  Real from Standard)   
    returns Boolean from Standard; 
    ---Purpose:
    --- Returns true if IsValidPointForFace returns true
    --- for both face aF1 and aF2
    ---
         
    IsValidBlockForFace (me:mutable;  
       aT1  :  Real  from Standard;      
       aT2  :  Real  from Standard;      
       aIC  :  Curve from IntTools; 
       aF   :  Face  from TopoDS; 
       aTol :  Real from Standard) 
    returns Boolean from Standard; 
    ---Purpose:
    --- Returns true if IsValidPointForFace returns true
    --- for some 3d point that lay on the curve aIC bounded by
    --- parameters aT1 and aT2
    ---

    IsValidBlockForFaces (me:mutable;  
       aT1  :  Real  from Standard;      
       aT2  :  Real  from Standard;      
       aIC  :  Curve from IntTools; 
       aF1  :  Face  from TopoDS; 
       aF2  :  Face  from TopoDS; 
       aTol :  Real from Standard) 
    returns Boolean from Standard;
    ---Purpose:
    --- Returns true if IsValidBlockForFace returns true
    --- for both faces aF1 and aF2
    ---
         
    IsVertexOnLine(me:mutable;  
       aV   :  Vertex from  TopoDS;  
       aIC  :  Curve from IntTools;  
       aTolC:  Real  from Standard; 
       aT   :out  Real  from Standard)   
    returns Boolean from Standard; 
    ---Purpose:
    --- Computes parameter of the vertex aV on
    --- the curve aIC.
    --- Returns true if the distance between vertex and
    --- curve is less than sum of tolerance of aV and aTolC,
    --- otherwise or if projection algorithm failed
    --- returns false (in this case aT isn't significant)
    --- 
        
    IsVertexOnLine(me:mutable;  
       aV   :  Vertex from  TopoDS; 
       aTolV:  Real  from Standard;  
       aIC  :  Curve from IntTools;  
       aTolC:  Real  from Standard; 
       aT   :out  Real  from Standard)   
    returns Boolean from Standard;
    ---Purpose:
    --- Computes parameter of the vertex aV on
    --- the curve aIC.
    --- Returns true if the distance between vertex and
    --- curve is less than sum of tolerance of aV and aTolC,
    --- otherwise or if projection algorithm failed
    --- returns false (in this case aT isn't significant)
    --- 

    ProjectPointOnEdge (me:mutable;  
       aP   : Pnt  from  gp;       
       aE   : Edge from  TopoDS;                    
       aT   :out Real from  Standard) 
    returns Boolean from Standard; 
    ---Purpose:
    --- Computes parameter of the point aP on
    --- the edge aE.
    --- Returns false if projection algorithm failed
    --- other wiese returns true.
    ---
     
fields 
    myAllocator  : BaseAllocator from BOPCol is protected;
    myFClass2dMap:DataMapOfShapeAddress from BOPCol is protected; 
    myProjPSMap  :DataMapOfShapeAddress from BOPCol is protected; 
    myProjPCMap  :DataMapOfShapeAddress from BOPCol is protected;    
    mySClassMap  :DataMapOfShapeAddress from BOPCol is protected;
    myProjPTMap  :DataMapOfTransientAddress from BOPCol is protected;    
    myHatcherMap :DataMapOfShapeAddress from BOPCol is protected; 
    myProjSDataMap:DataMapOfShapeAddress from BOPCol is protected; 
    myCreateFlag :Integer from Standard is protected; 
     
end Context;

