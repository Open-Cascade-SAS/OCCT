-- Created on: 1998-07-29
-- Created by: Administrateur Atelier XSTEP
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class EditSDR  from STEPEdit    inherits Editor  from IFSelect

    ---Purpose : EditSDR is an Editor fit for a Shape Definition Representation
    --           which designates a Product Definition

uses Transient, AsciiString, HAsciiString, InterfaceModel, EditForm

is

    Create returns EditSDR;

    Label (me) returns AsciiString;

    Recognize (me; form : EditForm) returns Boolean;

    StringValue (me; form : EditForm;  num : Integer)
    	returns HAsciiString from TCollection;

    Apply (me; form : EditForm; ent : Transient; model : InterfaceModel)
    	returns Boolean;

    Load (me; form : EditForm; ent : Transient; model : InterfaceModel)
    	returns Boolean;

end EditSDR;
