-- Created on: 1991-11-04
-- Created by: NW,JPB,CAL
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Edge from Aspect

	---Version:

	---Purpose: This class allows the definition of an edge.

	---Keywords: Edge, Visible, Invisible, Border, Line, Face

	---Warning:
	---References:

uses

	TypeOfEdge	from Aspect

raises

	EdgeDefinitionError	from Aspect

is

	Create
		returns Edge from Aspect;
	---Level: Public
	---Purpose: Creates an edge.

	Create ( AIndex1, AIndex2	: Integer from Standard;
		 AType			: TypeOfEdge from Aspect )
		returns Edge from Aspect
	---Level: Public
	---Purpose: Creates an edge from an index of vertices
	--	    in a table of vertices.
	--	    <AType> indicates if this edge is seen or not.
	--  Warning: Raises EdgeDefinitionError if AIndex1 == AIndex2.
	raises EdgeDefinitionError from Aspect;

	---------------------------------------------------
	-- Category: Methods to modify the class definition
	---------------------------------------------------

	SetValues ( me			: in out;
		    AIndex1, AIndex2	: Integer from Standard;
		    AType		: TypeOfEdge from Aspect )
	---Level: Public
	---Purpose: Updates the values of an edge <me>.
	--  Warning: Raises EdgeDefinitionError if AIndex1 == AIndex2.
	raises EdgeDefinitionError from Aspect;

	----------------------------
	-- Category: Inquire methods
	----------------------------

	Values ( me;
		 AIndex1, AIndex2	: out Integer from Standard;
		 AType			: out TypeOfEdge from Aspect );
	---Level: Public
	---Purpose: Returns the index of the vertices and the
	--	    type of edge <me>.
	---Category: Inquire methods

	FirstIndex ( me )
		returns Integer from Standard;
	---Level: Public
	---Purpose: Returns the index of the begin of the edge <me>.
	---Category: Inquire methods

	LastIndex ( me )
		returns Integer from Standard;
	---Level: Public
	---Purpose: Returns the index of the end of the edge <me>.
	---Category: Inquire methods

	Type ( me)
		returns TypeOfEdge from Aspect;
	---Level: Public
	---Purpose: Returns the type of the edge <me>.
	---Category: Inquire methods

--

fields

--
-- Class	:	Aspect_Edge
--
-- Purpose	:	Declaration of variables specific to edges
--
-- Reminder	:	An edge is defined by :
--			- two vertices referenced by indices
--			- its visibility
--

	-- indices of the vertices
	MyBegin		:	Integer from Standard;
	MyEnd		:	Integer from Standard;

	-- the visibility
	MyVisibility	:	TypeOfEdge from Aspect;

end Edge;
