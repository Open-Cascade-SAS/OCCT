-- Created on: 1993-05-04
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred generic class SITool from IntStart
    (ThePSurface as any)
                                   

	---Purpose: Template class for an additional tool on a bi-parametrised
	--          surface.


uses State from TopAbs

is

    NbSamplePoints(myclass; S: ThePSurface)

    	returns Integer from Standard;


    SamplePoint(myclass; S: ThePSurface; Index: Integer from Standard;
                U,V: out Real from Standard);


--    Classify(myclass; S: ThePSurface; U,V: Real from Standard)
--    
--    	returns State from TopAbs;


end SITool;
