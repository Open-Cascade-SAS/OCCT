-- Created on: 1997-02-11
-- Created by: Alexander BRIVIN and Dmitry TARASOV
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Normal from Vrml inherits  TShared  from  MMgt

	---Purpose: defines a Normal node of VRML specifying properties of geometry
	---          and its appearance.
    	--  This node defines a set of 3D surface normal vectors to be used by vertex-based shape
      	--  nodes (IndexedFaceSet, IndexedLineSet, PointSet) that follow it in the scene graph. This
      	--  node does not produce a visible result during rendering; it simply replaces the current
       	--  normals in the rendering state for subsequent nodes to use. This node contains one
       	--  multiple-valued field that contains the normal vectors. 
uses
 
  HArray1OfVec  from  TColgp 

is
 
    Create  (  aVector :  HArray1OfVec  from  TColgp  ) 
      returns  mutable Normal from Vrml;

    Create  returns  mutable  Normal  from  Vrml; 
    
    SetVector ( me  :  mutable;  aVector : HArray1OfVec  from  TColgp );
    Vector ( me )  returns  HArray1OfVec  from  TColgp;

    Print  ( me;  anOStream: in out OStream from Standard) returns OStream from Standard;
    ---C++:  return  & 

fields
 
    myVector  :  HArray1OfVec  from  TColgp;  -- Normal vector(s)

end Normal;
