-- Created on: 2000-09-07
-- Created by: TURIN  Anatoliy <ati@nnov.matra-dtv.fr>
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package StdLDrivers

uses  

    PDF,
    Standard,
    TCollection,
    CDM,
    PCDM,
    TDF,
    PDF,
    MDF,
    TDocStd,
    MDocStd,
    PDocStd
 
is 
    
    class DocumentRetrievalDriver;
    
    class DocumentStorageDriver;


    ---Category: Factory methods
    --           ==============================================================

    Factory (aGUID: GUID from Standard)
    returns Transient from Standard;
	---Purpose: Depending from the  ID, returns a list of  storage
	--          or retrieval attribute drivers. Used for plugin
		   
end PAppStdL;

