-- Created on: 1997-05-13
-- Created by: Fabien REUTER
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


package  StlAPI 

    	 ---Purpose : Offers the API for STL data manipulation.
    	 --         

uses 
 
    TopoDS,
    StlMesh
     
is 
    class Writer; 
    class Reader; 
    
    Write(aShape      : in Shape from TopoDS;  
          aFile       : in CString from Standard;
    	  aAsciiMode  : in Boolean from Standard = Standard_True);
	  ---Purpose : Convert and write shape to STL format.
	  --         file is written in binary if aAsciiMode is False
	  --         otherwise it is written in Ascii (by default)

    Read(aShape      : in out Shape from TopoDS;  
          aFile      : CString from Standard);
	  ---Purpose : Create a shape from a STL format.

end  StlAPI;
