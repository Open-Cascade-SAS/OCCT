-- Created on: 2008-12-28
-- Created by: Roman Lygin
-- Copyright (c) 2008-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

--            roman.lygin@gmail.com

generic class CurveCache from Extrema
    (Curve as any; -- Adaptor3d_Curve or Adaptor2d_Curve2d
     Pnt as any;   -- gp_Pnt or gp_Pnt2d
     ArrayOfPnt as Transient from Standard) -- TColgp_HArray1OfPnt or TColgp_HArray1OfPnt2d
inherits Transient from Standard

    ---Purpose:

uses
    Array1OfReal  from TColStd,
    HArray1OfReal from TColStd

raises NotDone from StdFail

is

    Create returns mutable CurveCache from Extrema;

    Create (theC: Curve; theUFirst, theULast: Real; theNbSamples: Integer;
        theToCalculate: Boolean)returns mutable CurveCache from Extrema;

    Create (theC: Curve; theUFirst, theULast: Real;
    	    IntervalsCN: Array1OfReal from TColStd;
	    StartIndex, EndIndex: Integer;
	    Coeff: Real)
    returns mutable CurveCache from Extrema;

    SetCurve (me: mutable; theC: Curve; theNbSamples: Integer;
        theToCalculate: Boolean);
    ---Purpose: Sets the \a theRank-th curve (1 or 2) and its parameters.
    --          Caches sample points for further reuse in Perform().

    SetCurve (me: mutable; theC: Curve;
        theUFirst, theULast: Real; theNbSamples: Integer; theToCalculate: Boolean);
        ---Purpose:

    SetRange (me: mutable; Uinf, Usup: Real; theToCalculate: Boolean);
    ---Purpose:

    CalculatePoints (me: mutable);
    ---Purpose: Calculates points along the curve and stores
    --          them in internal array for further reuse in Perform().

    IsValid (me) returns Boolean;
    ---C++: inline
    ---Purpose: Returns True if the points array has already been calculated
    --          for specified curve and range

    Parameters (me) returns HArray1OfReal from TColStd
        raises  NotDone from StdFail;
    ---C++: inline
    ---C++: return const &
    ---Purpose: Raises StdFail_NotDone if points have not yet been calculated.

    Points (me) returns ArrayOfPnt
        raises  NotDone from StdFail;
    ---C++: inline
    ---C++: return const &
    ---Purpose: Raises StdFail_NotDone if points have not yet been calculated.

    CurvePtr (me) returns Address from Standard;
    ---C++: inline
    ---Purpose:

    NbSamples (me) returns Integer;
    ---C++: inline
    ---Purpose:

    FirstParameter (me) returns Real;
    ---C++: inline
    ---Purpose:

    LastParameter (me) returns Real;
    ---C++: inline
    ---Purpose:

    TrimFirstParameter (me) returns Real;
    ---C++: inline
    ---Purpose: For bounded curves returns FirstParameter(), for unbounded - -1e-10.

    TrimLastParameter (me) returns Real;
    ---C++: inline
    ---Purpose: For bounded curves returns LastParameter(), for unbounded - 1e-10.

fields

    myC           : Address from Standard;
    myFirst       : Real;
    myLast        : Real;
    myTrimFirst   : Real;
    myTrimLast    : Real;
    myNbSamples   : Integer;
    myParamArray  : HArray1OfReal from TColStd;
    myPntArray    : ArrayOfPnt;
    myIsArrayValid: Boolean;

end;
