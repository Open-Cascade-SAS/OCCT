-- Created on: 1993-03-24
-- Created by: JCV
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class Point from Geom2d inherits Geometry from Geom2d

        --- Purpose : The abstract class Point describes the common
    	-- behavior of geometric points in 2D space.
    	-- The Geom2d package also provides the concrete
    	-- class Geom2d_CartesianPoint.

uses Pnt2d from gp

is


  Coord (me; X, Y : out Real) 
        --- Purpose : returns the Coordinates of <me>.
     is deferred;


  Pnt2d (me)  returns Pnt2d
        --- Purpose : returns a non persistent copy of <me>
     is deferred;


  X (me)  returns Real
        --- Purpose : returns the X coordinate of <me>.
     is deferred;


  Y (me)  returns Real
        --- Purpose : returns  the Y coordinate of <me>.
     is deferred;



  Distance (me; Other : Point)  returns Real;
        --- Purpose : computes the distance between <me> and <Other>.

  
  SquareDistance (me; Other : Point)  returns Real;
        --- Purpose : computes the square distance between <me> and <Other>.

end;

