-- Created on: 1998-01-26
-- Created by: Sergey ZARITCHNY
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class EllipseRadiusPresentation from DsgPrs 

	---Purpose: 

uses
    Presentation from Prs3d,
    Pnt          from gp,
    Elips        from gp, 
    OffsetCurve  from Geom,
    Drawer       from Prs3d,
    ArrowSide    from DsgPrs,
    ExtendedString from TCollection

is
      Add( myclass; aPresentation   : Presentation   from Prs3d;
    	    	    aDrawer         : Drawer         from Prs3d; 
		    theval          : Real           from Standard;
		    aText           : ExtendedString from TCollection; 
                    AttachmentPoint : Pnt            from gp;
    	    	    anEndOfArrow    : Pnt            from gp; 
		    aCenter         : Pnt            from gp; 
		    IsMaxRadius     : Boolean        from  Standard;
		    ArrowSide: ArrowSide             from DsgPrs);
		   ---Purpose: draws a  Radius  (Major  or  Minor)   
    	    	   -- representation for whole ellipse  case
		   
    Add( myclass; aPresentation   : Presentation   from Prs3d;
    	    	  aDrawer         : Drawer         from Prs3d; 
		  theval          : Real           from Standard;
		  aText           : ExtendedString from TCollection; 
		  anEllipse       : Elips          from gp;  
                  AttachmentPoint : Pnt            from gp; 
		  anEndOfArrow    : Pnt            from gp; 
		  aCenter         : Pnt            from gp;
		  uFirst          : Real           from Standard;  
		  IsInDomain      : Boolean        from Standard; 
		  IsMaxRadius     : Boolean        from Standard;
	          ArrowSide       : ArrowSide      from DsgPrs);
		   ---Purpose: draws a  Radius  (Major  or  Minor) representation     
    	    	   --  for arc of an ellipse  case 

		   
    Add( myclass; aPresentation   : Presentation   from Prs3d;
    	    	  aDrawer         : Drawer         from Prs3d; 
		  theval          : Real           from Standard;
		  aText           : ExtendedString from TCollection; 
    	    	  aCurve          : OffsetCurve    from Geom;
                  AttachmentPoint : Pnt            from gp; 
		  anEndOfArrow    : Pnt            from gp; 
		  aCenter         : Pnt            from gp;
		  uFirst          : Real           from Standard;  
		  IsInDomain      : Boolean        from Standard; 
		  IsMaxRadius     : Boolean        from Standard;
	          ArrowSide       : ArrowSide      from DsgPrs);
		   ---Purpose: draws a  Radius  (Major  or  Minor) representation     
    	    	   --  for arc of an offset  curve  from  ellipse

end EllipseRadiusPresentation;
