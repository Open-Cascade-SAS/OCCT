-- File:        QuasiUniformCurve.cdl
-- Created:     Mon Dec  4 12:02:30 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWQuasiUniformCurve from RWStepGeom

	---Purpose : Read & Write Module for QuasiUniformCurve

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     QuasiUniformCurve from StepGeom,
     EntityIterator from Interface

is

	Create returns RWQuasiUniformCurve;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable QuasiUniformCurve from StepGeom);

	WriteStep (me; SW : in out StepWriter; ent : QuasiUniformCurve from StepGeom);

	Share(me; ent : QuasiUniformCurve from StepGeom; iter : in out EntityIterator);

end RWQuasiUniformCurve;
