-- File:        OrientedFace.cdl
-- Created:     Fri Dec  1 11:11:23 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class OrientedFace from StepShape 

inherits Face from StepShape 

uses

	Boolean from Standard, 
	HArray1OfFaceBound from StepShape, 
	FaceBound from StepShape, 
	HAsciiString from TCollection
is

	Create returns mutable OrientedFace;
	---Purpose: Returns a OrientedFace


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aBounds : mutable HArray1OfFaceBound from StepShape) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aFaceElement : mutable Face from StepShape;
	      aOrientation : Boolean from Standard) is virtual;

	-- Specific Methods for Field Data Access --

	SetFaceElement(me : mutable; aFaceElement : mutable Face);
	FaceElement (me) returns mutable Face;
	SetOrientation(me : mutable; aOrientation : Boolean);
	Orientation (me) returns Boolean;
	SetBounds(me : mutable; aBounds : mutable HArray1OfFaceBound) is redefined;
	Bounds (me) returns mutable HArray1OfFaceBound is redefined;
	BoundsValue (me; num : Integer) returns mutable FaceBound is redefined;
	NbBounds (me) returns Integer is redefined;

fields

	faceElement : Face from StepShape;
	orientation : Boolean from Standard;

 -- 
 -- NB : field <bounds> inherited from classe <face> is redeclared.
 --      it shall appears in a physical file as a *.
 --

end OrientedFace;
