-- Created on: 2000-05-10
-- Created by: Andrey BETENEV
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1

class ExternalIdentificationItem from StepAP214
inherits SelectType from StepData

    ---Purpose: Representation of STEP SELECT type ExternalIdentificationItem

uses
    DocumentFile from StepBasic,
    ExternallyDefinedClass from StepAP214,
    ExternallyDefinedGeneralProperty from StepAP214,
    ProductDefinition from StepBasic

is
    Create returns ExternalIdentificationItem from StepAP214;
	---Purpose: Empty constructor

    CaseNum (me; ent: Transient) returns Integer;
	---Purpose: Recognizes a kind of ExternalIdentificationItem select type
	--          1 -> DocumentFile from StepBasic
	--          2 -> ExternallyDefinedClass from StepAP214
	--          3 -> ExternallyDefinedGeneralProperty from StepAP214
	--          4 -> ProductDefinition from StepBasic
	--          0 else

    DocumentFile (me) returns DocumentFile from StepBasic;
	---Purpose: Returns Value as DocumentFile (or Null if another type)

    ExternallyDefinedClass (me) returns ExternallyDefinedClass from StepAP214;
	---Purpose: Returns Value as ExternallyDefinedClass (or Null if another type)

    ExternallyDefinedGeneralProperty (me) returns ExternallyDefinedGeneralProperty from StepAP214;
	---Purpose: Returns Value as ExternallyDefinedGeneralProperty (or Null if another type)

    ProductDefinition (me) returns ProductDefinition from StepBasic;
	---Purpose: Returns Value as ProductDefinition (or Null if another type)

end ExternalIdentificationItem;
