-- Created on: 1994-06-16
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class FileName from HeaderSection 

inherits TShared from MMgt

uses

	HAsciiString from TCollection, 
	HArray1OfHAsciiString from Interface
is

	Create returns mutable FileName;
	---Purpose: Returns a FileName

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aTimeStamp : mutable HAsciiString from TCollection;
	      aAuthor : mutable HArray1OfHAsciiString from Interface;
	      aOrganization : mutable HArray1OfHAsciiString from Interface;
	      aPreprocessorVersion : mutable HAsciiString from TCollection;
	      aOriginatingSystem : mutable HAsciiString from TCollection;
	      aAuthorisation : mutable HAsciiString from TCollection);

	-- Specific Methods for Field Data Access --

	SetName(me : mutable; aName : mutable HAsciiString);
	Name (me) returns mutable HAsciiString;
	SetTimeStamp(me : mutable; aTimeStamp : mutable HAsciiString);
	TimeStamp (me) returns mutable HAsciiString;
	SetAuthor(me : mutable; aAuthor : mutable HArray1OfHAsciiString);
	Author (me) returns mutable HArray1OfHAsciiString;
	AuthorValue (me; num : Integer) returns mutable HAsciiString;
	NbAuthor (me) returns Integer;
	SetOrganization(me : mutable; aOrganization : mutable HArray1OfHAsciiString);
	Organization (me) returns mutable HArray1OfHAsciiString;
	OrganizationValue (me; num : Integer) returns mutable HAsciiString;
	NbOrganization (me) returns Integer;
	SetPreprocessorVersion(me : mutable; aPreprocessorVersion : mutable HAsciiString);
	PreprocessorVersion (me) returns mutable HAsciiString;
	SetOriginatingSystem(me : mutable; aOriginatingSystem : mutable HAsciiString);
	OriginatingSystem (me) returns mutable HAsciiString;
	SetAuthorisation(me : mutable; aAuthorisation : mutable HAsciiString);
	Authorisation (me) returns mutable HAsciiString;

fields

	name : HAsciiString from TCollection;
	timeStamp : HAsciiString from TCollection;
	author : HArray1OfHAsciiString from Interface;
	organization : HArray1OfHAsciiString from Interface;
	preprocessorVersion : HAsciiString from TCollection;
	originatingSystem : HAsciiString from TCollection;
	authorisation : HAsciiString from TCollection;

end FileName;
