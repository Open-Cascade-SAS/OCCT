-- File:        OuterBoundaryCurve.cdl
-- Created:     Fri Dec  1 11:11:23 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class OuterBoundaryCurve from StepGeom 

inherits BoundaryCurve from StepGeom 

uses

	HAsciiString from TCollection, 
	HArray1OfCompositeCurveSegment from StepGeom, 
	Logical from StepData
is

	Create returns mutable OuterBoundaryCurve;
	---Purpose: Returns a OuterBoundaryCurve


end OuterBoundaryCurve;
