-- Created on: 2001-09-11
-- Created by: Julia DOROVSKIKH
-- Copyright (c) 2001-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package XmlMXCAFDoc

        ---Purpose: Storage and Retrieval drivers for modelling attributes.
        --          Transient attributes are defined in package XCAFDoc

uses TopLoc,
     XmlMDF,
     XmlObjMgt,
     TDF,
     CDM,
     TopTools

is
    class AreaDriver;

    class CentroidDriver;

    class ColorDriver;

    class GraphNodeDriver;

    class LocationDriver;

    class VolumeDriver;

    class DatumDriver;
    class DimTolDriver;
    class MaterialDriver;

    class ColorToolDriver;
    class DocumentToolDriver;
    class LayerToolDriver;
    class ShapeToolDriver;
    class DimTolToolDriver;
    class MaterialToolDriver;

    AddDrivers (aDriverTable : ADriverTable  from XmlMDF;
                anMsgDrv     : MessageDriver from CDM);
        ---Purpose: Adds the attribute drivers to <aDriverTable>.

end XmlMXCAFDoc;
