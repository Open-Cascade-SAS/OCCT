-- Created by: Peter KURNEV
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ShapeSet from BOPTools 

	---Purpose: Implementation of some formal   
    	--          opereations with a set of shapes        

uses 
    Shape from TopoDS, 
    Edge from TopoDS,
    ShapeEnum from TopAbs,  
    BaseAllocator from BOPCol, 
    MapOfOrientedShape from BOPCol, 
    ListOfShape from BOPCol 
    
--raises

is 
    Create 
    	returns ShapeSet from BOPTools;  
    ---C++: alias "virtual ~BOPTools_ShapeSet();"  
    ---C++: inline 
     
    Create (theAllocator: BaseAllocator from BOPCol)
    	returns ShapeSet from BOPTools; 
    ---C++: inline   
     
    SetShape(me:out; 
    	    theS:Shape from TopoDS); 
    ---C++: inline  
     
    Shape(me) 
    	 returns Shape from TopoDS; 
    ---C++: return const & 
    ---C++: inline  
    
    Add(me:out; 
    	    theLS:ListOfShape from BOPCol);  
	    
    Add(me:out; 
    	    theShape:Shape from TopoDS); 
    ---C++: inline 

    Add(me:out; 
    	    theShape:Shape from TopoDS; 
    	    theType: ShapeEnum from TopAbs); 
	     
    AddEdge(me:out; 
    	    theEdge:Edge from TopoDS); 
    ---C++: inline 

    AddEdges(me:out; 
    	    theLS:ListOfShape from BOPCol);  

    AddEdges(me:out; 
    	    theFace:Shape from TopoDS); 
    ---C++: inline 
     
    Subtract(me:out; 
	    theSet:ShapeSet from BOPTools); 
    ---C++: alias operator -=
    ---C++: inline  
    
    Clear(me:out);
    ---C++: inline 
    
    Get(me; 
	    theLS:out ListOfShape from BOPCol);     
    ---C++: inline 
    
    Contains(me; 
	    theSet:ShapeSet from BOPTools) 
    	returns Boolean from Standard; 
    ---C++: inline
    
     
fields  
    myShape: Shape from TopoDS is protected;   
    myMap  : MapOfOrientedShape from BOPCol is protected;   
	    
end ShapeSet; 
