-- Created on: 1994-03-07
-- Created by: Joelle CHAUVET
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Modified:	Thu Jul  2 16:47:35 1998
--		add methods Generated and GeneratedShapes





class Generator from BRepFill

    	   ---Purpose: Compute a topological surface ( a  shell) using
    	   --          generating wires. The face of the shell will be
    	   --          ruled surfaces passing by the wires.
    	   --          The wires must have the same number of edges.
						    	

uses

    Wire            from TopoDS,
    Shell           from TopoDS,
    Shape           from TopoDS,
    SequenceOfShape from TopTools,
    ListOfShape from TopTools, 
    DataMapOfShapeListOfShape from TopTools


is 
    
    Create returns Generator from BRepFill;
    
    AddWire( me   : in out;
    	     Wire : in Wire from TopoDS)
    is static;
    
    Perform( me     : in out)
	---Purpose: Compute the  shell.
    is static;
    
    Shell(me)
	---C++: return const&
	---C++: inline      
    returns Shell from TopoDS
    is static;
    
    Generated (me )
        ---Purpose: Returns  all   the shapes created 
        ---C++ : return const &          
    returns DataMapOfShapeListOfShape from TopTools
    is static;			 
    
    GeneratedShapes (me ;
    	    	     SSection : Shape from TopoDS)
        ---Purpose: Returns   the  shapes  created  from   a  subshape
        --          <SSection>  of a  section.
        --	
        ---C++ : return const &          
    returns ListOfShape from TopTools
    is static;			 
    



fields
    myWires : SequenceOfShape from TopTools;
    myShell : Shell           from TopoDS;
    myMap   : DataMapOfShapeListOfShape from TopTools;  

end Generator;




