-- File:	TDF_DefaultDeltaOnRemoval.cdl
--      	-----------------------------
-- Author:	DAUTRY Philippe
--		<fid@fox.paris1.matra-dtv.fr>
---Copyright:	 MATRA DATAVISION 1997

---Version:	0.0
---History:	Version	Date		Purpose
--		0.0	Oct 10 1997	Creation


class DefaultDeltaOnRemoval from TDF
    inherits DeltaOnRemoval from TDF

	---Purpose: This class provides a default implementation of a
	--          TDF_DeltaOnRemoval.

uses

    Label     from TDF,
    Attribute from TDF
    
-- raises

is

    Create(anAttribute : Attribute from TDF);
	---Purpose: Creates a TDF_DefaultDeltaOnRemoval.

    Apply (me : mutable)
    	is redefined virtual;
    	---Purpose: Applies the delta to the attribute.

end DefaultDeltaOnRemoval;
