-- Created on: 1998-04-08
-- Created by: Andre LIEUTIER
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



package NLPlate

uses
     Plate, Geom, TCollection, TColStd,
     math, gp, TColgp,  GeomAbs
is

    class NLPlate;
-- Constraints Class
    deferred  class HGPPConstraint; 
    class  HPG0Constraint; 
    class  HPG0G1Constraint;
    class  HPG0G2Constraint;
    class  HPG0G3Constraint;
    class  HPG1Constraint;
    class  HPG2Constraint;
    class  HPG3Constraint;
--  

-- utilities and internal Classes
    class StackOfPlate instantiates Stack from TCollection  
                                       (Plate from Plate);   
    class SequenceOfHGPPConstraint instantiates Sequence from TCollection  
                                       (HGPPConstraint);   
end NLPlate;
