-- Created on: 1992-05-21
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



generic class IntConicCurveGen from IntCurve (
             TheImpTool     as any; -- as ImpTool from IntImpParGen
             ThePCurve      as any;
             ThePCurveTool  as any; -- as ParTool from IntImpParGen(ThePCurve)
	     TheProjPCur    as any) -- as ProjPCurGen(TheCurve,TheCurveTool)
 
inherits Intersection from IntRes2d
		       

	---Purpose: Generic algorithm to intersect a conic from gp and
	--          a parametric  curve.  This class  uses   the class
	--          IConicTool    from  IntCurve,    and  Domain  from
	--          IntCurve.  The  template class for  the PCurveTool
	--          is  given in  the package IntImpParGen  (ParTool).
	--          The  methods  used  to   know  the result  of  the
	--          intersection  are  inherited  from   the     class
	--          Intersection from IntRes2d.
	-- 
	--          This algorithm is called from the IntCurveCurveGen 
	--          class.

        ---Level: Internal

uses IConicTool from IntCurve,
     Lin2d   from gp,
     Circ2d  from gp,
     Elips2d from gp,
     Parab2d from gp,
     Hypr2d  from gp,
     Domain  from IntRes2d



        class TheIntersector    instantiates   Intersector from IntImpParGen(
	           TheImpTool,
		   ThePCurve,
		   ThePCurveTool,
    	    	   TheProjPCur);
        
is

    Create
    
	---Purpose: Empty constructor.

    	returns IntConicCurveGen from IntCurve;
	---C++:inline


    Create (L: Lin2d from gp; D1: Domain from IntRes2d;
            PCurve: ThePCurve; D2: Domain from IntRes2d;
    	    TolConf,Tol: Real from Standard)

	---Purpose: Intersection between a line and a parametric curve.

      	returns IntConicCurveGen from IntCurve;
	---C++:inline 


    Create (C: Circ2d from gp; D1: Domain from IntRes2d;
            PCurve: ThePCurve; D2: Domain from IntRes2d;
    	    TolConf,Tol: Real from Standard)

	---Purpose: Intersection between a line and a parametric curve.

    	returns IntConicCurveGen from IntCurve;



    Create (E: Elips2d from gp; D1: Domain from IntRes2d;
            PCurve: ThePCurve; D2: Domain from IntRes2d;
    	    TolConf,Tol: Real from Standard)

	---Purpose: Intersection between an ellipse and a parametric curve.

    	returns IntConicCurveGen from IntCurve;



    Create (Prb: Parab2d from gp; D1: Domain from IntRes2d;
            PCurve: ThePCurve; D2: Domain from IntRes2d;
    	    TolConf,Tol: Real from Standard)

	---Purpose: Intersection between a parabola and a parametric curve.

    	returns IntConicCurveGen from IntCurve;



    Create (H: Hypr2d from gp; D1: Domain from IntRes2d;
            PCurve: ThePCurve; D2: Domain from IntRes2d;
    	    TolConf,Tol: Real from Standard)

	---Purpose: Intersection between the main branch of an hyperbola
	--          and a parametric curve.

    	returns IntConicCurveGen from IntCurve;



    Perform (me: in out;
             L: Lin2d from gp; D1: Domain from IntRes2d;
             PCurve: ThePCurve; D2: Domain from IntRes2d;
    	     TolConf,Tol: Real from Standard)

	---Purpose: Intersection between a line and a parametric curve.
        ---C++:inline

    	is static;


    Perform (me: in out;
             C: Circ2d from gp; D1: Domain from IntRes2d;
             PCurve: ThePCurve; D2: Domain from IntRes2d;
       	     TolConf,Tol: Real from Standard)

	---Purpose: Intersection between a line and a parametric curve.
        ---C++:inline

    	is static;


    Perform (me: in out;
             E: Elips2d from gp; D1: Domain from IntRes2d;
             PCurve: ThePCurve; D2: Domain from IntRes2d;
       	     TolConf,Tol: Real from Standard)
        ---C++: inline
	---Purpose: Intersection between an ellipse and a parametric curve.

    	is static;


    Perform (me: in out;
             Prb: Parab2d from gp; D1: Domain from IntRes2d;
             PCurve: ThePCurve; D2: Domain from IntRes2d;
       	     TolConf,Tol: Real from Standard)
        ---C++: inline
	---Purpose: Intersection between a parabola and a parametric curve.

    	is static;


    Perform (me: in out; 
             H: Hypr2d from gp; D1: Domain from IntRes2d;
             PCurve: ThePCurve; D2: Domain from IntRes2d;
       	     TolConf,Tol: Real from Standard)

	---Purpose: Intersection between the main branch of an hyperbola
	--          and a parametric curve.
        ---C++: inline

    	is static;


    Perform (me: in out; 
             ICurve: IConicTool from IntCurve; D1: Domain from IntRes2d;
             PCurve: ThePCurve; D2: Domain from IntRes2d;
       	     TolConf,Tol: Real from Standard)
        ---C++:inline
	---Purpose: Intersection between a conic fom gp
	--          and a parametric curve.

    	is static private;


end IntConicCurveGen;
 
