-- Created on: 1994-12-16
-- Created by: Frederic MAUPAS
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Tool from StepToTopoDS

    ---Purpose: This Tool Class provides Information to build
    --          a Cas.Cad BRep from a ProSTEP Shape model.  

uses

    DataMapOfTRI                  from StepToTopoDS,
    PointPair                     from StepToTopoDS,
    PointVertexMap                from StepToTopoDS,
    PointEdgeMap                  from StepToTopoDS,
    TopologicalRepresentationItem from StepShape,
    CartesianPoint                from StepGeom,
    Edge                          from TopoDS,
    Vertex                        from TopoDS,
    Shape                         from TopoDS,
    Curve                         from Geom2d,
    Curve                         from Geom,
    Surface                       from Geom,
    TransientProcess              from Transfer
is

    Create returns Tool from StepToTopoDS;
    
    Create(Map : DataMapOfTRI from StepToTopoDS;
	   TP  : TransientProcess from Transfer)
    	returns Tool from StepToTopoDS;
    
    Init(me : in out;
    	 Map : DataMapOfTRI from StepToTopoDS;
	 TP  : TransientProcess from Transfer);

    IsBound(me   : in out;
    	    TRI  : TopologicalRepresentationItem from StepShape) 
    	returns Boolean from Standard;
	
    Bind(me  : in out;
	 TRI : TopologicalRepresentationItem from StepShape;
    	 S   : Shape from TopoDS);
	 
    Find(me  : in out;
     	 TRI : TopologicalRepresentationItem from StepShape) 
    	returns Shape from TopoDS;
    	---C++: return const &
    
    ClearEdgeMap(me : in out);
    
    IsEdgeBound(me : in out;
    	    	PP : PointPair from StepToTopoDS)
    	returns Boolean from Standard;
	
    BindEdge(me : in out;
    	     PP : PointPair from StepToTopoDS;
	     E  : Edge from TopoDS);
	     
    FindEdge(me : in out;
    	     PP : PointPair from StepToTopoDS)
	returns Edge from TopoDS;
	---C++: return const &
    
    ClearVertexMap(me : in out);
    	    	 
    IsVertexBound(me : in out;
    	    	  PG : CartesianPoint from StepGeom)
    	returns Boolean from Standard;
	
    BindVertex(me : in out;
    	       P  : CartesianPoint from StepGeom;
	       V  : Vertex from TopoDS);
	     
    FindVertex(me : in out;
    	       P  : CartesianPoint from StepGeom)
	returns Vertex from TopoDS;
	---C++: return const &


    ComputePCurve(me : in out;
    	    	  B  : Boolean from Standard);

    ComputePCurve(me) returns Boolean from Standard;    
    
    TransientProcess(me) returns TransientProcess from Transfer;

    -- Statistics

    AddContinuity  (me : in out; GeomSurf  : Surface from Geom);
    AddContinuity  (me : in out; GeomCurve : Curve   from Geom);
    AddContinuity  (me : in out; GeomCur2d : Curve   from Geom2d);

    
    C0Surf(me) returns Integer from Standard;
    C1Surf(me) returns Integer from Standard;
    C2Surf(me) returns Integer from Standard;

    C0Cur2(me) returns Integer from Standard;
    C1Cur2(me) returns Integer from Standard;
    C2Cur2(me) returns Integer from Standard;
    
    C0Cur3(me) returns Integer from Standard;
    C1Cur3(me) returns Integer from Standard;
    C2Cur3(me) returns Integer from Standard;
    
fields

    myDataMap   : DataMapOfTRI     from StepToTopoDS;
    
    myVertexMap : PointVertexMap   from StepToTopoDS;
    
    myEdgeMap   : PointEdgeMap     from StepToTopoDS;

    myComputePC : Boolean          from Standard;
    
    myTransProc : TransientProcess from Transfer;

    -- Statistics : 
    -- Surface continuity 
	     
    myNbC0Surf  : Integer             from Standard;
    myNbC1Surf  : Integer             from Standard;
    myNbC2Surf  : Integer             from Standard;

    -- Curve2d continuity 
	     
    myNbC0Cur2  : Integer             from Standard;
    myNbC1Cur2  : Integer             from Standard;
    myNbC2Cur2  : Integer             from Standard;    

    -- Curve3d continuity 
	     
    myNbC0Cur3  : Integer             from Standard;
    myNbC1Cur3  : Integer             from Standard;
    myNbC2Cur3  : Integer             from Standard;    

end Tool;
