-- Created on: 2001-12-13
-- Created by: Peter KURNEV
-- Copyright (c) 2001-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PntOnFace from IntTools 

	---Purpose: Contains a Face, a 3d point, corresponded UV parameters and a flag

uses
    Face from TopoDS, 
    Pnt  from  gp
--raises

is 
    Create 
    	returns PntOnFace from IntTools;  
	---Purpose:
	--- Empty constructor
	---

    Init(me:out;  
    	 aF: Face from TopoDS; 
	 aP: Pnt  from  gp; 
	 U : Real from  Standard;     
	 V : Real from  Standard); 
	---Purpose:
	--- Initializes me by aFace, a 3d point
	--- and it's UV parameters on face
	---
	
    SetFace(me:out; 
    	    aF:Face from TopoDS); 
	---Purpose:
	--- Modifier
	---
	
    SetPnt (me:out; 
    	    aP:Pnt  from  gp);
    	---Purpose:
	--- Modifier
	---

    SetParameters (me:out; 
	    	   U : Real from  Standard;     
	    	   V : Real from  Standard);
    	---Purpose:
	--- Modifier
	---
	
    SetValid(me:out; 
	     bF : Boolean from Standard); 
    	---Purpose:
	--- Modifier
	---
	    	 
    Valid(me) 
	returns Boolean from Standard; 
	---Purpose:
	--- Selector
	---
	 
    Face(me) 
    	returns Face from TopoDS; 
    	---C++:  return const & 
	---Purpose:
	--- Selector
	---
     
    Pnt (me) 
    	returns Pnt  from gp; 
    	---C++:  return const & 
	---Purpose:
	--- Selector
	---

    Parameters (me; 
	    	U :out Real from Standard;     
	    	V :out Real from Standard); 
    	---Purpose:
	--- Selector
	---
	  
    IsValid(me) 
	returns Boolean from Standard; 
	---Purpose:
	--- Selector

fields  

    myIsValid : Boolean from Standard;    
    myPnt : Pnt  from  gp; 
    myU   : Real from  Standard;        
    myV   : Real from  Standard;        
    myFace: Face from TopoDS; 
end PntOnFace;
