-- Created on: 1994-11-18
-- Created by: Marie Jose MARTZ
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class GeomVector from GeomToIGES inherits GeomEntity from GeomToIGES

    ---Purpose: This class implements the transfer of the Vector from Geom
    --          to IGES . These can be :
    --          . Vector
    --              * Direction
    --              * VectorWithMagnitude
  
uses
 
    Vector               from Geom,
    VectorWithMagnitude  from Geom,
    Direction            from Geom,
    Direction            from IGESGeom,
    GeomEntity           from GeomToIGES
     
is 
    
    Create returns GeomVector from GeomToIGES;


    Create(GE : GeomEntity from GeomToIGES)  
    	 returns GeomVector from GeomToIGES;
    ---Purpose : Creates a tool GeomVector ready to run and sets its
    --         fields as GE's.

    TransferVector   (me    : in out;
                      start : Vector from Geom)
    	 returns mutable Direction from IGESGeom;
    ---Purpose :  Transfert  a  GeometryEntity which  answer True  to  the
    --            member : BRepToIGES::IsGeomVector(Geometry).  If this
    --            Entity could not be converted, this member returns a NullEntity.


    TransferVector   (me    : in out;
                      start : VectorWithMagnitude from Geom)
    	 returns mutable Direction from IGESGeom;


    TransferVector   (me    : in out;
                      start : Direction from Geom)
    	 returns mutable Direction from IGESGeom;


end GeomVector;


