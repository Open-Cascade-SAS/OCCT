-- Created on: 1993-01-08
-- Created by: Philippe DAUTRY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



deferred generic class Builder from Sweep(TheShape as any)
    

	---Purpose: This  is   a  signature class  describing services
	--          strictly required    by  the    Swept   Primitives
	--          algorithms, from the Topology Data Structure .
	--          


uses

    Orientation from TopAbs
is

    MakeCompound (me; aCompound : out TheShape)
    	---Purpose: Returns an empty Compound.
    is deferred;

    MakeCompSolid (me; aCompSolid : out TheShape)
    	---Purpose: Returns an empty CompSolid.
    is deferred;

    MakeSolid (me; aSolid : out TheShape)
    	---Purpose: Returns an empty Solid.
    is deferred;

    MakeShell (me; aShell : out TheShape)
    	---Purpose: Returns an empty Shell.
    is deferred;

    MakeWire (me; aWire : out TheShape)
    	---Purpose: Returns an empty Wire.
    is deferred;
    
    Add(me; aShape1 : in out TheShape; 
	    aShape2 : in     TheShape;
    	    Orient  : in     Orientation from TopAbs)
    	---Purpose: Adds the Shape 1 in the Shape 2, set to
    	--          <Orient> orientation.
    is deferred;
    
    Add(me; aShape1 : in out TheShape; 
	    aShape2 : in     TheShape)
    	---Purpose: Adds the Shape 1 in the Shape 2.
    is deferred;

end Builder from Sweep;


