-- Created on: 1994-02-18
-- Created by: Remi LEQUETTE
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- modified by Michael KLOKOV  Wed Mar  6 15:01:25 2002

class Section from BRepAlgoAPI  
    inherits BooleanOperation from BRepAlgoAPI
      
    ---Purpose:  
    -- The algorithm is to build a Secton operation between arguments and tools. 
    -- The result of Section operation consists of vertices and edges. 
    -- The result of Section operation contains:
    -- 1. new vertices that are subjects of V/V, E/E, E/F, F/F interferences
    -- 2. vertices that are subjects of V/E, V/F interferences
    -- 3. new edges that are subjects of F/F interferences
    -- 4. edges that are Common Blocks

    -- The vertex is included in Section only when it is not shared 
    -- between the edges above 
    --  --  
   
    -- Default values:
    --   - geometries built are NOT approximated.
    --   - PCurves are NOT computed on both parts.
      
    -- Example of use:
    -- Standard_Boolean bRunParallel; 
    -- Standard_Integer iErr;
    -- BRepAlgoAPI_Section aSection; 
    -- //  
    -- bRunParallel=...;  //  turn  parallelism on/off 
    -- const TopTools_ListOfShape&  aLS=...;  //  Arguments 
    -- const TopTools_ListOfShape&  aLT=...;  //  Tools 
    -- // 
    -- aSection.SetRunParallel();  
    -- aSection.SetArguments(aLS);
    -- aSection.SetTools(aLT); 
    -- aSection.Approximation(Standard_True);
    -- // 
    -- aSection.Build();  // perform the algorithm     
    -- iErr=pBuilder->ErrorStatus();
    -- if (iErr) {
    --   // errors  occured 
    --   return 0;
    -- }  
    -- // 
    -- const TopoDS_Shape& aR=aSection.Shape();// the result 
    -- //... 
     
    
uses
    Pln   from gp,
    Shape from TopoDS,
    Surface from Geom,
    Curve   from Geom2d,
    PaveFiller from BOPAlgo, 
    Operation from BOPAlgo,
    ListOfShape from TopTools, 
    BaseAllocator from BOPCol
    
is
    Create 
        returns Section from BRepAlgoAPI;   
    ---C++: alias "Standard_EXPORT virtual ~BRepAlgoAPI_Section();"  
    --- Purpose: Empty constructor 
  
    Create (PF: PaveFiller from BOPAlgo)
        returns Section from BRepAlgoAPI;  
    --- Purpose: Empty constructor    
    -- <PF> - PaveFiller object that is carried out  
      
    Create(S1 : Shape from TopoDS; 
           S2 : Shape from TopoDS;
           PerformNow : Boolean = Standard_True) 
        returns Section from BRepAlgoAPI;
    ---Purpose: Constructor with two shapes  
    -- <S1>  -argument     
    -- <S2>  -tool   
    -- <PerformNow> - the flag: 
    -- if <PerformNow>=True - the algorithm is performed immediatly 
    -- Obsolete   
     
    Create (S1 : Shape from TopoDS;  
            S2 : Shape from TopoDS; 
            aDSF:PaveFiller from BOPAlgo;
            PerformNow : Boolean = Standard_True)  
        returns Section from BRepAlgoAPI;
    ---Purpose: Constructor with two shapes  
    -- <S1>  -argument     
    -- <S2>  -tool   
    -- <PF> - PaveFiller object that is carried out        
    -- <PerformNow> - the flag: 
    -- if <PerformNow>=True - the algorithm is performed immediatly 
    -- Obsolete   

    Create(S1 : Shape from TopoDS;  
           Pl : Pln from gp;
           PerformNow : Boolean = Standard_True) 
        returns Section from BRepAlgoAPI;
    ---Purpose: Constructor with two shapes  
    -- <S1>  - argument
    -- <Pl>  - tool  
    -- <PerformNow> - the flag: 
    -- if <PerformNow>=True - the algorithm is performed immediatly 
    -- Obsolete   
     

    Create(S1 : Shape from TopoDS;  
           Sf : Surface from Geom;
           PerformNow : Boolean = Standard_True) 
        returns Section from BRepAlgoAPI;
     ---Purpose: Constructor with two shapes   
     -- <S1>  - argument
     -- <Sf>  - tool  
     -- <PerformNow> - the flag: 
     -- if <PerformNow>=True - the algorithm is performed immediatly 
     -- Obsolete    
     

    Create(Sf : Surface from Geom;  
           S2 : Shape from TopoDS;
           PerformNow : Boolean = Standard_True) 
        returns Section from BRepAlgoAPI;
     ---Purpose: Constructor with two shapes   
     -- <Sf>  - argument
     -- <S2>  - tool  
     -- <PerformNow> - the flag: 
     -- if <PerformNow>=True - the algorithm is performed immediatly 
     -- Obsolete
 
    Create(Sf1 : Surface from Geom;  
           Sf2 : Surface from Geom;
           PerformNow : Boolean = Standard_True) 
        returns Section from BRepAlgoAPI;
     ---Purpose:  
     ---Purpose: Constructor with two shapes   
     -- <Sf1>  - argument
     -- <Sf2>  - tool  
     -- <PerformNow> - the flag: 
     -- if <PerformNow>=True - the algorithm is performed immediatly 
     -- Obsolete 

    Init1(me : out; 
            S1 : Shape from TopoDS);
    ---Purpose: initialize the argument  
    -- <S1>  - argument
    -- Obsolete 
     
    Init1(me : out; 
            Pl : Pln from gp); 
    ---Purpose: initialize the argument  
    -- <Pl>  - argument
    -- Obsolete  
        
    Init1(me : out; 
            Sf : Surface from Geom);
    ---Purpose: initialize the argument 
    -- <Sf>  - argument
    -- Obsolete 
     
    Init2(me : out; 
            S2 : Shape from TopoDS);
    ---Purpose: initialize the tool 
    -- <S2>  - tool
    -- Obsolete 
     
    Init2(me : out; 
            Pl : Pln from gp);
    ---Purpose: initialize the tool 
    -- <Pl>  - tool
    -- Obsolete  
 
    Init2(me : out; 
            Sf : Surface from Geom);
    ---Purpose: initialize the tool 
    -- <Sf>  - tool
    -- Obsolete   
    
    Approximation(me : out; 
        B : Boolean from Standard);
    ---Purpose:  
    --Defines an option for computation
    -- of further intersections. 
    -- By default, the underlying 3D geometry attached to each
    -- elementary edge of the result is:
    -- - analytic where possible, provided the corresponding
    --   geometry corresponds to a type of analytic curve defined in
    -- - or elsewhere, given as a succession of points grouped
    --   together in a BSpline curve of degree 1.  
    --   If Approx equals true, these edges will have an attached 3D
    --   geometry which is a BSpline approximation of the computed
    --   set of points.
    --   Note that as a result, approximations will be computed
    --   on edges built only on new intersection curves.
 
    ComputePCurveOn1(me : out; 
        B : Boolean from Standard);
    ---Purpose: 
    -- Indicates whether the P-Curve should be (or not)  
    -- performed on the argument. 
    -- By default, no parametric 2D curve (pcurve) is defined for the
    -- edges of the result.  
    -- If ComputePCurve1 equals true, further computations performed  
    -- to attach an P-Curve in the parametric space of the argument  
    -- to the constructed edges. 
    -- Obsolete   
 
    ComputePCurveOn2(me : out; 
            B : Boolean from Standard);
    ---Purpose:  
    -- Indicates whether the P-Curve should be (or not)  
    -- performed on the tool.  
    -- By default, no parametric 2D curve (pcurve) is defined for the
    -- edges of the result.  
    -- If ComputePCurve1 equals true, further computations performed  
    -- to attach an P-Curve in the parametric space of the tool  
    -- to the constructed edges.
    -- Obsolete   
     
    Build(me : in out) 
        is redefined;   
    ---Purpose: Performs the algorithm 
    -- Filling interference Data Structure (if it is necessary)
    -- Building the result of the operation. 
 
    HasAncestorFaceOn1(me;  
            E : Shape from TopoDS;
            F : out Shape from TopoDS)
        returns Boolean from Standard;
     ---Purpose:
     -- get the face of the first part giving section edge <E>.
     -- Returns True on the 3 following conditions :
     -- 1/ <E> is an edge returned by the Shape() metwod. 
     -- 2/ First part of section performed is a shape.
     -- 3/ <E> is built on a intersection curve (i.e <E>
     --   is not the result of common edges)
     -- When False, F remains untouched.
    -- Obsolete   
    
    HasAncestorFaceOn2(me;  
            E : Shape from TopoDS;
            F : out Shape from TopoDS)
        returns Boolean from Standard;
     ---Purpose:  Identifies the ancestor faces of
     -- the intersection edge E resulting from the last
     -- computation performed in this framework, that is, the faces of
     -- the two original shapes on which the edge E lies:
     -- -      HasAncestorFaceOn1 gives the ancestor face in the first shape, and
     -- -      HasAncestorFaceOn2 gives the ancestor face in the second shape.
     --   These functions return true if an ancestor face F is found, or false if not.
     --   An ancestor face is identifiable for the edge E if the following
     -- conditions are satisfied:
     -- -  the first part on which this algorithm performed its
     --    last computation is a shape, that is, it was not given as
     -- a surface or a plane at the time of construction of this
     -- algorithm or at a later time by the Init1 function,
     -- - E is one of the elementary edges built by the
     -- last computation of this section algorithm.
     -- To use these functions properly, you have to test the returned
     -- Boolean value before using the ancestor face: F is significant
     -- only if the returned Boolean value equals true.
    -- Obsolete   
     
    --
    --  protected methods 
    --
    Init(me: out; 
            PerformNow : Boolean) 
        is protected;
    
    SetAttributes (me:out) 
        is redefined protected;   
 
fields
    myParametersChanged : Boolean from Standard;
    myApprox            : Boolean from Standard;
    myComputePCurve1    : Boolean from Standard;
    myComputePCurve2    : Boolean from Standard;
    
end Section from BRepAlgoAPI;
