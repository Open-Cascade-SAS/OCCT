-- Created on: 1998-07-28
-- Created by: LECLERE Florence
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class FuseFace from TopOpeBRepBuild

	---Purpose: 

uses Shape                     from TopoDS,
     Face                      from TopoDS,
     Edge                      from TopoDS,
     Vertex                    from TopoDS,
     DataMapOfShapeListOfShape from TopTools,
     ListOfShape               from TopTools


is


    Create
    	returns FuseFace from TopOpeBRepBuild;
    	---C++: inline
    	--   
	
	
    Create(LIF : ListOfShape from TopTools;
   	   LRF : ListOfShape from TopTools;     
	   CXM : Integer from Standard)
	   
    	---C++: inline
    	--      
    	returns FuseFace from TopOpeBRepBuild;


    Init(me: in out; LIF : ListOfShape from TopTools;
	       	     LRF : ListOfShape from TopTools;
	    	     CXM : Integer from Standard)    
    	is static;


    PerformFace(me: in out)
  
    	is static;


    PerformEdge(me: in out)
  
    	is static;

    ClearEdge(me: in out)
    
    	is static;
	
    ClearVertex(me: in out)
    
    	is static;
	
    IsDone(me)
    
    	returns Boolean from Standard
	---C++: inline
	is static;	
	
    IsModified(me)
    
    	returns Boolean from Standard
	---C++: inline
	is static;	
	    
    LFuseFace(me)
    
        returns ListOfShape from TopTools
	---C++: return const&
    	is static;

    LInternEdge(me)
    
        returns ListOfShape from TopTools
	---C++: return const&
    	is static;
	
    LExternEdge(me)
    
        returns ListOfShape from TopTools
	---C++: return const&
    	is static;
	
    LModifEdge(me)
    
        returns ListOfShape from TopTools
	---C++: return const&
    	is static;
	
    LInternVertex(me)
    
        returns ListOfShape from TopTools
	---C++: return const&
    	is static;
	
    LExternVertex(me)
    
        returns ListOfShape from TopTools
	---C++: return const&
    	is static;
	
    LModifVertex(me)
    
        returns ListOfShape from TopTools
	---C++: return const&
    	is static;
	
		
fields

    myLIF      : ListOfShape               from TopTools;
    myLRF      : ListOfShape               from TopTools;
    myLFF      : ListOfShape               from TopTools;
    
    myLIE      : ListOfShape               from TopTools is protected;
    myLEE      : ListOfShape               from TopTools is protected;
    myLME      : ListOfShape               from TopTools is protected;
        
    myLIV      : ListOfShape               from TopTools is protected;
    myLEV      : ListOfShape               from TopTools is protected;
    myLMV      : ListOfShape               from TopTools is protected;

    myInternal : Boolean                   from Standard; 
    myModified : Boolean                   from Standard;
    myDone     : Boolean                   from Standard;
    
end FuseFace;    
