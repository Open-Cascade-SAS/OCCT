-- Created on: 1995-04-20
-- Created by: Tony GEORGIADES
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

--		Modified Tue Sep 19 1995 by Jean-Louis Frenkel
--		Modified Tue Jan 19 1999 by Louis Dusuzeau

package Resource
    ---Purpose: Resources management.
    --          A RESOURCE is a parameter saved on a file and used to
    --          initialize a variable.

uses
    TCollection,MMgt,SortTools,TColStd
is 

   enumeration FormatType is     
    	SJIS,
	EUC,
	ANSI,
	GB
   end FormatType ;
    	---Purpose:
    	-- List of non ASCII format types which may be
    	-- converted into the Unicode 16 bits format type.
    	-- Use the functions provided by the
    	-- Resource_Unicode class to convert a string
    	-- from one of these non ASCII format to Unicode, and vice versa.

   class DataMapOfAsciiStringAsciiString instantiates
    	 DataMap from TCollection(AsciiString from TCollection,
	    	    	    	 AsciiString from TCollection,
	    	    	    	 AsciiString from TCollection) ;

   class DataMapOfAsciiStringExtendedString instantiates
    	 DataMap from TCollection(AsciiString from TCollection,
	    	    	    	  ExtendedString from TCollection,
	    	    	    	  AsciiString from TCollection) ;
	 
   class QuickSortOfArray1 instantiates
    	 QuickSort from SortTools(AsciiString from TCollection,
    	    	    	    	  Array1OfAsciiString from TColStd,
	    	    	    	  LexicalCompare from Resource) ;
				  
---Class:
   class LexicalCompare ;
   
   class Manager;
   ---Purpose: Defines a resource structure and its management methods.

   class Unicode;

   exception NoSuchResource inherits NoSuchObject from Standard;

end Resource;
