-- Created on: 1991-09-02
-- Created by: NW,JPB,CAL
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


deferred class AspectMarker from Aspect

inherits

	TShared

	---Purpose: This class allows the definition of a group
	--	    of attributes for the primitive MARKER.
	--	    the attributes are:
	--		* Colour
	--		* Type
	--		* Scale factor
	--	    When any value of the group is modified
	--	    all graphic objects using the group are modified

uses

	Color		from Quantity,

	TypeOfMarker 	from Aspect

raises

	AspectMarkerDefinitionError 	from Aspect

is

	Initialize;
	---Level: Public
	---Purpose: Initialise the constructor for Graphic3d_AspectMarker3d.
	--
	-- defaults values :
	--
	--	Color	= Quantity_NOC_YELLOW;
	--	Type	= Aspect_TOM_X;
	--	Scale	= 1.0;

	Initialize ( AColor	: Color from Quantity;
		     AType	: TypeOfMarker from Aspect;
		     AScale	: Real from Standard )
	---Level: Public
	---Purpose: Initialise the values for the
	--	    constructor of Graphic3d_AspectMarker3d.
	--  Warning: Raises AspectMarkerDefinitionError if the
	--	    scale is a negative value.
	raises AspectMarkerDefinitionError from Aspect;

	---------------------------------------------------
	-- Category: Methods to modify the class definition
	---------------------------------------------------

	SetColor ( me		: mutable;
		   AColor	: Color from Quantity );
	---Level: Public
	---Purpose: Modifies the colour of <me>.
	---Category: Methods to modify the class definition

	SetScale ( me		: mutable;
		   AScale	: Real from Standard )
	---Level: Public
	---Purpose: Modifies the scale factor of <me>.
	--	    Marker type Aspect_TOM_POINT is not affected
	--	    by the marker size scale factor. It is always
	--	    the smallest displayable dot.
	--  Warning: Raises AspectMarkerDefinitionError if the
	--	    scale is a negative value.
	raises AspectMarkerDefinitionError from Aspect;

	SetType ( me	: mutable;
		  AType	: TypeOfMarker from Aspect );
	---Level: Public
	---Purpose: Modifies the type of marker <me>.
	---Category: Methods to modify the class definition

	----------------------------
	-- Category: Inquire methods
	----------------------------

	Values ( me;
		 AColor	: out Color from Quantity;
		 AType	: out TypeOfMarker from Aspect;
		 AScale	: out Real from Standard );
	---Level: Public
	---Purpose: Returns the current values of the group <me>.
	---Category: Inquire methods

--

fields

--
-- Class	:	Aspect_AspectMarker
--
-- Purpose	:	Declaration of variables specific to the context of
--			drawing markers
--
-- Reminder	:	A drawing context for markers is defined by :
--			- the colour
--			- the type
--			- the scale
--

	-- the colour
	MyColor	:	Color from Quantity;

	-- the type
	MyType	:	TypeOfMarker from Aspect;

	-- the scale
	MyScale	:	Real from Standard;

end AspectMarker;
