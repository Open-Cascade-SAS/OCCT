-- Created on: 1995-12-06
-- Created by: Frederic MAUPAS
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class BoxCharacteristicSelect from StepVisual

    -- Hand made Select Type

uses

    Real from Standard
    
is

    Create returns BoxCharacteristicSelect;
    
    TypeOfContent(me) returns Integer from Standard;
    -- 1 box_height,
    -- 2 box_width,
    -- 3 box_slant_angle,
    -- 4 box_rotate_angle)

    SetTypeOfContent(me : in out; aType : Integer from Standard);
    
    RealValue(me) returns Real from Standard;
    
    SetRealValue(me : in out; aValue : Real from Standard);
    
fields

    theRealValue     : Real from Standard;
    theTypeOfContent : Integer from Standard;
    
end BoxCharacteristicSelect;
