-- Created on: 2000-08-11
-- Created by: Andrey BETENEV
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Style from XCAFPrs 

    ---Purpose: Represents a set of styling settings applicable to 
    --          a (sub)shape

uses
    Color from Quantity

is

    Create returns Style from XCAFPrs;  

    IsSetColorSurf (me) returns Boolean;  
    GetColorSurf (me) returns Color from Quantity;  
    SetColorSurf (me: in out; col: Color from Quantity);  
    UnSetColorSurf (me: in out);  
    	---Purpose: Manage surface color setting

    IsSetColorCurv (me) returns Boolean;  
    GetColorCurv (me) returns Color from Quantity;  
    SetColorCurv (me: in out; col: Color from Quantity);  
    UnSetColorCurv (me: in out);  
    	---Purpose: Manage curve color setting

    SetVisibility(me: in out; visibility: Boolean from Standard);
    IsVisible(me) returns Boolean;
    	---Purpose: Manage visibility
	--          Note: Setting visibility to False makes colors undefined
	--          This is necessary for HashCode

    IsEqual (me; other: Style from XCAFPrs) returns Boolean;
    	---Purpose: Returs True if styles are the same
	---C++: alias operator ==

    ---Purpose: Methods for using Style as key in maps

    HashCode(myclass; S : Style from XCAFPrs; Upper : Integer) returns Integer;
	---Purpose: Returns a HasCode value  for  the  Key <K>  in the
	--          range 0..Upper.
	
    IsEqual(myclass; S1, S2 : Style from XCAFPrs) returns Boolean;
	---Purpose: Returns True  when the two  keys are the same. Two
	--          same  keys  must   have  the  same  hashcode,  the
	--          contrary is not necessary.
	
fields

--    defColor:     Boolean;
    defColorSurf: Boolean;
    defColorCurv: Boolean;
    myVisibility: Boolean from Standard;

--    myColor:     Color from Quantity;
    myColorSurf: Color from Quantity;
    myColorCurv: Color from Quantity;
    

end Style;
