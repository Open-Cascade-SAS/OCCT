-- Created on: 2000-08-15
-- Created by: Andrey BETENEV
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Reader from STEPCAFControl 
-- inherits Reader from STEPControl

    ---Purpose: Provides a tool to read STEP file and put it into
    --          DECAF document. Besides transfer of shapes (including 
    --          assemblies) provided by STEPControl, supports also 
    --          colors and part names
    --
    --          This reader supports reading files with external references
    --          i.e. multifile reading
    --          It behaves as usual Reader (from STEPControl) for the main
    --          file (e.g. if it is single file)
    --          Results of reading other files can be accessed by name of the
    --          file or by iterating on a readers

uses
    AsciiString from TCollection,
    WorkSession from XSControl,
    ReturnStatus from IFSelect,
    Shape from TopoDS,
    Document from TDocStd,
    Reader from STEPControl,
    NextAssemblyUsageOccurrence from StepRepr,
    DictionaryOfExternFile from STEPCAFControl,
    ExternFile from STEPCAFControl,
    ExternRefs from STEPConstruct,
    Tool from STEPConstruct,
    DataMapOfShapePD from STEPCAFControl,
    DataMapOfPDExternFile from STEPCAFControl,
    DataMapOfShapeLabel from XCAFDoc,
    MapOfShape from TopTools,
    ShapeTool from XCAFDoc,
    Label from TDF,
    LabelSequence from TDF,
    HSequenceOfTransient from TColStd,
    RepresentationItem from StepRepr,
    TransientProcess from Transfer,
    ConnectedFaceSet from StepShape

is

    Create returns Reader;
    	---Purpose: Creates a reader with an empty
-- STEP model and sets ColorMode, LayerMode, NameMode and
-- PropsMode to Standard_True.

    Create (WS : mutable WorkSession from XSControl;
    	    	 scratch : Boolean = Standard_True) returns Reader;
    	---Purpose: Creates a reader tool and attaches it to an already existing Session
    	-- 	    Clears the session if it was not yet set for STEP

    Init (me: in out; WS : mutable WorkSession from XSControl;
    	       	      scratch : Boolean = Standard_True);
    	---Purpose: Clears the internal data structures and attaches to a new session
    	--          Clears the session if it was not yet set for STEP

    ReadFile (me : in out; filename : CString) 
    returns ReturnStatus from IFSelect;
        ---Purpose: Loads a file and returns the read status
	--          Provided for use like single-file reader

    NbRootsForTransfer (me: in out) returns Integer;
    	---Purpose: Returns number of roots recognized for transfer
	--          Shortcut for Reader().NbRootsForTransfer()

    TransferOneRoot (me: in out; num: Integer; doc: in out Document from TDocStd) 
    returns Boolean;
    	---Purpose: Translates currently loaded STEP file into the document
	--          Returns True if succeeded, and False in case of fail
	--          Provided for use like single-file reader

    Transfer (me: in out; doc: in out Document from TDocStd) 
    returns Boolean;
    	---Purpose: Translates currently loaded STEP file into the document
	--          Returns True if succeeded, and False in case of fail
	--          Provided for use like single-file reader

    Perform (me: in out; filename: AsciiString from TCollection; 
    	    	         doc: in out Document from TDocStd) returns Boolean;

    Perform (me: in out; filename: CString; doc: in out Document from TDocStd) 
    returns Boolean;
    	---Purpose: Translate STEP file given by filename into the document
	--          Return True if succeeded, and False in case of fail

    ---Scope: Access to fields
    
    ExternFiles (me) returns DictionaryOfExternFile from STEPCAFControl;
    	---Purpose: Returns data on external files
	--          Returns Null handle if no external files are read
	---C++: return const &
	
    ExternFile (me; name: CString; ef: out ExternFile from STEPCAFControl)
    returns Boolean;
    	---Purpose: Returns data on external file by its name
	--          Returns False if no external file with given name is read
	
    ChangeReader (me: in out) returns Reader from STEPControl;
    	---Purpose: Returns basic reader 
	---C++: return &

    Reader (me) returns Reader from STEPControl;
    	---Purpose: Returns basic reader as const
	---C++: return const &

    ---Scope: Internal methods

    Transfer (me: in out; rd: in out Reader from STEPControl; 
    	    	    	  num: Integer;
                          doc: in out Document from TDocStd;
			  Lseq: out LabelSequence from TDF;
    	    	    	  asOne: Boolean = Standard_False)
    returns Boolean is protected;
    	---Purpose: Translates STEP file already loaded into the reader 
        --          into the document
	--          If num==0, translates all roots, else only root number num
	--          Returns True if succeeded, and False in case of fail
	--          If asOne is True, in case of multiple results composes
        --          them into assembly. Fills sequence of produced labels

    AddShape (me; S: Shape from TopoDS; STool: ShapeTool from XCAFDoc;
                  NewShapesMap : MapOfShape from TopTools;
    	    	  ShapePDMap: DataMapOfShapePD from STEPCAFControl;
    	    	  PDFileMap : DataMapOfPDExternFile from STEPCAFControl;
    	    	  ShapeLabelMap: in out DataMapOfShapeLabel from XCAFDoc)
    returns Label from TDF is protected;
    	---Purpose: Add a shape to a document
	--          Depending on a case, this shape can be added as one, or
	--          as assembly, or (in case if it is associated with external
	--          reference) taken as that referred shape

    ReadExternFile (me: in out; file, fullpath: CString; doc: in out Document from TDocStd) 
    returns ExternFile from STEPCAFControl is protected;
    	---Purpose: Reads (or if returns already read) extern file with 
	--          given name

    ReadColors (me; WS: WorkSession from XSControl;
                    doc: in out Document from TDocStd;
		    PDFileMap : DataMapOfPDExternFile from STEPCAFControl;
    	    	    ShapeLabelMap: DataMapOfShapeLabel from XCAFDoc)
    returns Boolean is protected;
    	---Purpose: Reads style assignments from STEP model and sets
	--          corresponding color assignments in the DECAF document

    ReadNames (me; WS: WorkSession from XSControl; 
                   doc: in out Document from TDocStd;
    	    	   PDFileMap : DataMapOfPDExternFile from STEPCAFControl;
    	    	   ShapeLabelMap: DataMapOfShapeLabel from XCAFDoc) 
    returns Boolean is protected;
    	---Purpose: Reads names of parts defined in the STEP model and 
	--          assigns them to corresponding labels in the DECAF document

    ReadValProps (me; WS: WorkSession from XSControl; 
                      doc: in out Document from TDocStd;
    	    	      PDFileMap : DataMapOfPDExternFile from STEPCAFControl;
    	    	      ShapeLabelMap: DataMapOfShapeLabel from XCAFDoc)
    returns Boolean is protected;
    	---Purpose: Reads validation properties assigned to shapes in the STEP 
        --          model and assigns them to corresponding labels in the DECAF 
        --          document

    ReadLayers (me; WS: WorkSession from XSControl; 
                   doc: in out Document from TDocStd) 
    returns Boolean is protected;
    	---Purpose: Reads layers of parts defined in the STEP model and 
	--          set reference between shape and layers in the DECAF document

    ReadSHUOs (me; WS: WorkSession from XSControl;
                   doc: in out Document from TDocStd;
    	    	   PDFileMap : DataMapOfPDExternFile from STEPCAFControl;
    	    	   ShapeLabelMap: DataMapOfShapeLabel from XCAFDoc)
    returns Boolean is protected;
    	---Purpose: Reads SHUO for instances defined in the STEP model and 
	--          set reference between shape instances from different assemblyes 

    ReadGDTs (me; WS: WorkSession from XSControl;
                  doc: in out Document from TDocStd)
    returns Boolean is protected;
    	---Purpose: Reads D&GT for instances defined in the STEP model and 
	--          set reference between shape instances from different assemblyes 

    ReadMaterials (me; WS: WorkSession from XSControl;
                       doc: in out Document from TDocStd;
    	               SeqPDS : HSequenceOfTransient from TColStd)
    returns Boolean is protected;
    	---Purpose: Reads materials for instances defined in the STEP model and 
	--          set reference between shape instances from different assemblyes 

    SettleShapeData(me; theItem: RepresentationItem from StepRepr;
                        theLab: out Label from TDF;
                        theShapeTool: ShapeTool from XCAFDoc;
                        theTP: TransientProcess from Transfer)
    returns Label from TDF is protected;
    --- Purpose: Populates the sub-Label of the passed TDF Label with shape
     --          data associated with the given STEP Representation Item,
     --          including naming and topological information.

    ExpandSubShapes(me; theShapeTool: ShapeTool from XCAFDoc;
                        theShapeLabelMap: DataMapOfShapeLabel from XCAFDoc;
                        theShapePDMap: DataMapOfShapePD from STEPCAFControl)
    is protected;
    --- Purpose: Given the maps of already translated shapes, this method
     --          expands their correspondent Labels in XDE Document so that
     --          to have a dedicated sub-Label for each sub-shape coming
     --          with associated name in its STEP Representation Item.

    ExpandManifoldSolidBrep(me; theLab: out Label from TDF;
                                theItem: RepresentationItem from StepRepr;
                                theTP: TransientProcess from Transfer;
                                theShapeTool: ShapeTool from XCAFDoc)
    is protected;
    ---  Purpose: Expands the topological structure of Manifold Solid BRep
     --           STEP entity to OCAF sub-tree. Entities having no names
     --           associated via their Representation Items are skipped.

    ExpandSBSM(me; theLab: out Label from TDF;
               theItem: RepresentationItem from StepRepr;
               theTP: TransientProcess from Transfer;
               theShapeTool: ShapeTool from XCAFDoc)
    is protected;
    ---  Purpose: Expands the topological structure of Shell-Based Surface
     --           Model STEP entity to OCAF sub-tree. Entities having no names
     --           associated via their Representation Items are skipped.

    ExpandShell(me; theShell: ConnectedFaceSet from StepShape;
                    theLab: out Label from TDF;
                    theTP: TransientProcess from Transfer;
                    theShapeTool: ShapeTool from XCAFDoc)
    is protected;
    ---  Purpose: Expands STEP Shell structure to OCAF sub-tree. Entities
     --           having no names associated via their Representation Items
     --           are skipped.

    FindInstance (myclass; NAUO: NextAssemblyUsageOccurrence from StepRepr;
                      STool: ShapeTool from XCAFDoc;
     	    	      Tool: Tool from STEPConstruct; 
    	    	      PDRFileMap : DataMapOfPDExternFile from STEPCAFControl;
    	    	      ShapeLabelMap: DataMapOfShapeLabel from XCAFDoc)
    returns Label from TDF;
    	---Purpose: Returns label of instance of an assembly component
	--          corresponding to a given NAUO

    --- Work with fileds for different mode of reading STEP file.

    SetColorMode(me: in out; colormode: Boolean from Standard);
    	---Purpose: Set ColorMode for indicate read Colors or not.

    GetColorMode(me) returns Boolean;

    SetNameMode(me: in out; namemode: Boolean from Standard);
    	---Purpose: Set NameMode for indicate read Name or not.
    
    GetNameMode(me) returns Boolean;

    SetLayerMode(me: in out; layermode: Boolean from Standard);
    	---Purpose: Set LayerMode for indicate read Layers or not.

    GetLayerMode(me) returns Boolean; 

    
    SetPropsMode(me: in out; propsmode: Boolean from Standard);
    	---Purpose: PropsMode for indicate read Validation properties or not.

    GetPropsMode(me) returns Boolean;
	
    SetSHUOMode(me: in out; shuomode: Boolean from Standard);
    	---Purpose: Set SHUO mode for indicate write SHUO or not.

    GetSHUOMode(me) returns Boolean;
	
    SetGDTMode(me: in out; gdtmode: Boolean from Standard);
    	---Purpose: Set GDT mode for indicate write GDT or not.

    GetGDTMode(me) returns Boolean;
	
    SetMatMode(me: in out; matmode: Boolean from Standard);
    	---Purpose: Set Material mode

    GetMatMode(me) returns Boolean;
	
fields

    myReader : Reader from STEPControl;
    myFiles  : DictionaryOfExternFile from STEPCAFControl;
    myColorMode : Boolean;
    myNameMode  : Boolean;
    myLayerMode : Boolean;
    myPropsMode : Boolean;
    mySHUOMode  : Boolean;
    myGDTMode   : Boolean;
    myMatMode   : Boolean;

end Reader;
