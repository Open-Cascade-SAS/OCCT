-- Created on: 1997-02-10
-- Created by: Odile Olivier
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

--  SAV : OCC218 06/03/02 : Add(...) overloaded to take into account arrow & text
--                          aspects.

class XYZAxisPresentation from DsgPrs
    	---Purpose: A framework for displaying the axes of an XYZ trihedron.
uses

    Presentation from Prs3d,
    LineAspect   from Prs3d,
    Pnt          from gp,
    Dir          from gp,
    ArrowAspect from Prs3d,
    TextAspect from Prs3d

is

    Add(myclass;
    	aPresentation: Presentation from Prs3d;
    	anLineAspect : LineAspect from Prs3d;
    	aDir         : Dir from gp;
	aVal         : Real from Standard;
	aText        : CString from Standard;
    	aPfirst      : Pnt    from gp;
    	aPlast       : Pnt    from gp);
	 
    	---Purpose: Draws each axis of a trihedron displayed in the
    	-- presentation aPresentation and with lines shown by
    	-- the values of aLineAspect. Each axis is defined by:
    	-- -   the first and last points aPfirst and aPlast
    	-- -   the direction aDir and
    	-- -   the value aVal which provides a value for length.
    	--  The value for length is provided so that the trihedron
    	-- can vary in length relative to the scale of shape display.
    	-- Each axis will be identified as X, Y, or Z by the text aText.


    Add(myclass;
    	aPresentation : Presentation from Prs3d;
    	aLineAspect   : LineAspect from Prs3d;
    	anArrowAspect : ArrowAspect from Prs3d;
    	aTextAspect   : TextAspect from Prs3d;
    	aDir          : Dir from gp;
	aVal          : Real from Standard;
	aText         : CString from Standard;
    	aPfirst       : Pnt    from gp;
    	aPlast        : Pnt    from gp);
	 
    	---Purpose: draws the presentation X ,Y ,Z axis

end XYZAxisPresentation;
