-- Created on: 1992-09-23
-- Created by: Christian CAILLET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Cumulate  from IFGraph  inherits GraphContent

    	---Purpose : this class evaluates effect of cumulated sub-parts :
    	--           overlapping, forgotten entities
    	--           Results are kept in a Graph, several question can be set
    	--           Basic Iteration gives entities which are part of Cumulation

uses Transient, EntityIterator, Graph

is

    Create (agraph : Graph) returns Cumulate;
    ---Purpose : creates empty Cumulate, ready to work

    GetFromEntity (me : in out; ent : any Transient);
    ---Purpose : adds an entity and its shared ones to the list

    GetFromIter (me : in out; iter : EntityIterator);
    ---Purpose : adds a list of entities (as an iterator) as such, that is,
    --           without their shared entities (use AllShared to have them)

    ResetData (me : in out);
    ---Purpose : Allows to restart on a new data set

    	-- --   Results   -- --
    	--   More-Next-Value-Entity give all entities taken into the Cumulation
    	--   other informations are provided, as EntityIterator : hence they
    	--   are available for other evaluations

    Evaluate (me : in out) is redefined;
    ---Purpose : Evaluates the result of cumulation

    Overlapped (me) returns EntityIterator;
    ---Purpose : returns entities which are taken several times

    Forgotten (me) returns EntityIterator;
    ---Purpose : returns entities which are not taken

    PerCount (me; count : Integer = 1) returns EntityIterator;
    ---Purpose : Returns entities taken a given count of times
    --           (0 : same as Forgotten, 1 : same as no Overlap : default)

    NbTimes (me; ent : Transient) returns Integer;
    ---Purpose : returns number of times an Entity has been counted
    --           (0 means forgotten, more than 1 means overlap, 1 is normal)

    HighestNbTimes (me) returns Integer;
    ---Purpose : Returns the highest number of times recorded for every Entity
    --           (0 means empty, 1 means no overlap)

fields

    thegraph : Graph;

end Cumulate;
