-- Created on: 1995-09-21
-- Created by: Philippe GIRODENGO
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package StlMesh 

	---Purpose: Implements a  basic  mesh data-structure  for  the
	--          needs of the application fast prototyping.
	--          

uses  

    MMgt,  
    TCollection,  
    TColStd,  
    gp,  
    TColgp

is

    class Mesh;
    	---Purpose: Mesh definition.  The mesh contains one or several
    	--          domains. Each  mesh   domain  contains a  set   of
    	--          triangles. Each domain can have its own deflection
    	--          value.


    class MeshExplorer;
    	---Purpose: Provides   facilities to explore  the triangles of
    	--          each mesh domain.
    

    class MeshDomain;
    	---Purpose: Set of triangles defined with three vertices and a
    	--          given orientation. Internal class used to classify
    	--          the triangles of each domain.


    class MeshTriangle;
        ---Purpose: triangle defined with three vertices and a given 
        --          orientation

    

    class SequenceOfMeshDomain  instantiates
          Sequence from TCollection (MeshDomain from StlMesh);



    class SequenceOfMeshTriangle  instantiates
          Sequence from TCollection (MeshTriangle from StlMesh);
    
    
    class SequenceOfMesh instantiates
    	  Sequence from TCollection (Mesh from StlMesh);
	  ---Purpose: Sequence of meshes
    
    Merge (mesh1, mesh2 : in Mesh) returns Mesh;
    ---Purpose: Make a merge of two Mesh and returns a new Mesh.
    --          Very useful if you want to merge partMesh and CheckSurfaceMesh
    --          for example

end StlMesh;
