-- File:        SiUnitAndRatioUnit.cdl
-- Created:     Mon Dec  4 12:02:36 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWSiUnitAndRatioUnit from RWStepBasic

	---Purpose : Read & Write Module for SiUnitAndRatioUnit

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     SiUnitAndRatioUnit from StepBasic

is

	Create returns RWSiUnitAndRatioUnit;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable SiUnitAndRatioUnit from StepBasic);

	WriteStep (me; SW : in out StepWriter; ent : SiUnitAndRatioUnit from StepBasic);

end RWSiUnitAndRatioUnit;
