-- Created on: 1993-07-06
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Curve3D from PBRep inherits GCurve from PBRep

	---Purpose: Representation of a curve by a 3D curve.

uses

    Location from PTopLoc,
    Curve    from PGeom

is

    Create(C  : Curve    from PGeom;
    	   CF : Real     from Standard;
	   CL : Real     from Standard;
    	   L  : Location from PTopLoc) 
    returns mutable Curve3D from PBRep;
    	---Purpose : CF is curve first param
    	--           CL is curve last param
    	--           As far as they can't be computed from a Persistent Curve
    	--          they are given in the Curve3D constructor

    Curve3D(me) returns Curve from PGeom
    is static;

    IsCurve3D(me) returns Boolean
	 ---Purpose: Returns True.
    is redefined;
	
fields
    
    myCurve3D : Curve from PGeom;

end Curve3D;
