-- File:      HLRAppli_ReflectLines.cdl
-- Created:   05.12.12 15:53:35
-- Created by: Julia GERASIMOVA
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class ReflectLines from HLRAppli

        ---Purpose : This class builds reflect lines on a shape
        --         according to the axes of view defined by user.
        --         Reflect lines are represented by edges in 3d.


uses
    Shape from TopoDS,
    Projector from HLRAlgo
    
is 
    Create(aShape : Shape from TopoDS)
    ---Purpose: Constructor
    --
    returns ReflectLines from HLRAppli;
    
    SetAxes(me: in out;
    	    Nx,  Ny,  Nz  : Real from Standard;
    	    XAt, YAt, ZAt : Real from Standard;
	    XUp, YUp, ZUp : Real from Standard);
	---Purpose: Sets the normal to the plane of visualisation,
	--          the coordinates of the view point and
	--          the coordinates of the vertical direction vector.

    Perform(me: in out);
    
    GetResult(me)
    returns Shape from TopoDS;
	---Purpose: returns resulting compound of reflect lines
	--          represented by edges in 3d
   
fields

    myProjector : Projector from HLRAlgo;
    myShape     : Shape     from TopoDS;
    myCompound  : Shape     from TopoDS;
    
end ReflectLines;
