-- Created on: 1993-04-20
-- Created by: Modelistation
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class CLPropsATool from HLRBRep

uses
    Curve from HLRBRep,
    Pnt2d from gp,
    Vec2d from gp

is
    Value(myclass; A :     Address from Standard;
                   U :     Real    from Standard;
                   P : out Pnt2d   from gp);
    	---Purpose: Computes the  point <P> of  parameter <U>   on the
    	--          Curve from HLRBRep <C>.
    	--
    	---C++: inline          
         	
    D1   (myclass; A  :     Address from Standard;
                   U  :     Real    from Standard;
                   P  : out Pnt2d   from gp;
                   V1 : out Vec2d   from gp);
    	---Purpose: Computes the point <P>  and  first derivative <V1>
    	--          of parameter <U> on the curve <C>.
    	--
    	---C++: inline          

    D2   (myclass; A      :     Address from Standard;
                   U      :     Real    from Standard;
                   P      : out Pnt2d   from gp;
                   V1, V2 : out Vec2d from gp);
    	---Purpose: Computes the point <P>,  the first derivative <V1>
    	--          and second derivative <V2> of parameter <U> on the
    	--          curve <C>.
    	--
    	---C++: inline          
    
    D3   (myclass; A          :     Address from Standard;
                   U          :     Real    from Standard; 
                   P          : out Pnt2d   from gp;
                   V1, V2, V3 : out Vec2d   from gp);
    	---Purpose: Computes the point <P>, the first derivative <V1>,
    	--          the second derivative  <V2>   and third derivative
    	--          <V3> of parameter <U> on the curve <C>.
    	--
    	---C++: inline          

    Continuity(myclass; A : Address from Standard)
    returns Integer from Standard;
     	---Purpose: returns the order  of continuity of the curve <C>.
     	--          returns 1 :  first  derivative only is  computable
     	--          returns 2  : first and  second derivative only are
     	--          computable.  returns  3 : first,  second and third
     	--          are computable.
    	--
    	---C++: inline          

    FirstParameter(myclass; A : Address from Standard)
    returns Real from Standard;
     	---Purpose: returns the first parameter bound of the curve.
     	--          
    	---C++: inline          
     
    LastParameter(myclass; A : Address from Standard)
    returns Real from Standard;
	---Purpose: returns the  last  parameter bound  of  the curve.
	--          FirstParameter must be less than LastParamenter.
    	--
    	---C++: inline          

end CLPropsATool;
