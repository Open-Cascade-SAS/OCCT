-- Created on: 2000-05-30
-- Created by: Sergey MOZOKHIN
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



package VrmlAPI 

	---Purpose: API for writing to VRML 1.0

uses
    TopoDS,
    VrmlConverter,
    Vrml,
    Quantity
is
    enumeration RepresentationOfShape
    	---Purpose: Identifies the representation of the shape written
    	-- to a VRML file. The available options are :
    	-- -      VrmlAPI_ShadedRepresentation :
    	--    the shape is translated with a shaded representation.
    	-- -      VrmlAPI_WireFrameRepresentation :
    	--   the shape is translated with a wireframe representation.
    	-- -      VrmlAPI_BothRepresentation : the shape is translated
    	--   to VRML format with both representations : shaded and
    	--    wireframe. This is the default option.
        
    is
	    ShadedRepresentation,
	    WireFrameRepresentation,
	    BothRepresentation
    end RepresentationOfShape;

    class Writer;
    	---Purpose: With help of this class user can change parameters of writing.
    
    Write(aShape: Shape from TopoDS; aFileName: CString from Standard);
    	---Purpose: Converts the shape aShape to VRML format and writes it
    	-- to the file identified by aFileName using default parameters.
    
end VrmlAPI;
