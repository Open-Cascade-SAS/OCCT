-- Created by: NW,JPB,CAL
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class AspectLine3d from Graphic3d inherits AspectLine from Aspect

	---Version:

	---Purpose: Creates and updates a group of attributes
	--	    for 3d line primitives. This group contains the
	--	    colour, the type of line, and its thickness.
	

uses

	Color		from Quantity,

	TypeOfLine	from Aspect

is

	Create
		returns mutable AspectLine3d from Graphic3d;
	---Level: Public
	---Purpose: Creates a context table for line primitives
	--	    defined with the following default values:
	--
	--	    Colour	: NOC_YELLOW
	--	    Line type	: TOL_SOLID
	--	    Width	: 1.0

	Create ( AColor	: Color from Quantity;
		 AType	: TypeOfLine from Aspect;
		 AWidth	: Real from Standard )
		returns mutable AspectLine3d from Graphic3d;
	---Level: Public
	---Purpose: Creates a context table for line primitives
	--	    defined with the specified values.
	--  Warning: <AWidth> is the "linewidth scale factor".
	--	    The nominal line width is 1 pixel. The width of
	--	    the line is determined by applying the linewidth scale
	--	    factor to this nominal line width.
	--	    The supported linewidths vary by 1-pixel units.

--

-- fields

--
-- Class	:	Graphic3d_AspectLine3d
--
-- Purpose	:	Declaration of context-specific variables
--			for drawing 3d lines
--
-- Reminder	:	A context for drawing 3d lines inherits:
--			- the colour
--			- the type of line
--			- the thickness
--			defined by AspectLine.
--

end AspectLine3d;
