-- Created on: 1996-03-29
-- Created by: Laurent BOURESCHE
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Constant from Law inherits Function from Law

	---Purpose: Loi constante

uses
    Array1OfReal    from TColStd,
    Shape           from GeomAbs
      
raises OutOfRange from Standard

is

    Create returns mutable Constant from Law;
    
    

    Set(me: mutable; Radius,PFirst,PLast : Real from Standard)
    ---Purpose: Set the radius and the range of the constant Law.
    is static;
		
    Continuity(me) returns Shape from GeomAbs
    	---Purpose: Returns GeomAbs_CN
    is redefined static;
    
    NbIntervals(me; S : Shape from GeomAbs) returns Integer    
	---Purpose: Returns  1
    is redefined static;
    
    Intervals(me; T : in out Array1OfReal from TColStd; 
    	          S : Shape from GeomAbs)
    raises
    	OutOfRange from Standard 
    is redefined static;

    Value(me: mutable; X: Real from Standard)
    ---Purpose: Returns the value at parameter X.
    returns Real from Standard;

    D1(me: mutable; X: Real from Standard; F,D: out Real from Standard);
    ---Purpose: Returns the value and the first derivative at parameter X.

    D2(me: mutable; X: Real from Standard; 
       F,D, D2: out Real from Standard);
    ---Purpose: Returns the value, first and second derivatives 
    --          at parameter X.
    
        
    Trim(me; PFirst, PLast, Tol :Real from Standard) returns Function   
    is redefined static;
    
    Bounds(me: mutable; PFirst,PLast : out Real from Standard);
    ---Purpose: Returns the parametric bounds of the function.

fields

radius : Real from Standard;
first  : Real from Standard;
last   : Real from Standard;

end Constant;
