-- File:        DescriptiveRepresentationItem.cdl
-- Created:     Mon Dec  4 12:02:25 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWDescriptiveRepresentationItem from RWStepRepr

	---Purpose : Read & Write Module for DescriptiveRepresentationItem

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     DescriptiveRepresentationItem from StepRepr

is

	Create returns RWDescriptiveRepresentationItem;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable DescriptiveRepresentationItem from StepRepr);

	WriteStep (me; SW : in out StepWriter; ent : DescriptiveRepresentationItem from StepRepr);

end RWDescriptiveRepresentationItem;
