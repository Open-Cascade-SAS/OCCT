-- Created on: 2003-02-04
-- Created by: data exchange team
-- Copyright (c) 2003-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class ElementOrElementGroup from StepFEA
inherits SelectType from StepData

    ---Purpose: Representation of STEP SELECT type ElementOrElementGroup

uses
    ElementRepresentation from StepFEA,
    ElementGroup from StepFEA

is
    Create returns ElementOrElementGroup from StepFEA;
	---Purpose: Empty constructor

    CaseNum (me; ent: Transient) returns Integer;
	---Purpose: Recognizes a kind of ElementOrElementGroup select type
	--          1 -> ElementRepresentation from StepFEA
	--          2 -> ElementGroup from StepFEA
	--          0 else

    ElementRepresentation (me) returns ElementRepresentation from StepFEA;
	---Purpose: Returns Value as ElementRepresentation (or Null if another type)

    ElementGroup (me) returns ElementGroup from StepFEA;
	---Purpose: Returns Value as ElementGroup (or Null if another type)

end ElementOrElementGroup;
