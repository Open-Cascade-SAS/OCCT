-- File:	AIS_PerpendicularRelation.cdl
-- Created:	Thu Dec  5 09:40:49 1996
-- Author:	Jean-Pierre COMBE/Odile Olivier
--		<odl@sacadox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1996

class PerpendicularRelation from AIS inherits Relation from AIS
    	---Purpose: A framework to display constraints of perpendicularity
    	-- between two or more interactive datums. These
    	-- datums can be edges or faces.
uses Shape                 from TopoDS,
     Presentation          from Prs3d,
     PresentationManager3d from PrsMgr,
     Selection             from SelectMgr,
     Pnt                   from gp,
     Dir                   from gp,
     Projector             from Prs3d,
    Transformation        from Geom,
     PresentationManager2d from PrsMgr,
     GraphicObject         from Graphic2d,     
     Plane                 from Geom

is
    Create (aFShape     : Shape          from TopoDS;
    	    aSShape     : Shape          from TopoDS;
	    aPlane      : Plane          from Geom)
	---Purpose:  Constructs an object to display constraints of
    	-- perpendicularity on shapes.
    	-- This object is defined by a first shape aFShape, a
    	-- second shape aSShape, and a plane aPlane.
    	-- aPlane is the plane of reference to show and test the
    	-- perpendicular relation between two shapes, at least
    	-- one of which has a revolved surface.
    returns mutable PerpendicularRelation from AIS;

    Create (aFShape     : Shape          from TopoDS;
    	    aSShape     : Shape          from TopoDS)
	---Purpose:  Constructs an object to display constraints of
    	-- perpendicularity on shapes.
    	-- This object is defined by a first shape aFShape and a
    	-- second shape aSShape.
    returns mutable PerpendicularRelation from AIS;

-- -- Methods from PresentableObject

    Compute(me            : mutable;
    	    aPresentationManager: PresentationManager3d from PrsMgr;
    	    aPresentation : mutable Presentation from Prs3d;
    	    aMode         : Integer from Standard= 0) 
    is redefined static private;
    
    Compute(me:mutable;
    	        aProjector: Projector from Prs3d;
                aPresentation: mutable Presentation from Prs3d)
    is redefined static private;     

    Compute(me:mutable;
    	    aPresentationManager: PresentationManager2d from PrsMgr;
            aPresentation: mutable GraphicObject from Graphic2d;
            aMode: Integer from Standard = 0)
    is redefined static private;	    

    Compute(me            : mutable;
    	    aProjector    : Projector from Prs3d;
    	    aTrsf         : Transformation from Geom;
	    aPresentation : mutable Presentation from Prs3d)
    is redefined;
    	---Purpose: computes the presentation according to a point of view
    	--          given by <aProjector>. 
    	--          To be Used when the associated degenerated Presentations 
    	--          have been transformed by <aTrsf> which is not a Pure
    	--          Translation. The HLR Prs can't be deducted automatically
    	--          WARNING :<aTrsf> must be applied
    	--           to the object to display before computation  !!!

-- Methods from SelectableObject

    ComputeSelection(me         : mutable;
    	    	     aSelection : mutable Selection from SelectMgr;
    	    	     aMode      : Integer from Standard)is private;


--
--     Computation private methods
--

    ComputeTwoFacesPerpendicular(me: mutable;
    	    	    	         aPresentation : mutable Presentation from Prs3d)
    is private;
    
    ComputeTwoEdgesPerpendicular(me: mutable;
    	    	    	         aPresentation : mutable Presentation from Prs3d)
    is private;
    

fields

    myFAttach     : Pnt from gp;
    mySAttach     : Pnt from gp;
    
end PerpendicularRelation;


