-- Created on: 1991-05-16
-- Created by: Isabelle GRIGNON
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class IntLinTorus from IntAna 

	---Purpose: Intersection between a line and a torus.

uses Lin          from gp,
     Torus        from gp,
     Pnt          from gp

raises NotDone    from StdFail,
       OutOfRange from Standard


is

    Create
    
    	returns IntLinTorus from IntAna;

    Create(L : Lin from gp; T : Torus from gp)
    
    	---Purpose: Creates the intersection between a line and a torus.

    	returns IntLinTorus from IntAna;


    Perform(me: in out; L : Lin from gp; T : Torus from gp)
    
    	---Purpose: Intersects a line and a torus.

    	is static;


    IsDone(me)
    
	---Purpose: Returns True if the computation was successful.
	--          
	---C++: inline

    	returns Boolean from Standard
	
	is static;


    NbPoints(me)
    
    	---Purpose: Returns the number of intersection points.
	--          
	---C++: inline

    	returns Integer from Standard
	
	raises NotDone     from StdFail
    	--     The exception NotDone is raised if IsDone returns False. 

	is static;


    Value(me; Index : Integer from Standard)
    
    	---Purpose: Returns the intersection point of range Index.
	--          
	---C++: inline
	---C++: return const&

    	returns Pnt from gp

    	raises NotDone    from StdFail,
               OutOfRange from Standard
    	--     The exception NotDone is raised if IsDone returns False. 
    	--     The exception OutOfRange is raised if Index <= 0 or
    	--        Index > NbPoints
	
	is static;


    ParamOnLine(me; Index : Integer from Standard)
    
    	---Purpose: Returns the parameter on the line of the intersection
    	--          point of range Index.
	--          
	---C++: inline

    	returns Real from Standard

    	raises NotDone    from StdFail,
               OutOfRange from Standard
    	--     The exception NotDone is raised if IsDone returns False. 
    	--     The exception OutOfRange is raised if Index <= 0 or
    	--        Index > NbPoints
	
	is static;


    ParamOnTorus(me; Index : Integer from Standard;
                     FI,THETA: out Real from Standard)
    
    	---Purpose: Returns the parameters on the torus of the intersection
    	--          point of range Index.
	--          
	---C++: inline

    	raises NotDone    from StdFail,
               OutOfRange from Standard
    	--     The exception NotDone is raised if IsDone returns False. 
    	--     The exception OutOfRange is raised if Index <= 0 or
    	--        Index > NbPoints
	
	is static;


fields

    done    : Boolean      from Standard;
    nbpt    : Integer      from Standard;
    thePoint: Pnt          from gp [4];
    theParam: Real         from Standard [4];
    theFi   : Real         from Standard [4];
    theTheta: Real         from Standard [4];

end IntLinTorus;
