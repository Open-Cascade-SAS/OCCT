-- Created on: 1991-02-21
-- Created by: Isabelle GRIGNON
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class   ExtPElS from Extrema
    	---Purpose: It calculates all the extremum distances
    	--          between a point and a surface.
    	--          These distances can be minimum or maximum.

uses   	POnSurf  from Extrema,
    	Cone     from gp,
	Pln      from gp,
    	Cylinder from gp,
    	Pnt      from gp,
    	Sphere   from gp,
    	Torus    from gp

raises  NotDone from StdFail,
    	OutOfRange

is
    Create returns ExtPElS;
    
    Create (P: Pnt; S: Cylinder; Tol: Real) returns ExtPElS;
      	---Purpose: It calculates all the distances between a point 
      	--          and a cylinder from gp.
      	--          Tol is used to test if the point is on the axis.

    Perform(me: in out; P: Pnt; S: Cylinder; Tol: Real) 
    is static;

    Create (P: Pnt; S: Pln; Tol: Real) returns ExtPElS;
      	---Purpose: It calculates all the distances between a point 
      	--          and a plane from gp.
      	--          Tol is used to test if the point is on the plane.

    Perform(me: in out; P: Pnt; S: Pln; Tol: Real) 
    is static;


    Create (P: Pnt; S: Cone; Tol: Real) returns ExtPElS;
      	---Purpose: It calculates all the distances between a point 
      	--          and a cone from gp.
      	--          Tol is used to test if the point is at the apex or
      	--          on the axis.

    Perform(me: in out;P: Pnt; S: Cone; Tol: Real)
    is static;
    
    Create (P: Pnt; S: Torus; Tol: Real) returns ExtPElS;
      	---Purpose: It calculates all the distances between a point 
      	--          and a torus from gp.
      	--          Tol is used to test if the point is on the axis.
    
    Perform(me: in out; P: Pnt; S: Torus; Tol: Real)
    is static;

    Create (P: Pnt; S: Sphere; Tol: Real) returns ExtPElS;
      	---Purpose: It calculates all the distances between a point 
      	--          and a sphere from gp.
      	--          Tol is used to test if the point is at the center.
    
    Perform(me: in out; P: Pnt; S: Sphere; Tol: Real)
    is static;


    IsDone (me) returns Boolean
    	---Purpose: Returns True if the distances are found.
    	is static;
    
    NbExt (me) returns Integer
    	---Purpose: Returns the number of extremum distances.
    	raises  NotDone from StdFail
	    	-- if IsDone(me)=False.
    	is static;

    SquareDistance (me; N: Integer) returns Real
    	---Purpose: Returns the value of the Nth resulting square distance.
    	raises  NotDone from StdFail,
    	    	-- if IsDone(me)=False.
    	        OutOfRange
		-- if N < 1 or N > NbPoints(me).
    	is static;

    Point (me; N: Integer) returns POnSurf
        ---C++: return const &
    	---Purpose: Returns the point of the Nth resulting distance.
    	raises  NotDone from StdFail,
    	    	-- if IsDone(me)=False.
    	        OutOfRange
		-- if N < 1 or N > NbPoints(me).
    	is static;

fields
    myDone : Boolean;
    myNbExt: Integer;
    mySqDist: Real [4];
    myPoint: POnSurf from Extrema [4];

end ExtPElS;
