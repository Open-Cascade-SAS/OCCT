-- Created by: TCL
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Straightness from Prs2d inherits Tolerance from Prs2d

uses

	GraphicObject   from Graphic2d,
	Drawer          from Graphic2d,
	Length	        from Quantity,
    FStream         from Aspect 

is
	-------------------------
	-- Category: Constructors
	-------------------------

	Create( aGO                    : GraphicObject from Graphic2d;
		    aX, aY                 : Real          from Standard;
		    aLength                : Real          from Standard = 3.0;
            anAngle                : Real          from Standard = 0.0 );
	---Level: Public
	---Purpose: Creates a tolerance straightness with the center at <aX>, <aY>; 
	--          length of this is <aLength>;
	--          reference point is <aXPosition>, <aYPosition>
	---Category: Constructor

    --------------------------
	-- Category: Draw and Pick
	--------------------------

	Draw( me : mutable; aDrawer: Drawer from Graphic2d ) is static protected;
	---Level: Internal
	---Purpose: Draws the straightness <me>.

	Save( me; aFStream: in out FStream from Aspect ) is virtual;

end Straightness from Prs2d;
