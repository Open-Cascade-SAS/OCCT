-- Created on: 1999-10-08
-- Created by: Vladislav ROMASHKO
-- Copyright (c) 1999-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Fillet from QANewBRepNaming inherits TopNaming from QANewBRepNaming

	---Purpose: For topological naming of a fillet

uses

     MakeFillet from BRepFilletAPI,
     Shape      from TopoDS,
     Label      from TDF

is

    Create returns Fillet from QANewBRepNaming;

    Create(ResultLabel : Label from TDF)
    returns Fillet from QANewBRepNaming;

    Init(me : in out; ResultLabel : Label from TDF);


    Load (me; part     :        Shape      from TopoDS;
    	      mkFillet : in out MakeFillet from BRepFilletAPI);
      ---Purpose: Loads a fillet in a data framework

    DeletedFaces(me)
    ---Purpose: Returns a label for deleted faces of the part.
    returns Label from TDF;

    ModifiedFaces(me)
    ---Purpose: Returns a label for modified faces of the part.
    returns Label from TDF;

    FacesFromEdges(me)
    ---Purpose: Returns a label for faces generated from edges of the part.
    returns Label from TDF;

    FacesFromVertices(me)
    ---Purpose: Returns a label for faces generated from vertices of the part.
    returns Label from TDF;

    WRFace1(me)
    ---Purpose: Returns a label for WorkAround Face number 1
    returns Label from TDF;

    WRFace2(me)
    ---Purpose: Returns a label for WorkAround Face number 2
    returns Label from TDF;

    WREdge1(me)
    ---Purpose: Returns a label for WorkAround Edge number 1
    returns Label from TDF;

    WREdge2(me)
    ---Purpose: Returns a label for WorkAround Edge number 2
    returns Label from TDF;


end Fillet;
