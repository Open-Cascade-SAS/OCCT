-- Created on: 1998-05-12
-- Created by: Philippe NOUAILLE
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class AppFuncRstRst from BRepBlend inherits AppFuncRoot from BRepBlend
	---Purpose: Function to approximate by AppSurface for Edge/Face          
	---Level: Advanced

uses 
 Line            from BRepBlend,
 Point           from Blend,
 AppFunction     from Blend,
 RstRstFunction  from Blend,
 Vector          from math

 
raises OutOfRange from  Standard

is   
     
   Create(Line : in out Line from BRepBlend;
    	  Func  : in  out RstRstFunction from Blend; 
          Tol3d: Real;
          Tol2d: Real)
   returns AppFuncRstRst from BRepBlend;

   Point(me;
    	 Func  : AppFunction from Blend; 
	 Param : Real;
	 Sol   : Vector from math;
	 Pnt   : in out Point from Blend);
	
   Vec(me;
       Sol : in out Vector from math;
       Pnt : Point from Blend);
	
end AppFuncRstRst;
