-- Created on: 1995-04-05
-- Created by: Christophe MARION
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class OutLiner from HLRTest inherits Drawable3D from Draw
	---Purpose: 

uses
    OStream,
    Display     from Draw,
    Interpretor from Draw,
    OutLiner    from HLRTopoBRep,
    Shape       from TopoDS

is
    Create(S : Shape from TopoDS)
    returns mutable OutLiner from HLRTest; 
    
    OutLiner(me) returns OutLiner from HLRTopoBRep;
	---C++: inline

    DrawOn(me; dis : in out Display from Draw);
	---Purpose: Does nothhing,
    
    Copy(me) returns mutable Drawable3D from Draw
	---Purpose: For variable copy.
    is redefined;
	
    Dump(me; S : in out OStream)
	---Purpose: For variable dump.
    is redefined;

    Whatis(me; I : in out Interpretor from Draw)
	---Purpose: For variable whatis command. Set  as a result  the
	--          type of the variable.
    is redefined;

fields
    myOutLiner : OutLiner from HLRTopoBRep;

end OutLiner;
