-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class EIR from TopOpeBRepDS 

---Purpose:  EdgeInterferenceReducer

uses

    Shape       from TopoDS,
    Edge        from TopoDS,
    ListOfShape from TopTools,
    IndexedMapOfShape from TopTools,
    Config                            from TopOpeBRepDS,
    Interference                      from TopOpeBRepDS,
    ListOfInterference                from TopOpeBRepDS,
    ListIteratorOfListOfInterference  from TopOpeBRepDS,
    ListOfShapeOn1State               from TopOpeBRepDS,
    DataMapOfShapeListOfShapeOn1State from TopOpeBRepDS,
    HDataStructure                    from TopOpeBRepDS

is

    Create(HDS:HDataStructure) returns EIR from TopOpeBRepDS;
    ProcessEdgeInterferences(me : in out);
    ProcessEdgeInterferences(me : in out; I : Integer);

fields

    myHDS : HDataStructure;
    
end EIR from TopOpeBRepDS;
