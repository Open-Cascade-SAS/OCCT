-- File:	IGESDimen_ToolDimensionTolerance.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolDimensionTolerance  from IGESDimen

    ---Purpose : Tool to work on a DimensionTolerance. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses DimensionTolerance from IGESDimen,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolDimensionTolerance;
    ---Purpose : Returns a ToolDimensionTolerance, ready to work


    ReadOwnParams (me; ent : mutable DimensionTolerance;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : DimensionTolerance;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : DimensionTolerance;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a DimensionTolerance <ent>, from
    --           its specific (own) parameters

    OwnCorrect (me; ent : mutable DimensionTolerance) returns Boolean  is static;
    ---Purpose : Sets automatic unambiguous Correction on a DimensionTolerance
    --           (NbPropertyValues forced to 8)

    DirChecker (me; ent : DimensionTolerance) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : DimensionTolerance;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : DimensionTolerance; entto : mutable DimensionTolerance;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : DimensionTolerance;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolDimensionTolerance;
