-- Created on: 1992-11-18
-- Created by: Christian CAILLET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class SelectAnyType  from IFSelect  inherits SelectExtract

    ---Purpose : A SelectAnyType sorts the Entities of which the Type is Kind
    --           of a given Type : this Type for Match is specific of each
    --           class of SelectAnyType

uses Type, InterfaceModel

is

    TypeForMatch (me) returns Type  is deferred;
    ---Purpose : Returns the Type which has to be matched for select

    Sort (me; rank : Integer; ent : Transient; model : InterfaceModel)
    	returns Boolean;
    ---Purpose : Returns True for an Entity (model->Value(num)) which is kind
    --           of the choosen type, given by the method TypeForMatch.
    --           Criterium is IsKind.

end SelectAnyType;
