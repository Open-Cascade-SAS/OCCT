-- Created on: 1996-10-11
-- Created by: Christian CAILLET
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SelectSubordinate  from IGESSelect  inherits SelectExtract

    ---Purpose : This selections uses Subordinate Status as sort criterium
    --           It is an integer number which can be :
    --           0 Independant
    --           1 Physically Dependant
    --           2 Logically Dependant
    --           3 Both (recorded)
    --           + to sort :
    --           4 : 1 or 3  ->  at least Physically
    --           5 : 2 or 3  ->  at least Logically
    --           6 : 1 or 2 or 3 -> any kind of dependance
    --             (corresponds to 0 reversed)

uses AsciiString from TCollection, Transient, InterfaceModel
 
is
 
    Create (status : Integer) returns SelectSubordinate;
    ---Purpose : Creates a SelectSubordinate with a status to be sorted

    Status (me) returns Integer;
    ---Purpose : Returns the status used for sorting
 
    Sort (me; rank : Integer; ent : Transient; model : InterfaceModel)
        returns Boolean;
    ---Purpose : Returns True if <ent> is an IGES Entity with Subordinate
    --           Status matching the criterium

    ExtractLabel (me) returns AsciiString from TCollection;
    ---Purpose : Returns the Selection criterium : "IGES Entity, Independant"
    --           etc...

fields

    thestatus : Integer;

end SelectSubordinate;
