-- Created on: 2000-09-08
-- Created by: data exchange team
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Volume from XCAFDoc inherits Attribute from TDF

	---Purpose: 

uses
     Attribute       from TDF,
     Label           from TDF,
     GUID            from Standard,
     Real            from Standard,
     RelocationTable from TDF
    
is
    Create returns Volume from XCAFDoc;
    
    ---Purpose: class methods
    --          =============

    GetID (myclass) 
    	---C++: return const &  
    returns GUID from Standard;

    ID (me)
    	---C++: return const & 
    returns GUID from Standard;

    Set (me: mutable; vol: Real from Standard);
    	---Purpose: Sets a value of volume

    Set (myclass ; label : Label from TDF; vol: Real from Standard)
    returns Volume from XCAFDoc;
        ---Purpose: Find, or create, an Volume attribute and set its value

    Get (me)
    returns Real from Standard;
    
    Get (myclass ; label : Label from TDF; vol: in out Real from Standard)
    returns Boolean from Standard;
        ---Purpose: Returns volume as argument
	--          returns false if no such attribute at the <label>

    Restore (me: mutable; With : Attribute from TDF);

    NewEmpty(me)
    returns mutable Attribute from TDF;

    Paste (me; Into : mutable Attribute from TDF;
	       RT   : mutable RelocationTable from TDF);    

    Dump(me; anOS : in out OStream from Standard)
    returns OStream from Standard
    is redefined;
    ---C++: return &

fields

    myValue     : Real     from Standard;

end Volume from XCAFDoc;
