-- Created on: 2000-08-31
-- Created by: Andrey BETENEV
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class OperLibrary from ShapeProcess 

    ---Purpose: Provides a set of following operators
    --
    --          DirectFaces
    --          FixShape
    --          SameParameter
    --          SetTolerance
    --          SplitAngle
    --          BSplineRestriction
    --          ElementaryToRevolution
    --          SurfaceToBSpline
    --          ToBezier
    --          SplitContinuity
    --          SplitClosedFaces
    --          FixWireGaps
    --          FixFaceSize
    --          DropSmallEdges
    --          FixShape
    --          SplitClosedEdges

uses

    Shape               from TopoDS,
    UOperator           from ShapeProcess,
    ShapeContext        from ShapeProcess,
    Modification        from BRepTools,
    DataMapOfShapeShape from TopTools

is

    Init (myclass);
    	---Purpose: Registers all the operators

    ApplyModifier (myclass; S: Shape from TopoDS;
    	    	    	    context: ShapeContext from ShapeProcess;
			    M: Modification from BRepTools;
			    map: in out DataMapOfShapeShape from TopTools)
    	---Purpose: Applies BRepTools_Modification to a shape,
	--          taking into account sharing of components of compounds.
    returns Shape from TopoDS;

end OperLibrary;
