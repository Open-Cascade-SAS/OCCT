-- Created on: 1997-07-28
-- Created by: Pierre CHALAMET
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Modified :	GG 10/01/2000 IMP 
--		Add NumberOfTextures() and TextureName() methods
--		Add Name() method

class  TextureEnv  from  Graphic3d 
    
inherits  TextureRoot  from  Graphic3d 
 

    ---Purpose: This class provides environment texture usable only in Visual3d_ContextView

uses 
    NameOfTextureEnv  from  Graphic3d, 
    StructureManager  from  Graphic3d 

raises
    OutOfRange from Standard

is 
    Create(SM  :  StructureManager  from  Graphic3d; 
           aFileName  :  CString  from  Standard)
	returns  mutable TextureEnv  from  Graphic3d;    
    ---Purpose: Creates an environment texture from a file

    Create(SM  	:  StructureManager  from  Graphic3d;
    	   aName:  NameOfTextureEnv  from  Graphic3d)  
	returns  mutable  TextureEnv  from  Graphic3d; 
    ---Purpose: Creates an environment texture from a predefined texture name set.

    Name(me) returns NameOfTextureEnv from Graphic3d;
    ---Purpose:
    -- Returns the name of the predefined textures or NOT_ENV_UNKNOWN
    -- when the name is given as a filename.
    ---Level: Public

    NumberOfTextures(myclass) returns Integer from Standard;
    ---Purpose:
    -- Returns the number of predefined textures.
    ---Level: Public

    TextureName(myclass; aRank: Integer from Standard)
	returns CString from Standard
	raises OutOfRange from Standard;
    ---Purpose:
    -- Returns the name of the predefined texture of rank <aRank>
    ---Trigger: when <aRank> is < 1 or > NumberOfTextures.
    ---Level: Public

fields
    myName: NameOfTextureEnv from Graphic3d;
     
end  TextureEnv; 

