-- Created on: 1993-06-24
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class InterferenceTool from TopOpeBRepDS
     
uses

    Curve        from Geom2d,
    Orientation  from TopAbs,
    Transition   from TopOpeBRepDS,
    Interference from TopOpeBRepDS,
    Config       from TopOpeBRepDS,
    Kind         from TopOpeBRepDS
    
is

    MakeEdgeInterference(myclass;
			 T : Transition from TopOpeBRepDS;
	      	    	 SK : Kind; SI : Integer;
   	    	    	 GK : Kind; GI : Integer;
	      	    	 P : Real from Standard) 
    returns any Interference from TopOpeBRepDS;

    MakeCurveInterference(myclass;
    	     		  T : Transition from TopOpeBRepDS;
	      	    	  SK : Kind; SI : Integer;
    	    	    	  GK : Kind; GI : Integer;
	      	    	  P : Real from Standard) 
    returns any Interference from TopOpeBRepDS;

    DuplicateCurvePointInterference(myclass; I : Interference from TopOpeBRepDS)
    ---Purpose :  duplicate I in a new interference with Complement() transition.
    returns any Interference from TopOpeBRepDS;

    MakeFaceCurveInterference(myclass;
		    	      Transition : Transition from TopOpeBRepDS;
	      	    	      FaceI, CurveI : Integer from Standard;
	      	    	      PC : Curve from Geom2d) 
    returns any Interference from TopOpeBRepDS;

    MakeSolidSurfaceInterference(myclass;
    	      	    	    	 Transition : Transition from TopOpeBRepDS;
	      	    	    	 SolidI, SurfaceI : Integer from Standard)
    returns any Interference from TopOpeBRepDS;

    MakeEdgeVertexInterference(myclass;
    	      	    	       Transition : Transition from TopOpeBRepDS;
	      	    	       EdgeI, VertexI : Integer from Standard;
    	      	    	       VertexIsBound : Boolean from Standard;
    	      	    	       Config : Config from TopOpeBRepDS;
    	      	    	       param : Real from Standard)
    returns any Interference from TopOpeBRepDS;

    MakeFaceEdgeInterference(myclass;
    	      	    	       Transition : Transition from TopOpeBRepDS;
	      	    	       FaceI, EdgeI : Integer from Standard;
    	      	    	       EdgeIsBound : Boolean from Standard;
    	      	    	       Config : Config from TopOpeBRepDS)
    returns any Interference from TopOpeBRepDS;

    Parameter(myclass; CPI : Interference from TopOpeBRepDS)
    returns Real from Standard;

    Parameter(myclass; CPI : mutable Interference from TopOpeBRepDS; 
                       Par : Real from Standard);
    
end InterferenceTool from TopOpeBRepDS;
