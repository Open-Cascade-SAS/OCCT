-- Created on: 2000-05-10
-- Created by: Andrey BETENEV
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1

class ExternalSource from StepBasic
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity ExternalSource

uses
    SourceItem from StepBasic

is
    Create returns ExternalSource from StepBasic;
	---Purpose: Empty constructor

    Init (me: mutable; aSourceId: SourceItem from StepBasic);
	---Purpose: Initialize all fields (own and inherited)

    SourceId (me) returns SourceItem from StepBasic;
	---Purpose: Returns field SourceId
    SetSourceId (me: mutable; SourceId: SourceItem from StepBasic);
	---Purpose: Set field SourceId

fields
    theSourceId: SourceItem from StepBasic;

end ExternalSource;
