-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class FontSelect from StepVisual inherits SelectType from StepData

	-- <FontSelect> is an EXPRESS Select Type construct translation.
	-- it gathers : PreDefinedTextFont, ExternallyDefinedTextFont

uses

	PreDefinedTextFont,
	ExternallyDefinedTextFont
is

	Create returns FontSelect;
	---Purpose : Returns a FontSelect SelectType

	CaseNum (me; ent : Transient) returns Integer;
	---Purpose: Recognizes a FontSelect Kind Entity that is :
	--        1 -> PreDefinedTextFont
	--        2 -> ExternallyDefinedTextFont
	--        0 else

	PreDefinedTextFont (me) returns any PreDefinedTextFont;
	---Purpose : returns Value as a PreDefinedTextFont (Null if another type)

	ExternallyDefinedTextFont (me) returns any ExternallyDefinedTextFont;
	---Purpose : returns Value as a ExternallyDefinedTextFont (Null if another type)


end FontSelect;

