-- Created on: 1992-03-25
-- Created by: Isabelle GRIGNON
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Couple from IntSurf

	---Purpose: creation d 'un couple de 2 entiers

is

     Create
     	returns Couple from IntSurf;
     	---C++: inline

     Create(Index1, Index2 : Integer from Standard)
    	---C++: inline
    	returns Couple from IntSurf;
	
     
     First(me) returns Integer from Standard
     ---Purpose: returns the first element 
     ---C++: inline
     is static;


     Second (me) returns Integer from Standard
     ---Purpose: returns the Second element 
     ---C++: inline
     is static;


fields

    firstInteger  : Integer from Standard;
    secondInteger : Integer from Standard;

end Couple;


