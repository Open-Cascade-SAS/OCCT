-- Created on: 1997-02-28
-- Created by: Christophe LEYNADIER
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


private class TypedCallBack from Storage 

inherits TShared from MMgt

uses CallBack from Storage,
     AsciiString from TCollection
     
is
    Create returns mutable TypedCallBack from Storage;

    Create(aTypeName : AsciiString from TCollection; aCallBack : CallBack from Storage)
    	returns mutable TypedCallBack from Storage;

    SetType(me : mutable; aType : AsciiString from TCollection);
    Type(me) returns AsciiString from TCollection;
    
    SetCallBack(me : mutable; aCallBack : CallBack from Storage);
    CallBack(me) returns CallBack from Storage;

    SetIndex(me : mutable; anIndex : Integer from Standard);
    Index(me) returns Integer from Standard;
    
    fields
    
    	myType     : AsciiString from TCollection;
	myCallBack : CallBack from Storage;
    	myIndex    : Integer from Standard;
	
end;
