-- Created on: 1993-03-08
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Update:      Frederic Maupas


package PTopoDS 

	---Purpose: The package PTopoDS provides persistent classes to
	--          store Topological Data Structures in Data Base.
	--          
	--          The  structure  of  this  persistent  topology  is
	--          similar  to   the  transient  topology   (see  its
	--          documentation for more comprehension of this one).
	--          But some differences occure:
	--          
	--          * The class Model and derivatives disappear;
	--          
	--          * The "free"  information  disappears,  because  a 
	--          TShape stored in the Data Base is always "frozen";
	--          

	--          * The class HShape  inherits  from ExternShareable  from
	--          ObjMgt,  so that an intance of HShape  may be
	--          shared by a TShape even if the HShape is not in the
	--          same Container.
	--          
	--          * The class Shape1 inherits from Storable from
	--          Standard.
	--          
	--          Note that the  use of this topology is managed  by
	--          the package MgtTopoDS.
	--          
	--          About the question of "Location", see the  package
	--          PTopLoc  itself;  about  naming,  referencing  and
	--          using persistent  Shapes outsing  the  topological
	--          world, see the package TopoDB.

uses

    ObjMgt,
    Standard,
    TopAbs,      -- basic enumerations : ShapeEnum, Orientation
    PTopLoc,     -- Persistent local coordinate systems
    PCollection,
    TCollection
    
is

    ---Category: Old version of Shape/TShape.
    --           ============================

    class HShape;
	---Purpose: A reference (even outside the same container) to a
	--          Topological shape with Location, Orientation.
	
    deferred class TShape;
    	-- inherits ExternShareable from ObjMgt
	---Purpose: A topological shape is a structure made from other
	--          shapes.  This is a deferred class  used to support
	--          topological objects.
	
    deferred class TVertex;
	---Purpose: A TVertex  is a topological  point in two or three
	--          dimensions.
	
    class Vertex;
	---Purpose: A Vertex  is  a TVertex  with a  Location   and an
	--          Orientation.
	--          It inherits HShape
	
    deferred class TEdge;
	---Purpose: A topological part  of a  curve  in 2D or 3D,  the
	--          boundary    is   a   set  of oriented    Vertices.
	
    class Edge;
	---Purpose: A Edge  is a   TEdge    with  a Location  and   an
	--          Orientation.
	--          It inherits HShape
	
    class TWire;
	---Purpose: A set of Edges making a wire  structure, it can be
	--          a wireframe or a composite line.
	
    class Wire;
	---Purpose: A  Wire is  a   TWire  with  a  Location  and   an
	--          Orientation.
	--          It inherits HShape
	
    class TFace;
	---Purpose: A  topological part  of a  surface  or of  the  2D
	--          space. The boundary is a set of wires and edges.
	
    class Face;
	---Purpose: A Face  is   a   TFace with a   Location  and   an
	--          Orientation.
	--          It inherits HShape
	
    class TShell;
	---Purpose: A set of Faces or Shells, a topological surface or
	--          any faces structure.

    class Shell;
	---Purpose: A  Shell is a  TShell   with  a   Location  and an
	--          Orientation.
	--          It inherits HShape
	
    class TSolid;
	---Purpose: A Topological part of 3D  space, bounded by Shells
	--          and Faces.

    class Solid;
	---Purpose: A  Solid  is  a TSolid  with   a  Location and  an
	--          Orientation.
	--          It inherits HShape
	
    class TCompSolid;
	---Purpose: A structure of Solids sharing Faces.
	
    class CompSolid;
	---Purpose: A CompSolid is a TCompSolid with a Location and an
	--          Orientation.
	--          It inherits HShape
	
    class TCompound;
	---Purpose: A TCompound is an all-purpose set of Shapes.
	
    class Compound;
	---Purpose: A Compound is a  TCompound with a Location  and an
	--          Orientation.
	--          It inherits HShape
	

    class HArray1OfHShape instantiates HArray1 from PCollection
    	(HShape from PTopoDS);


    ---Category: New version of Shape/TShape.
    --           ============================

    class Shape1;
	---Purpose: A reference to a Topological TShape with Location,
	--          Orientation.
	
    deferred class TShape1;
    	-- inherits ExternShareable from ObjMgt
	---Purpose: A topological shape is a structure made from other
	--          shapes.  This is a deferred class  used to support
	--          topological objects.
	
    deferred class TVertex1;
	---Purpose: A TVertex  is a topological  point in two or three
	--          dimensions.
	
    deferred class TEdge1;
	---Purpose: A topological part  of a  curve  in 2D or 3D,  the
	--          boundary    is   a   set  of oriented    Vertices.
	
    class TWire1;
	---Purpose: A set of Edges making a wire  structure, it can be
	--          a wireframe or a composite line.
	
    class TFace1;
	---Purpose: A  topological part  of a  surface  or of  the  2D
	--          space. The boundary is a set of wires and edges.
	
    class TShell1;
	---Purpose: A set of Faces or Shells, a topological surface or
	--          any faces structure.

    class TSolid1;
	---Purpose: A Topological part of 3D  space, bounded by Shells
	--          and Faces.

    class TCompSolid1;
	---Purpose: A structure of Solids sharing Faces.
	
    class TCompound1;
	---Purpose: A TCompound is an all-purpose set of Shapes.
	

    class HArray1OfShape1 instantiates HArray1 from PCollection
    	(Shape1 from PTopoDS);

end PTopoDS;
