-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class CurveStyle from StepVisual 

inherits TShared from MMgt

uses

	HAsciiString from TCollection, 
	CurveStyleFontSelect from StepVisual, 
	SizeSelect from StepBasic, 
	Colour from StepVisual
is

	Create returns mutable CurveStyle;
	---Purpose: Returns a CurveStyle

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aCurveFont : CurveStyleFontSelect from StepVisual;
	      aCurveWidth : SizeSelect from StepBasic;
	      aCurveColour : mutable Colour from StepVisual) is virtual;

	-- Specific Methods for Field Data Access --

	SetName(me : mutable; aName : mutable HAsciiString);
	Name (me) returns mutable HAsciiString;
	SetCurveFont(me : mutable; aCurveFont : CurveStyleFontSelect);
	CurveFont (me) returns CurveStyleFontSelect;
	SetCurveWidth(me : mutable; aCurveWidth : SizeSelect);
	CurveWidth (me) returns SizeSelect;
	SetCurveColour(me : mutable; aCurveColour : mutable Colour);
	CurveColour (me) returns mutable Colour;

fields

	name : HAsciiString from TCollection;
	curveFont : CurveStyleFontSelect from StepVisual; -- a SelectType
	curveWidth : SizeSelect from StepBasic; -- a SelectType
	curveColour : Colour from StepVisual;

end CurveStyle;
