-- File:        ApprovalRole.cdl
-- Created:     Mon Dec  4 12:02:23 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWApprovalRole from RWStepBasic

	---Purpose : Read & Write Module for ApprovalRole

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     ApprovalRole from StepBasic

is

	Create returns RWApprovalRole;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable ApprovalRole from StepBasic);

	WriteStep (me; SW : in out StepWriter; ent : ApprovalRole from StepBasic);

end RWApprovalRole;
