-- Created on: 1994-05-27
-- Created by: Christian CAILLET
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



deferred class Transformer  from IFSelect  inherits TShared

    ---Purpose : A Transformer defines the way an InterfaceModel is transformed
    --           (without sending it to a file).
    --           In order to work, each type of Transformer defines it method
    --           Perform, it can be parametred as needed.
    --           
    --           It receives a Model (the data set) as input. It then can :
    --           - edit this Model on the spot (i.e. alter its content : by
    --             editing entities, or adding/replacing some ...)
    --           - produce a copied Model, which detains the needed changes
    --             (typically on the same type, but some or all entities beeing
    --              rebuilt or converted; or converted from a protocol to
    --              another one)

uses AsciiString from TCollection,
     CheckIterator, Graph, Protocol from Interface, InterfaceModel

is

    Perform (me : mutable; G : Graph; protocol : Protocol from Interface;
    	     checks : in out CheckIterator;
    	     newmod : out mutable InterfaceModel)  returns Boolean  is deferred;
    ---Purpose : Performs a Transformation (defined by each sub-class) :
    --         <G> gives the input data (especially the starting model) and
    --           can be used for queries (by Selections, etc...)
    --         <protocol> allows to work with General Services as necessary
    --           (it applies to input data)
    --           If the change corresponds to a conversion to a new protocol,
    --           see also the method ChangeProtocol
    --         <checks> stores produced checks messages if any
    --         <newmod> gives the result of the transformation :
    --         - if it is Null (i.e. has not been affected), the transformation
    --           has been made on the spot, it is assumed to cause no change
    --           to the graph of dependances
    --         - if it equates the starting Model, it has been transformed on
    --           the spot (possibiliy some entities were replaced inside it)
    --         - if it is new, it corresponds to a new data set which replaces
    --           the starting one
    --         
    --         <me> is mutable to allow results for ChangeProtocol to be
    --           memorized if needed, and to store informations useful for
    --           the method Updated
    --         
    --         Returns True if Done, False if an Error occured : in this case,
    --           if a new data set has been produced, the transformation
    --           is ignored, else data may be corrupted.

    ChangeProtocol (me; newproto : in out Protocol from Interface)
    	returns Boolean  is virtual;
    ---Purpose : This methods allows to declare that the Protocol applied to
    --           the new Model has changed. It applies to the last call to
    --           Perform.
    --           
    --           Returns True if the Protocol has changed, False else.
    --           The provided default keeps the starting Protocol. This method
    --           should be redefined as required by the effect of Perform.

    Updated (me; entfrom : Transient; entto : out mutable Transient)
    	returns Boolean  is deferred;
    ---Purpose : This method allows to know what happened to a starting
    --           entity after the last Perform. If <entfrom> (from starting
    --           model) has one and only one known item which corresponds in
    --           the new produced model, this method must return True and
    --           fill the argument <entto>. Else, it returns False.

    Label (me) returns AsciiString from TCollection  is deferred;
    ---Purpose : Returns a text which defines the way a Transformer works
    --           (to identify the transformation it performs)

end Transformer;
