-- Created on: 1993-05-06
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class Polygo from IntPatch

	---Purpose: 

inherits Polygon2d from Intf

uses Pnt2d from gp,
     Box2d from Bnd

raises OutOfRange from Standard

is

    Initialize (theError : Real from Standard = 0.0)
        returns Polygo from IntPatch;

    Error (me) returns Real from Standard;
    ---C++: inline

    NbPoints (me) returns Integer is deferred;

    Point (me; Index : Integer) returns Pnt2d from gp is deferred;

    DeflectionOverEstimation (me)
    returns Real from Standard is redefined virtual;
    ---C++: inline
    ---Purpose: Returns the tolerance of the polygon.

    NbSegments (me)
    returns Integer from Standard is redefined virtual;
    ---C++: inline
    ---Purpose: Returns the number of Segments in the polyline.

    Segment (me; theIndex : in Integer from Standard;
                 theBegin, theEnd : in out Pnt2d from gp)
        raises OutOfRange from Standard is redefined virtual;
    ---C++: inline
    ---Purpose: Returns the points of the segment <Index> in the Polygon.

    Dump (me);

fields

    myError : Real from Standard is protected;

end Polygo;
