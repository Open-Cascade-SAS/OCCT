-- Created on: 1992-06-04
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class CurveTool from Geom2dGcc

	---Purpose: 

uses Curve from Geom2dAdaptor,
     Pnt2d from gp,
     Vec2d from gp

is

    FirstParameter(myclass; C: Curve from Geom2dAdaptor)
    	returns Real;

    LastParameter(myclass; C: Curve from Geom2dAdaptor)
    	returns Real;

    EpsX (myclass                           ; 
    	  C       : Curve from Geom2dAdaptor;
    	  Tol     : Real  from Standard     )
    	returns Real;

    NbSamples(myclass                    ;
    	      C       : Curve from Geom2dAdaptor)
    	returns Integer;

    Value (myclass; C: Curve from Geom2dAdaptor; X: Real)
    	returns Pnt2d from gp;

    D1 (myclass; C: Curve from Geom2dAdaptor; U: Real ; 
                 P: out Pnt2d; T: out Vec2d);

    D2 (myclass; C: Curve from Geom2dAdaptor; U: Real ; 
                 P: out Pnt2d; T,N: out Vec2d);

    D3 (myclass; C: Curve from Geom2dAdaptor; U: Real ; 
                 P: out Pnt2d; T,N,dN: out Vec2d);

end CurveTool;

