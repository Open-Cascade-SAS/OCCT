-- Created on: 1999-07-12
-- Created by: Denis PASCAL
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




private class Owner from TDocStd inherits Attribute from TDF

	---Purpose: 

uses Attribute from TDF,
     GUID      from Standard, 
     RelocationTable from TDF, 
     Data      from TDF,
     Label     from TDF,
     Document  from TDocStd

is 

    ---Purpose: class methods
    --          =============

    GetID (myclass)   
    	---C++: return const &  
    returns GUID from Standard;

    SetDocument (myclass; indata : Data from TDF; doc : Document from TDocStd);
    
    GetDocument (myclass; ofdata : Data from TDF)
    returns Document from TDocStd;

    ---Purpose: Owner methods
    --          ===============
    
    Create
    returns mutable Owner from TDocStd;  
    
    SetDocument (me : mutable; document : Document from TDocStd);    

    GetDocument (me)
    returns Document from TDocStd;
    
    ---Category: methodes de TDF_Attribute
    --           =========================
    
    ID (me)
    	---C++: return const & 
    returns GUID from Standard;

    Restore (me: mutable; With : Attribute from TDF);

    NewEmpty (me)
    returns mutable Attribute from TDF;

    Paste (me; Into : mutable Attribute from TDF;
	       RT   : mutable RelocationTable from TDF);    

    Dump(me; anOS : in out OStream from Standard)
    	returns OStream from Standard
    	is redefined;
	---C++: return &

fields

    myDocument : Document from TDocStd;

end Owner;
