-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ShapeAspect from StepRepr 

inherits TShared from MMgt

uses

	HAsciiString from TCollection, 
	ProductDefinitionShape from StepRepr, 
	Logical from StepData
is

	Create returns mutable ShapeAspect;
	---Purpose: Returns a ShapeAspect

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aDescription : mutable HAsciiString from TCollection;
	      aOfShape : mutable ProductDefinitionShape from StepRepr;
	      aProductDefinitional : Logical from StepData) is virtual;

	-- Specific Methods for Field Data Access --

	SetName(me : mutable; aName : mutable HAsciiString);
	Name (me) returns mutable HAsciiString;
	SetDescription(me : mutable; aDescription : mutable HAsciiString);
	Description (me) returns mutable HAsciiString;
	SetOfShape(me : mutable; aOfShape : mutable ProductDefinitionShape);
	OfShape (me) returns mutable ProductDefinitionShape;
	SetProductDefinitional(me : mutable; aProductDefinitional : Logical);
	ProductDefinitional (me) returns Logical;

fields

	name : HAsciiString from TCollection;
	description : HAsciiString from TCollection;
	ofShape : ProductDefinitionShape from StepRepr;
	productDefinitional : Logical from StepData;

end ShapeAspect;
