-- File:        PlanarExtent.cdl
-- Created:     Fri Dec  1 11:11:24 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class PlanarExtent from StepVisual 

inherits GeometricRepresentationItem from StepGeom

uses

	Real from Standard, 
	HAsciiString from TCollection
is

	Create returns mutable PlanarExtent;
	---Purpose: Returns a PlanarExtent


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aSizeInX : Real from Standard;
	      aSizeInY : Real from Standard) is virtual;

	-- Specific Methods for Field Data Access --

	SetSizeInX(me : mutable; aSizeInX : Real);
	SizeInX (me) returns Real;
	SetSizeInY(me : mutable; aSizeInY : Real);
	SizeInY (me) returns Real;

fields

	sizeInX : Real from Standard;
	sizeInY : Real from Standard;

end PlanarExtent;
