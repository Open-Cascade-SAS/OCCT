-- File:	STEPCAFControl_ActorWrite.cdl
-- Created:	Thu Oct  5 19:34:41 2000
-- Author:	Andrey BETENEV
--		<abv@doomox.nnov.matra-dtv.fr>
---Copyright:	 Matra Datavision 2000


class ActorWrite from STEPCAFControl inherits ActorWrite from STEPControl

    ---Purpose: Extends ActorWrite from STEPControl by analysis of
    --          whether shape is assembly (based on information from DECAF)

uses
    Shape from TopoDS,
    MapOfShape from TopTools

is

    Create returns mutable ActorWrite;

    IsAssembly (me; S: in out Shape from TopoDS) returns Boolean is redefined;
    	---Purpose: Check whether shape S is assembly
	--          Returns True if shape is registered in assemblies map

    SetStdMode (me: mutable; stdmode: Boolean = Standard_True);
    	---Purpose: Set standard mode of work 
	--          In standard mode Actor (default) behaves exactly as its 
        --          ancestor, also map is cleared

    ClearMap (me: mutable);
    	---Purpose: Clears map of shapes registered as assemblies

    RegisterAssembly (me: mutable; S: Shape from TopoDS);
    	---Purpose: Registers shape to be written as assembly
	--          The shape should be TopoDS_Compound (else does nothing)

fields

    myStdMode: Boolean;
    myMap: MapOfShape from TopTools;

end ActorWrite;
