-- Created on: 1993-07-12
-- Created by: Yves FRICAUD
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class SketchExplorer from MAT2d

	---Purpose: SketchExplorer  is  an iterator on  a  sketch.   A
	--          sketch is a set of contours, each contour is a set
	--          of curves from Geom2d.

uses

    Curve           from Geom2d
is
    
    NumberOfContours(me)
	--- Purpose : Returns the number of contours in the figure.
    returns Integer;
       
    Init(me : in out ; ContourIndex : Integer );
	--- Purpose : Initializes the curves explorer on the contour
	--            of range <ContourIndex>.           
   
    More(me) returns Boolean from Standard;
       	--- Purpose: Returns False if  there is no  more curves on the
       	--           current contour.
    
    Next(me : in out);
	--- Purpose  : Moves to the next curve of the current contour.
    
    Value(me) returns Curve from Geom2d; 
        --- Purpose : Returns the current curve on the current contour.
    

end SketchExplorer;




