-- Created on: 1995-02-08
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class LineTool from GeomInt

	---Purpose: 

uses Line  from IntPatch,
     Point from IntPatch,
     Pnt2d from gp

is


    NbVertex(myclass; L: Line from IntPatch)
    
    	returns Integer from Standard;


    Vertex(myclass; L:Line from IntPatch; I: Integer from Standard)
    
    	returns Point from IntPatch;
	---C++: return const&
	
    FirstParameter(myclass; L: Line from IntPatch)
    
    	returns Real from Standard;


    LastParameter(myclass; L: Line from IntPatch)
    
    	returns Real from Standard;


end LineTool;
