-- File:        Representation.cdl
-- Created:     Mon Dec  4 12:02:31 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWRepresentation from RWStepRepr

	---Purpose : Read & Write Module for Representation

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     Representation from StepRepr,
     EntityIterator from Interface

is

	Create returns RWRepresentation;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable Representation from StepRepr);

	WriteStep (me; SW : in out StepWriter; ent : Representation from StepRepr);

	Share(me; ent : Representation from StepRepr; iter : in out EntityIterator);

end RWRepresentation;
