-- File:	MXCAFDoc_LocationRetrievalDriver.cdl
-- Created:	Tue Aug 15 15:16:37 2000
-- Author:	data exchange team
--		<det@strelox.nnov.matra-dtv.fr>
---Copyright:	 Matra Datavision 2000


class LocationRetrievalDriver from MXCAFDoc inherits ARDriver from MDF

	---Purpose: 

uses
    RRelocationTable from MDF,
    Attribute        from PDF,
    Attribute        from TDF,
    MessageDriver    from CDM

is
--    Create -- Version 0
--    returns mutable LocationRetrievalDriver from MXCAFDoc;
    Create (theMsgDriver : MessageDriver from CDM)
    returns mutable LocationRetrievalDriver from MXCAFDoc;
    
    VersionNumber(me) returns Integer from Standard;
    ---Purpose: Returns the version number from which the driver
    --          is available: 0.

    SourceType(me) returns Type from Standard;
    ---Purpose: Returns the type: XCAFDoc_Location

    NewEmpty (me)  returns mutable Attribute from TDF;

    Paste(me;
    	  Source     :         Attribute from PDF;
    	  Target     : mutable Attribute from TDF;
    	  RelocTable : RRelocationTable from MDF);

end LocationRetrievalDriver;

    
