-- Created on: 1999-06-22
-- Created by: data exchange team
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ApplySequence from ShapeProcessAPI 

    ---Purpose: Applies one of the sequence read from resource file.

uses
    
    ShapeEnum           from TopAbs,
    Shape               from TopoDS,
    DataMapOfShapeShape from TopTools,
    Printer             from Message,
    ShapeContext        from ShapeProcess,
    AsciiString         from TCollection
is

    Create (rscName: CString; seqName: CString = "") returns ApplySequence from ShapeProcessAPI;
    	---Purpose: Creates an object and loads resource file and sequence of
    	--          operators given by their names.
    
    Context (me: in out) returns ShapeContext from ShapeProcess;
    	---C++ : return &
	---Purpose: Returns object for managing resource file and sequence of
    	--          operators.
    
    PrepareShape (me: in out; shape  : Shape from TopoDS;
    	    	    	      fillmap: Boolean = Standard_False;
			      until  : ShapeEnum from TopAbs = TopAbs_SHAPE)
    returns Shape from TopoDS;
    	---Purpose: Performs sequence of operators stored in myRsc.
	--          If <fillmap> is True adds history "shape-shape" into myMap
	--          for shape and its subshapes until level <until> (included).
    	--          If <until> is TopAbs_SHAPE,  all the subshapes are considered.
	
    ClearMap (me: in out);
    	---Purpose: Clears myMap with accumulated history.
	
    Map (me) returns DataMapOfShapeShape from TopTools;
    	---C++: return const &
	---Purpose: Returns myMap with accumulated history.

    PrintPreparationResult (me);
    	---Purpose: Prints result of preparation onto the messenger of the context.
	--          Note that results can be accumulated from previous preparations
	--          it method ClearMap was not called before PrepareShape.
	---Remark: At the moment outputs information only on shells and faces.
    
fields

    myContext: ShapeContext from ShapeProcess;
    myMap    : DataMapOfShapeShape from TopTools;
    mySeq    : AsciiString from TCollection;

end ApplySequence;
