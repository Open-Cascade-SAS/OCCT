-- Created on: 1993-03-09
-- Created by: JCV
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class BSplineSurface from Geom inherits BoundedSurface from Geom

        ---Purpose : Describes a BSpline surface.
    	-- In each parametric direction, a BSpline surface can be:
    	-- - uniform or non-uniform,
    	-- - rational or non-rational,
    	-- - periodic or non-periodic.
    	-- A BSpline surface is defined by:
    	-- - its degrees, in the u and v parametric directions,
    	-- - its periodic characteristic, in the u and v parametric directions,
    	-- - a table of poles, also called control points (together
    	--   with the associated weights if the surface is rational), and
    	-- - a table of knots, together with the associated multiplicities.
    	--   The degree of a Geom_BSplineSurface is limited to
    	-- a value (25) which is defined and controlled by the
    	-- system. This value is returned by the function MaxDegree.
    	--       Poles and Weights
    	-- Poles and Weights are manipulated using two associative double arrays:
    	-- - the poles table, which is a double array of gp_Pnt points, and
    	-- - the weights table, which is a double array of reals.
    	-- The bounds of the poles and weights arrays are:
    	-- - 1 and NbUPoles for the row bounds (provided
    	--   that the BSpline surface is not periodic in the u
    	--   parametric direction), where NbUPoles is the
    	--   number of poles of the surface in the u parametric direction, and
    	-- - 1 and NbVPoles for the column bounds (provided
    	--   that the BSpline surface is not periodic in the v
    	--   parametric direction), where NbVPoles is the
    	--   number of poles of the surface in the v parametric direction.
    	--   The poles of the surface are the points used to shape
    	-- and reshape the surface. They comprise a rectangular network.
    	-- If the surface is not periodic:
    	-- - The points (1, 1), (NbUPoles, 1), (1,
    	--   NbVPoles), and (NbUPoles, NbVPoles)
    	--   are the four parametric "corners" of the surface.
    	-- - The first column of poles and the last column of
    	--   poles define two BSpline curves which delimit the
    	--   surface in the v parametric direction. These are the
    	--   v isoparametric curves corresponding to the two
    	--   bounds of the v parameter.
    	-- - The first row of poles and the last row of poles
    	--   define two BSpline curves which delimit the surface
    	--   in the u parametric direction. These are the u
    	--   isoparametric curves corresponding to the two bounds of the u parameter.
    	-- If the surface is periodic, these geometric properties are not verified.
    	-- It is more difficult to define a geometrical significance
    	-- for the weights. However they are useful for
    	-- representing a quadric surface precisely. Moreover, if
    	-- the weights of all the poles are equal, the surface has
    	-- a polynomial equation, and hence is a "non-rational surface".
    	-- The non-rational surface is a special, but frequently
    	-- used, case, where all poles have identical weights.
    	-- The weights are defined and used only in the case of
    	-- a rational surface. The rational characteristic is
    	-- defined in each parametric direction. A surface can be
    	-- rational in the u parametric direction, and
    	-- non-rational in the v parametric direction.
    	--        Knots and Multiplicities
    	-- For a Geom_BSplineSurface the table of knots is
    	-- made up of two increasing sequences of reals, without
    	-- repetition, one for each parametric direction. The
    	-- multiplicities define the repetition of the knots.
    	-- A BSpline surface comprises multiple contiguous
    	-- patches, which are themselves polynomial or rational
    	-- surfaces. The knots are the parameters of the
    	-- isoparametric curves which limit these contiguous
    	-- patches. The multiplicity of a knot on a BSpline
    	-- surface (in a given parametric direction) is related to
    	-- the degree of continuity of the surface at that knot in
    	-- that parametric direction:
    	-- Degree of continuity at knot(i) = Degree - Multi(i) where:
    	-- - Degree is the degree of the BSpline surface in
    	--   the given parametric direction, and
    	-- - Multi(i) is the multiplicity of knot number i in
    	--   the given parametric direction.
    	-- There are some special cases, where the knots are
    	-- regularly spaced in one parametric direction (i.e. the
    	-- difference between two consecutive knots is a constant).
    	-- - "Uniform": all the multiplicities are equal to 1.
    	-- - "Quasi-uniform": all the multiplicities are equal to 1,
    	--   except for the first and last knots in this parametric
    	--   direction, and these are equal to Degree + 1.
    	-- - "Piecewise Bezier": all the multiplicities are equal to
    	--   Degree except for the first and last knots, which
    	--   are equal to Degree + 1. This surface is a
    	--   concatenation of Bezier patches in the given
    	--   parametric direction.
    	-- If the BSpline surface is not periodic in a given
    	-- parametric direction, the bounds of the knots and
    	-- multiplicities tables are 1 and NbKnots, where
    	-- NbKnots is the number of knots of the BSpline
    	-- surface in that parametric direction.
    	-- If the BSpline surface is periodic in a given parametric
    	-- direction, and there are k periodic knots and p
    	-- periodic poles in that parametric direction:
    	-- - the period is such that:
    	-- period = Knot(k+1) - Knot(1), and
    	-- - the poles and knots tables in that parametric
    	--   direction can be considered as infinite tables, such that:
    	-- Knot(i+k) = Knot(i) + period, and
    	-- Pole(i+p) = Pole(i)
    	-- Note: The data structure tables for a periodic BSpline
    	-- surface are more complex than those of a non-periodic one.
        -- References :
        --  . A survey of curve and surface methods in CADG Wolfgang BOHM
        --    CAGD 1 (1984)
        --  . On de Boor-like algorithms and blossoming Wolfgang BOEHM
        --    cagd 5 (1988)
        --  . Blossoming and knot insertion algorithms for B-spline curves
        --    Ronald N. GOLDMAN
        --  . Modelisation des surfaces en CAO, Henri GIAUME Peugeot SA   
        --  . Curves and Surfaces for Computer Aided Geometric Design,
        --    a practical guide Gerald Farin



uses  Array1OfInteger      from TColStd,
      Array1OfReal         from TColStd,
      Array2OfReal         from TColStd, 
      HArray1OfInteger     from TColStd,
      HArray1OfReal        from TColStd,
      HArray2OfReal        from TColStd,
      Array1OfPnt          from TColgp, 
      Array2OfPnt          from TColgp,
      Ax1                  from gp, 
      Ax2                  from gp,
      HArray2OfPnt         from TColgp, 
      Pnt                  from gp,
      Trsf                 from gp,
      Vec                  from gp, 
      BSplKnotDistribution from GeomAbs,
      Curve                from Geom,
      Geometry             from Geom,
      Shape                from GeomAbs,
      Mutex                from Standard

raises ConstructionError   from Standard,
       DimensionError      from Standard,
       DomainError         from Standard,
       OutOfRange          from Standard,
       NoSuchObject        from Standard,
       RangeError          from Standard,
       UndefinedDerivative from Geom



is
      


  Create (Poles                        : Array2OfPnt     from TColgp; 
          UKnots, VKnots               : Array1OfReal    from TColStd; 
          UMults, VMults               : Array1OfInteger from TColStd; 
          UDegree, VDegree             : Integer;
    	  UPeriodic                    : Boolean = Standard_False;
    	  VPeriodic                    : Boolean = Standard_False)
     returns BSplineSurface
     
    	---Purpose : Creates  a non-rational b-spline surface (weights
        --         default value is 1.).
     raises ConstructionError;
    	---Purpose: The following conditions must be verified.
    	--   0 < UDegree <= MaxDegree.
        --   UKnots.Length() == UMults.Length() >= 2
        --   UKnots(i) < UKnots(i+1) (Knots are increasing)
        --   1 <= UMults(i) <= UDegree
    	--   On a   non  uperiodic   surface    the  first and    last 
    	--   umultiplicities  may  be     UDegree+1  (this   is   even
    	--   recommanded if you want the curve  to start and finish on
        --   the first and last pole).
    	--   On a uperiodic     surface  the first    and   the   last
        --   umultiplicities must be the same.
        --   on non-uperiodic surfaces
    	--     Poles.ColLength() == Sum(UMults(i)) - UDegree - 1 >= 2
        --   on uperiodic surfaces 
    	--   Poles.ColLength() == Sum(UMults(i)) except the first or last
    	--   The previous conditions for U holds  also for V, with the
        --   RowLength of the poles.




  Create (Poles                        : Array2OfPnt     from TColgp; 
    	  Weights                      : Array2OfReal    from TColStd;
          UKnots, VKnots               : Array1OfReal    from TColStd; 
          UMults, VMults               : Array1OfInteger from TColStd; 
          UDegree, VDegree             : Integer;
    	  UPeriodic                    : Boolean = Standard_False;
    	  VPeriodic                    : Boolean = Standard_False)
     returns BSplineSurface
     
        ---Purpose : Creates  a non-rational b-spline surface (weights
        --         default value is 1.).
        --  
     raises ConstructionError;
    	---Purpose: The following conditions must be verified.
        --  0 < UDegree <= MaxDegree.
        --  
        --  UKnots.Length() == UMults.Length() >= 2
        --  
        --  UKnots(i) < UKnots(i+1) (Knots are increasing)
        --  1 <= UMults(i) <= UDegree
        --  
        --   On a   non  uperiodic   surface    the  first and    last
        --   umultiplicities  may  be     UDegree+1  (this   is   even
        --   recommanded if you want the curve  to start and finish on
        --   the first and last pole).
        --   
        --   On a uperiodic     surface  the first    and   the   last
        --   umultiplicities must be the same.
        --   
        --   on non-uperiodic surfaces
        --   
        --     Poles.ColLength() == Sum(UMults(i)) - UDegree - 1 >= 2
        --     
        --   on uperiodic surfaces 
        --   
        --     Poles.ColLength() == Sum(UMults(i)) except the first or
        --     last
        --     
        --   
        --   The previous conditions for U holds  also for V, with the
        --   RowLength of the poles.



  ExchangeUV (me : mutable);
    	---Purpose: Exchanges the u and v parametric directions on
    	-- this BSpline surface.
    	-- As a consequence:
    	-- - the poles and weights tables are transposed,
    	-- - the knots and multiplicities tables are exchanged,
    	-- - degrees of continuity, and rational, periodic and
    	--   uniform characteristics are exchanged, and
    	-- - the orientation of the surface is inverted.

  SetUPeriodic (me : mutable);
	---Purpose: Sets the surface U periodic.

  SetVPeriodic (me : mutable);
	---Purpose:  Modifies this surface to be periodic in the u (or v)
    	-- parametric direction.
    	-- To become periodic in a given parametric direction a
    	-- surface must be closed in that parametric direction,
    	-- and the knot sequence relative to that direction must be periodic.
    	-- To generate this periodic sequence of knots, the
    	-- functions FirstUKnotIndex and LastUKnotIndex (or
    	-- FirstVKnotIndex and LastVKnotIndex) are used to
    	-- compute I1 and I2. These are the indexes, in the
    	-- knot array associated with the given parametric
    	-- direction, of the knots that correspond to the first and
    	-- last parameters of this BSpline surface in the given
    	-- parametric direction. Hence the period is:
    	-- Knots(I1) - Knots(I2)
    	-- As a result, the knots and poles tables are modified.
    	-- Exceptions
    	-- Standard_ConstructionError if the surface is not
    	-- closed in the given parametric direction.
	         
	      
	     
        
  PeriodicNormalization(me ;  U,V : in out Real) ; 
       
        ---Purpose : returns the parameter normalized within
        --         the period if the surface is periodic : otherwise
        --         does not do anything

  SetUOrigin (me : mutable; Index : Integer)
    	---Purpose: Assigns the knot of index Index in the knots table in
    	-- the corresponding parametric direction to be the
    	-- origin of this periodic BSpline surface. As a
    	-- consequence, the knots and poles tables are modified.
    	-- Exceptions
    	-- Standard_NoSuchObject if this BSpline surface is
    	-- not periodic in the given parametric direction.
    	-- Standard_DomainError if Index is outside the
    	-- bounds of the knots table in the given parametric direction.
    raises NoSuchObject,
    	   DomainError;
	
  SetVOrigin (me : mutable; Index : Integer)
    	---Purpose: Assigns the knot of index Index in the knots table in
    	-- the corresponding parametric direction to be the
    	-- origin of this periodic BSpline surface. As a
    	-- consequence, the knots and poles tables are modified.
    	-- Exceptions
    	-- Standard_NoSuchObject if this BSpline surface is
    	-- not periodic in the given parametric direction.
    	-- Standard_DomainError if Index is outside the
    	-- bounds of the knots table in the given parametric direction.
    raises NoSuchObject,
    	   DomainError;
	

  SetUNotPeriodic (me : mutable);

  SetVNotPeriodic (me : mutable);
    	---Purpose: Modifies this surface to be periodic in the u (or v) parametric direction.
    	-- To become periodic in a given parametric direction a
    	-- surface must be closed in that parametric direction,
    	-- and the knot sequence relative to that direction must be periodic.
    	-- To generate this periodic sequence of knots, the
    	-- functions FirstUKnotIndex and LastUKnotIndex (or
    	-- FirstVKnotIndex and LastVKnotIndex) are used to
    	-- compute I1 and I2. These are the indexes, in the
    	-- knot array associated with the given parametric
    	-- direction, of the knots that correspond to the first and
    	-- last parameters of this BSpline surface in the given
    	-- parametric direction. Hence the period is:
    	-- Knots(I1) - Knots(I2)
    	-- As a result, the knots and poles tables are modified.
    	-- Exceptions
    	-- Standard_ConstructionError if the surface is not
    	-- closed in the given parametric direction.

  UReverse (me : mutable);
    
  VReverse (me : mutable);
        ---Purpose: Changes the orientation of this BSpline surface in the
    	-- u (or v) parametric direction. The bounds of the
    	-- surface are not changed but the given parametric
    	-- direction is reversed. Hence the orientation of the
    	-- surface is reversed.
    	-- The knots and poles tables are modified.
    
  UReversedParameter (me; U : Real) returns Real;
  
  VReversedParameter (me; V : Real) returns Real;
	---Purpose: Computes the u (or v) parameter on the modified
    	-- surface, produced by reversing its u (or v) parametric
    	-- direction, for the point of u parameter U, (or of v
    	-- parameter V) on this BSpline surface.
    	-- For a BSpline surface, these functions return respectively:
    	-- - UFirst + ULast - U, or
    	-- - VFirst + VLast - V,
    	-- where UFirst, ULast, VFirst and VLast are
    	-- the values of the first and last parameters of this
    	-- BSpline surface, in the u and v parametric directions.


  IncreaseDegree (me : mutable; UDegree, VDegree : Integer);
    	---Purpose : Increases the degrees of this BSpline surface to
    	-- UDegree and VDegree in the u and v parametric
    	-- directions respectively. As a result, the tables of poles,
    	-- weights and multiplicities are modified. The tables of
    	-- knots is not changed.
    	-- Note: Nothing is done if the given degree is less than
    	-- or equal to the current degree in the corresponding
    	-- parametric direction.
    	-- Exceptions
    	-- Standard_ConstructionError if UDegree or
    	-- VDegree is greater than
    	-- Geom_BSplineSurface::MaxDegree().


  InsertUKnots (me : mutable; Knots : Array1OfReal    from TColStd; 
    	    	    	      Mults : Array1OfInteger from TColStd;
    	    	    	      ParametricTolerance : Real = 0.0;
    	    	    	      Add : Boolean = Standard_True);
			     
  InsertVKnots (me : mutable; Knots : Array1OfReal    from TColStd; 
    	    	    	      Mults : Array1OfInteger from TColStd;
    	    	    	      ParametricTolerance : Real = 0.0;
    	    	    	      Add : Boolean = Standard_True);
			     
        ---Purpose: Inserts into the knots table for the corresponding
    	-- parametric direction of this BSpline surface:
    	-- - the value U, or V, with the multiplicity M (defaulted to 1), or
    	-- - the values of the array Knots, with their respective
    	-- multiplicities, Mults.
    	-- If the knot value to insert already exists in the table, its multiplicity is:
    	-- - increased by M, if Add is true (the default), or
    	-- - increased to M, if Add is false.
    	-- The tolerance criterion used to check the equality of
    	-- the knots is the larger of the values ParametricTolerance and
	-- Standard_Real::Epsilon(val), where val is the knot value to be inserted.
    	-- Warning
    	-- - If a given multiplicity coefficient is null, or negative, nothing is done.
    	-- - The new multiplicity of a knot is limited to the degree of this BSpline surface in the
    	--   corresponding parametric direction.
    	-- Exceptions
    	-- Standard_ConstructionError if a knot value to
    	-- insert is outside the bounds of this BSpline surface in
    	-- the specified parametric direction. The comparison
    	-- uses the precision criterion ParametricTolerance.
   
     
  RemoveUKnot(me : mutable; Index     : Integer; 
    	    	    	   M         : Integer;
    	    	    	   Tolerance : Real) returns Boolean
  raises OutOfRange;
			   
  RemoveVKnot(me : mutable; Index     : Integer; 
    	    	    	   M         : Integer;
    	    	    	   Tolerance : Real) returns Boolean
  raises OutOfRange;
			   
        ---Purpose : Reduces to M the multiplicity of the knot of index
    	-- Index in the given parametric direction. If M is 0, the knot is removed.
    	-- With a modification of this type, the table of poles is also modified.
    	-- Two different algorithms are used systematically to
    	-- compute the new poles of the surface. For each
    	-- pole, the distance between the pole calculated
    	-- using the first algorithm and the same pole
    	-- calculated using the second algorithm, is checked. If
    	-- this distance is less than Tolerance it ensures that
    	-- the surface is not modified by more than Tolerance.
    	-- Under these conditions, the function returns true;
    	-- otherwise, it returns false.
    	-- A low tolerance prevents modification of the
    	-- surface. A high tolerance "smoothes" the surface.
    	-- Exceptions
    	-- Standard_OutOfRange if Index is outside the
    	-- bounds of the knots table of this BSpline surface.         

     
  IncreaseUMultiplicity (me : mutable; UIndex : Integer; M : Integer)
        ---Purpose :
        --  Increases the multiplicity of the knot of range UIndex 
        --  in the UKnots sequence.
        --  M is the new multiplicity. M must be greater than the
        --  previous multiplicity and lower or equal to the degree
        --  of the surface in the U parametric direction.
     raises ConstructionError,
        ---Purpose : Raised if M is not in the range [1, UDegree]
            OutOfRange;
        ---Purpose : 
        --  Raised if UIndex is not in the range [FirstUKnotIndex,
        --  LastUKnotIndex] given by the methods with the same name.


  IncreaseUMultiplicity (me : mutable; FromI1, ToI2 : Integer; M : Integer)
        ---Purpose :
        --  Increases until order M the multiplicity of the set of knots
        --  FromI1,...., ToI2 in the U direction. This method can be used 
        --  to make a B_spline surface into a PiecewiseBezier B_spline
        --  surface.
        --  If <me> was uniform, it can become non uniform.
     raises OutOfRange,
        ---Purpose :
        --  Raised if FromI1 or ToI2 is out of the range [FirstUKnotIndex,
        --  LastUKnotIndex].
            ConstructionError;
        ---Purpose : 
        --  M should be greater than the previous multiplicity of the 
        --  all the knots FromI1,..., ToI2 and lower or equal to the
        --   Degree of the surface in the U parametric direction.


  IncrementUMultiplicity (me : mutable; FromI1, ToI2 : Integer; Step : Integer)
        ---Purpose :
        --  Increments the multiplicity of the consecutives uknots FromI1..ToI2
        --  by step.   The multiplicity of each knot FromI1,.....,ToI2 must be
        --  lower or equal to the UDegree of the B_spline.
     raises OutOfRange,
        ---Purpose :
        --  Raised if FromI1 or ToI2 is not in the range
        --  [FirstUKnotIndex, LastUKnotIndex] 
            ConstructionError;
       ---Purpose :
        --  Raised if one knot has a multiplicity greater than UDegree.


  IncreaseVMultiplicity (me : mutable; VIndex : Integer; M : Integer)
        ---Purpose :
        --  Increases the multiplicity of a knot in the V direction.
        --  M is the new multiplicity.
     raises ConstructionError,
        ---Purpose :
        --  M should be greater than the previous multiplicity and lower 
        --  than the degree of the surface in the V parametric direction.
            OutOfRange;
        ---Purpose :
        --  Raised if VIndex is not in the range [FirstVKnotIndex, 
        --  LastVKnotIndex] given by the methods with the same name.


  IncreaseVMultiplicity (me : mutable; FromI1, ToI2 : Integer; M : Integer)
        ---Purpose :
        --  Increases until order M the multiplicity of the set of knots
        --  FromI1,...., ToI2 in the V direction. This method can be used to
        --  make a BSplineSurface into a PiecewiseBezier B_spline
        --  surface. If <me> was uniform, it can become non-uniform.
     raises OutOfRange,
        ---Purpose :
        --  Raised if FromI1 or ToI2 is out of the range [FirstVKnotIndex,
        --  LastVKnotIndex] given by the methods with the same name.
            ConstructionError;
        ---Purpose : 
        --  M should be greater than the previous multiplicity of the
        --  all the knots FromI1,..., ToI2 and lower or equal to the
        --  Degree of the surface in the V parametric direction.


  IncrementVMultiplicity (me : mutable; FromI1, ToI2 : Integer; Step : Integer)
        ---Purpose :
        --  Increments the multiplicity of the consecutives vknots FromI1..ToI2
        --  by step.  The multiplicity of each knot FromI1,.....,ToI2 must be
        --  lower or equal to the VDegree of the B_spline.
     raises OutOfRange,
        ---Purpose :
        --  Raised if FromI1 or ToI2 is not in the range
        --  [FirstVKnotIndex, LastVKnotIndex] 
            ConstructionError;
        ---Purpose :
        --  Raised if one knot has a multiplicity greater than VDegree.


  InsertUKnot (me : mutable; U : Real; M : Integer; ParametricTolerance : Real;
     	    	    	     Add : Boolean = Standard_True)
        ---Purpose:
        --  Inserts a knot value in the sequence of UKnots. If U is a knot
        --  value this method increases the multiplicity of the knot if the
        --  previous multiplicity was lower than M else it does nothing. The
        --  tolerance criterion is ParametricTolerance. ParametricTolerance
        --  should be greater or equal than Resolution from package gp.
     raises ConstructionError;
        ---Purpose :
        --  Raised if U is out of the bounds [U1, U2] given by the methods 
        --  Bounds, the criterion ParametricTolerance is used.
        --  Raised if M is not in the range [1, UDegree].


  InsertVKnot (me : mutable; V : Real; M : Integer; ParametricTolerance : Real;
                             Add : Boolean = Standard_True)
        ---Purpose :
        --  Inserts a knot value in the sequence of VKnots. If V is a knot
        --  value this method increases the multiplicity of the knot if the
        --  previous multiplicity was lower than M otherwise it does nothing.
        --  The tolerance criterion is ParametricTolerance.
        --  ParametricTolerance should be greater or equal than Resolution
        --  from package gp.
     raises ConstructionError;
        ---Purpose :
        --  raises if V is out of the Bounds [V1, V2] given by the methods 
        --  Bounds, the criterion ParametricTolerance is used.
        --  raises if M is not in the range [1, VDegree].


  Segment (me : mutable; U1, U2, V1, V2 : Real)
        ---Purpose :
        --  Segments the surface between U1 and U2 in the U-Direction.
        --                       between V1 and V2 in the V-Direction.
        --  The control points are modified, the first and the last point
        --  are not the same.
        -- Warnings :
        --  Even if <me> is not closed it can become closed after the 
        --  segmentation for example if U1 or U2 are out of the bounds 
        --  of the surface <me> or if the surface makes loop.
    raises DomainError from Standard;
	---Purpose: raises if U2 < U1 or V2 < V1


  CheckAndSegment (me : mutable; U1, U2, V1, V2 : Real)
        ---Purpose :
        --  Segments the surface between U1 and U2 in the U-Direction.
        --                       between V1 and V2 in the V-Direction.
        --                       
        --  same as Segment but do nothing if U1 and U2 (resp. V1 and V2) are
        --  equal to the bounds in U (resp. in V) of <me>. 
        --  For example, if <me> is periodic in V, it will be always periodic
        --  in V after the segmentation if the bounds in V are unchanged
        --  
        -- Warnings : 
        --  Even if <me> is not closed it can become closed after the 
        --  segmentation for example if U1 or U2 are out of the bounds 
        --  of the surface <me> or if the surface makes loop.
    raises DomainError from Standard;
	---Purpose: raises if U2 < U1 or V2 < V1


  SetUKnot (me : mutable; UIndex : Integer; K : Real)
        ---Purpose :  Substitutes the UKnots of range UIndex with K.
     raises OutOfRange,
        ---Purpose :
        --  Raised if UIndex < 1 or UIndex > NbUKnots
            ConstructionError;
	---Purpose :
	--  Raised if K >= UKnots(UIndex+1) or K <= UKnots(UIndex-1)


  SetUKnots (me : mutable; UK : Array1OfReal from TColStd)
	---Purpose :  Changes all the U-knots of the surface.
        --  The multiplicity of the knots are not modified.
     raises ConstructionError,
	---Purpose : 
	--  Raised if there is an index such that UK (Index+1) <= UK (Index).
            OutOfRange;
        ---Purpose : 
        --  Raised if  UK.Lower() < 1 or UK.Upper() > NbUKnots


  SetUKnot (me : mutable; UIndex : Integer; K : Real; M : Integer)
        ---Purpose :  
        --  Changes the value of the UKnots of range UIndex and 
        --  increases its multiplicity.
     raises OutOfRange,
        ---Purpose :
        --  Raised if UIndex is not in the range [FirstUKnotIndex,
        --  LastUKnotIndex] given by the methods with the same name.
            ConstructionError;
	---Purpose :
	--  Raised if K >= UKnots(UIndex+1) or K <= UKnots(UIndex-1)
        --  M must be lower than UDegree and greater than the previous 
        --  multiplicity of the knot of range UIndex.


  SetVKnot (me : mutable; VIndex : Integer; K : Real)
        ---Purpose :  Substitutes the VKnots of range VIndex with K.
     raises OutOfRange,
        ---Purpose :
        --  Raised if VIndex < 1 or VIndex > NbVKnots
            ConstructionError;
	---Purpose :
	--  Raised if K >= VKnots(VIndex+1) or K <= VKnots(VIndex-1)


  SetVKnots (me : mutable; VK : Array1OfReal from TColStd)
	---Purpose :  Changes all the V-knots of the surface.
        --  The multiplicity of the knots are not modified.
     raises ConstructionError,
	---Purpose : 
	--  Raised if there is an index such that VK (Index+1) <= VK (Index).
            OutOfRange;
        ---Purpose : 
        --  Raised if  VK.Lower() < 1 or VK.Upper() > NbVKnots



  SetVKnot (me : mutable; VIndex : Integer; K : Real; M : Integer)
        ---Purpose :  
        --  Changes the value of the VKnots of range VIndex and increases 
        --  its multiplicity.
     raises OutOfRange,
        ---Purpose :
        --  Raised if VIndex is not in the range [FirstVKnotIndex,
        --  LastVKnotIndex] given by the methods with the same name.
            ConstructionError;
	---Purpose :
	--  Raised if K >= VKnots(VIndex+1) or K <= VKnots(VIndex-1)
        --  M must be lower than VDegree and greater than the previous 
        --  multiplicity of the knot of range VIndex.


  LocateU (me;
           U                   : Real; 
           ParametricTolerance : Real;
           I1, I2              : in out Integer;
           WithKnotRepetition  : Boolean = Standard_False);
        ---Purpose :
        --  Locates the parametric value U in the sequence of UKnots.
        --  If "WithKnotRepetition" is True we consider the knot's
        --  representation with repetition of multiple knot value,
        --  otherwise  we consider the knot's representation with
        --  no repetition of multiple knot values.
        --  UKnots (I1) <= U <= UKnots (I2)
        --  . if I1 = I2  U is a knot value (the tolerance criterion 
        --    ParametricTolerance is used).
        --  . if I1 < 1  => U < UKnots(1) - Abs(ParametricTolerance)
        --  . if I2 > NbUKnots => U > UKnots(NbUKnots)+Abs(ParametricTolerance)


  LocateV (me; 
           V                   : Real; 
           ParametricTolerance : Real;
           I1, I2              : in out Integer;
           WithKnotRepetition  : Boolean = Standard_False);
        ---Purpose :
        --  Locates the parametric value U in the sequence of knots.
        --  If "WithKnotRepetition" is True we consider the knot's
        --  representation with repetition of multiple knot value,
        --  otherwise  we consider the knot's representation with
        --  no repetition of multiple knot values.
        --  VKnots (I1) <= V <= VKnots (I2)
        --  . if I1 = I2  V is a knot value (the tolerance criterion 
        --    ParametricTolerance is used).
        --  . if I1 < 1  => V < VKnots(1) - Abs(ParametricTolerance)
        --  . if I2 > NbVKnots => V > VKnots(NbVKnots)+Abs(ParametricTolerance)







        ---Purpose :  poles insertion and removing
        --  The following methods are available only if the surface
        --  is Uniform or QuasiUniform in the considered direction
        --  The knot repartition is modified.




        ----Purpose : poles and weights modifications

  SetPole (me : mutable; UIndex, VIndex : Integer; P : Pnt)
        ---Purpose :
        --  Substitutes the pole of range (UIndex, VIndex) with P.
        --  If the surface is rational the weight of range (UIndex, VIndex)
        --  is not modified.
     raises OutOfRange;
        ---Purpose :
        --  Raised if UIndex < 1 or UIndex > NbUPoles or VIndex < 1 or
        --  VIndex > NbVPoles.


  SetPole (me : mutable; UIndex, VIndex : Integer; P : Pnt; Weight : Real)
        ---Purpose :
        --  Substitutes the pole and the weight of range (UIndex, VIndex)
        --  with P and W.
     raises OutOfRange,
        ---Purpose :
        --  Raised if UIndex < 1 or UIndex > NbUPoles or VIndex < 1 or
        --  VIndex > NbVPoles.
            ConstructionError;
	---Purpose : Raised if Weight <= Resolution from package gp.


  SetPoleCol (me : mutable; VIndex : Integer; CPoles : Array1OfPnt from TColgp)
         ---Purpose :
         --  Changes a column of poles or a part of this column.
     raises OutOfRange,
        ---Purpose : Raised if Vindex < 1 or VIndex > NbVPoles.
            ConstructionError;
	---Purpose :
	--  Raised if CPoles.Lower() < 1 or CPoles.Upper() > NbUPoles.


  SetPoleCol (me : mutable; VIndex : Integer; CPoles : Array1OfPnt from TColgp;
              CPoleWeights : Array1OfReal from TColStd)
         ---Purpose :
         --  Changes a column of poles or a part of this column with the
         --  corresponding weights. If the surface was rational it can
         --  become non rational. If the surface was non rational it can
         --  become rational.
     raises OutOfRange,
        ---Purpose : Raised if Vindex < 1 or VIndex > NbVPoles.
            ConstructionError;
	---Purpose :
	--  Raised if CPoles.Lower() < 1 or CPoles.Upper() > NbUPoles
	--  Raised if the bounds of CPoleWeights are not the same as the
	--  bounds of CPoles.
	--  Raised if one of the weight value of CPoleWeights is lower or
	--  equal to Resolution from package gp.


  SetPoleRow (me : mutable; UIndex : Integer; CPoles : Array1OfPnt from TColgp;
              CPoleWeights : Array1OfReal from TColStd)
         ---Purpose :
         --  Changes a row of poles or a part of this row with the
         --  corresponding weights. If the surface was rational it can
         --  become non rational. If the surface was non rational it can
         --  become rational.
     raises OutOfRange,
        ---Purpose : Raised if Uindex < 1 or UIndex > NbUPoles.
            ConstructionError;
	---Purpose :
	--  Raised if CPoles.Lower() < 1 or CPoles.Upper() > NbVPoles
	--  raises if the bounds of CPoleWeights are not the same as the
	--  bounds of CPoles.
	--  Raised if one of the weight value of CPoleWeights is lower or
	--  equal to Resolution from package gp.


  SetPoleRow (me : mutable; UIndex : Integer; CPoles : Array1OfPnt from TColgp)
         ---Purpose :
         --  Changes a row of poles or a part of this row.
     raises OutOfRange,
        ---Purpose : Raised if Uindex < 1 or UIndex > NbUPoles.
            ConstructionError;
	---Purpose :
	--  Raised if CPoles.Lower() < 1 or CPoles.Upper() > NbVPoles.


  SetWeight (me : mutable; UIndex, VIndex : Integer; Weight : Real)
        ---Purpose :
        --  Changes the weight of the pole of range UIndex, VIndex.
        --  If the surface was non rational it can become rational.
        --  If the surface was rational it can become non rational.
     raises OutOfRange,
        ---Purpose : 
        --  Raised if UIndex < 1 or UIndex > NbUPoles or VIndex < 1 or
        --  VIndex > NbVPoles
            ConstructionError;
        ---Purpose : 
        --  Raised if weight is lower or equal to Resolution from 
        --  package gp


  SetWeightCol (me : mutable; VIndex : Integer;
    	        CPoleWeights : Array1OfReal from TColStd)
        ---Purpose :
        --  Changes a column of weights of a part of this column.
     raises OutOfRange,
        ---Purpose : 
        --  Raised if VIndex < 1 or VIndex > NbVPoles
            ConstructionError;
	---Purpose :
	--  Raised if CPoleWeights.Lower() < 1 or 
	--            CPoleWeights.Upper() > NbUPoles.
        --  Raised if a weight value is lower or equal to Resolution
        --  from package gp.


  SetWeightRow (me : mutable; UIndex : Integer;
    	        CPoleWeights : Array1OfReal from TColStd)
        ---Purpose :  
        --  Changes a row of weights or a part of this row.
     raises OutOfRange,
        ---Purpose : 
        --  Raised if UIndex < 1 or UIndex > NbUPoles
            ConstructionError;
	---Purpose :
	--  Raised if CPoleWeights.Lower() < 1 or 
	--            CPoleWeights.Upper() > NbVPoles.
        --  Raised  if a weight value is lower or equal to Resolution
        --  from package gp.

  MovePoint(me: mutable; U, V : Real; P: Pnt;
    	    UIndex1, UIndex2, VIndex1, VIndex2: Integer;
            UFirstIndex, ULastIndex, VFirstIndex, VLastIndex: out Integer)
      ---Purpose: Move a point with parameter U and V to P.
      --          given u,v  as parameters)  to  reach a  new position
      --          UIndex1, UIndex2, VIndex1, VIndex2:
      --                  indicates the poles which can be moved      
      --          if Problem in BSplineBasis calculation, no change
      --          for the curve and
      --              UFirstIndex, VLastIndex = 0
      --              VFirstIndex, VLastIndex = 0
     raises OutOfRange;
        ---Purpose:
        --  Raised if UIndex1 < UIndex2 or VIndex1 < VIndex2 or
        --            UIndex1 < 1 || UIndex1 > NbUPoles or
        --            UIndex2 < 1 || UIndex2 > NbUPoles
        --            VIndex1 < 1 || VIndex1 > NbVPoles or
        --            VIndex2 < 1 || VIndex2 > NbVPoles



        ---Purpose : characteristics of the surface

  IsUClosed (me)  returns Boolean;
        ---Purpose :
        --  Returns true if the first control points row and the last
        --  control points row are identical. The tolerance criterion
        --  is Resolution from package gp.

  IsVClosed (me)   returns Boolean;
        ---Purpose :
        --  Returns true if the first control points column and the
        --  last last control points column are identical. 
        --  The tolerance criterion is Resolution from package gp.


  IsCNu (me; N : Integer)  returns Boolean
        ---Purpose :
        --  Returns True if the order of continuity of the surface in the 
        --  U direction  is N.
     raises RangeError;
        ---Purpose : Raised if N < 0.


  IsCNv (me; N : Integer)   returns Boolean
        ---Purpose :
        --  Returns True if the order of continuity of the surface 
        --  in the V direction  is N.
     raises RangeError;
        ---Purpose : Raised if N < 0.


  IsUPeriodic (me)  returns Boolean;
        ---Purpose :
        --  Returns True if the surface is closed in the U direction
        --  and if the B-spline has been turned into a periodic surface
        --  using the function SetUPeriodic.


  IsURational (me)   returns Boolean;
        ---Purpose :
        --  Returns False if for each row of weights all the weights
        --  are identical.
        --  The tolerance criterion is resolution from package gp.
        --  Example :
        --                 |1.0, 1.0, 1.0|
        --   if Weights =  |0.5, 0.5, 0.5|   returns False
        --                 |2.0, 2.0, 2.0|


  IsVPeriodic (me)  returns Boolean;
        ---Purpose :
        --  Returns True if the surface is closed in the V direction
        --  and if the B-spline has been turned into a periodic 
        --  surface using the function SetVPeriodic.


  IsVRational (me)  returns Boolean;
        ---Purpose :
        --  Returns False if for each column of weights all the weights 
        --  are identical.
        --  The tolerance criterion is resolution from package gp.
        --- Examples :
        --                 |1.0, 2.0, 0.5|
        --   if Weights =  |1.0, 2.0, 0.5|   returns False
        --                 |1.0, 2.0, 0.5|

  IsCacheValid(me;  UParameter, VParameter : Real) returns Boolean ;
  
        ---Purpose :
        --           Tells whether the Cache is valid for the
        --           given parameter 
        -- Warnings : the parameter must be normalized within
        -- the period if the curve is periodic. Otherwise
        -- the answer will be false
        -- 
        
  Bounds (me; U1, U2, V1, V2 : out Real);
        ---Purpose :
        --  Returns the parametric bounds of the surface.
        --- Warnings :
        --  These parametric values are the bounds of the array of
        --  knots UKnots and VKnots only if the first knots and the
        --  last knots have a multiplicity equal to UDegree + 1 or
        --  VDegree + 1


  Continuity (me)   returns Shape from GeomAbs;
        ---Purpose :
        --  Returns the continuity of the surface : 
        --  C0 : only geometric continuity,
        --  C1 : continuity of the first derivative all along the Surface,
        --  C2 : continuity of the second derivative all along the Surface,
        --  C3 : continuity of the third derivative all along the Surface,
        --  CN : the order of continuity is infinite.
        --  A B-spline surface is infinitely continuously differentiable 
        --  for the couple of parameters U, V such thats U != UKnots(i) 
        --  and V != VKnots(i). The continuity of the surface at a knot 
        --  value depends on the multiplicity of this knot.
        --- Example :
        --  If the surface is C1 in the V direction and C2 in the U 
        --  direction this function returns Shape = C1.


  FirstUKnotIndex (me)   returns Integer;
        ---Purpose :
        --  Computes the Index of the UKnots which gives the first 
        --  parametric value of the surface in the U direction.
        --  The UIso curve corresponding to this value is a 
        --  boundary curve of the surface.


  FirstVKnotIndex (me)   returns Integer;
        ---Purpose :
        --  Computes the Index of the VKnots which gives the
        --  first parametric value of the surface in the V direction.
        --  The VIso curve corresponding to this knot is a boundary
        --  curve of the surface.
     
     
  LastUKnotIndex (me)   returns Integer;
        ---Purpose :
        --  Computes the Index of the UKnots which gives the 
        --  last parametric value of the surface in the U direction.
        --  The UIso curve corresponding to this knot is a boundary 
        --  curve of the surface.
     
     
  LastVKnotIndex (me)   returns Integer;
        ---Purpose :
        --  Computes the Index of the VKnots which gives the 
        --  last parametric value of the surface in the V direction.
        --  The VIso curve corresponding to this knot is a
        --  boundary curve of the surface.


  NbUKnots (me)   returns Integer;
        ---Purpose :  Returns the number of knots in the U direction. 

  NbUPoles (me)  returns Integer;
        ---Purpose : Returns number of poles in the U direction.

  NbVKnots (me)  returns Integer;
        ---Purpose : Returns the number of knots in the V direction.

  NbVPoles (me)  returns Integer;
        ---Purpose : Returns the number of poles in the V direction.


  Pole (me; UIndex, VIndex : Integer)   returns Pnt
        ---Purpose: 
        --  Returns the pole of range (UIndex, VIndex).
     raises OutOfRange;
        ---Purpose :
        --  Raised if UIndex < 1 or UIndex > NbUPoles or VIndex < 1 or
        --  VIndex > NbVPoles.


  Poles (me; P : out Array2OfPnt from TColgp)
       ---Purpose : Returns the poles of the B-spline surface.
     raises DimensionError;
       ---Purpose :
       --  Raised if the length of P in the U and V direction
       --  is not equal to NbUpoles and NbVPoles.
  Poles (me)
  returns Array2OfPnt from TColgp
       ---Purpose : Returns the poles of the B-spline surface.
       ---C++ : return const &
  is static;


  UDegree (me)  returns Integer;
        ---Purpose :
        --  Returns the degree of the normalized B-splines Ni,n in the U
        --  direction.


  UKnot (me; UIndex : Integer)  returns Real
        ---Purpose :
        --  Returns the Knot value of range UIndex.
     raises OutOfRange;
        ---Purpose : Raised if UIndex < 1 or UIndex > NbUKnots


  UKnotDistribution (me)   returns BSplKnotDistribution from GeomAbs;
        ---Purpose :
        --  Returns NonUniform or Uniform or QuasiUniform or 
        --  PiecewiseBezier.  If all the knots differ by a
        --  positive constant from the preceding knot in the U 
        --  direction the B-spline surface can be :
        --  - Uniform if all the knots are of multiplicity 1,
        --  - QuasiUniform if all the knots are of multiplicity 1
        --    except for the first and last knot which are of 
        --    multiplicity Degree + 1,
        --  - PiecewiseBezier if the first and last knots have 
        --    multiplicity Degree + 1 and if interior knots have
        --    multiplicity Degree
        --  otherwise the surface is non uniform in the U direction 
        --  The tolerance criterion is Resolution from package gp.


  UKnots (me; Ku : out Array1OfReal from TColStd)
       	---Purpose : Returns the knots in the U direction.
     raises DimensionError;
       	---Purpose :
       	--  Raised if the length of Ku is not equal to the number of knots
       	--  in the U direction.
  UKnots (me)
  returns Array1OfReal from TColStd
       ---Purpose : Returns the knots in the U direction.
       ---C++ : return const &
  is static;


  UKnotSequence (me; Ku : out Array1OfReal from TColStd)
        ---Purpose : Returns the uknots sequence.
        --  In this sequence the knots with a multiplicity greater than 1
        --  are repeated.
        --- Example :
        --  Ku = {k1, k1, k1, k2, k3, k3, k4, k4, k4}
     raises DimensionError;
        ---Purpose :
        --  Raised if the length of Ku is not equal to NbUPoles + UDegree + 1
  UKnotSequence (me)
  returns Array1OfReal from TColStd
        ---Purpose : Returns the uknots sequence.
        --  In this sequence the knots with a multiplicity greater than 1
        --  are repeated.
        --- Example :
        --  Ku = {k1, k1, k1, k2, k3, k3, k4, k4, k4}
        ---C++ : return const &
  is static;


  UMultiplicity (me; UIndex : Integer)   returns Integer
        ---Purpose :
        --  Returns the multiplicity value of knot of range UIndex in 
        --  the u direction.
     raises OutOfRange;
        ---Purpose : Raised if UIndex < 1 or UIndex > NbUKnots.


  UMultiplicities (me; Mu : out Array1OfInteger from TColStd)
       	---Purpose : 
       	--  Returns the multiplicities of the knots in the U direction.
     raises DimensionError;
       	---Purpose :
       	--  Raised if the length of Mu is not equal to the number of
       	--  knots in the U direction.
  UMultiplicities (me)
  returns Array1OfInteger from TColStd
       ---Purpose : Returns the multiplicities of the knots in the U direction.
       ---C++ : return const &
  is static;


  VDegree (me)  returns Integer;
        ---Purpose : 
        --  Returns the degree of the normalized B-splines Ni,d in the 
        --  V direction.


  VKnot (me; VIndex : Integer)   returns Real
        ---Purpose : Returns the Knot value of range VIndex.
     raises OutOfRange;
        --- Purpse : Raised if VIndex < 1 or VIndex > NbVKnots


  VKnotDistribution (me)  returns BSplKnotDistribution from GeomAbs;
        ---Purpose :
        --  Returns NonUniform or Uniform or QuasiUniform or
        --  PiecewiseBezier. If all the knots differ by a positive
        --  constant from the preceding knot in the V direction the
        --  B-spline surface can be :
        --  - Uniform if all the knots are of multiplicity 1,
        --  - QuasiUniform if all the knots are of multiplicity 1 
        --    except for the first and last knot which are of 
        --    multiplicity Degree + 1,
        --  - PiecewiseBezier if the first and last knots have
        --    multiplicity  Degree + 1 and if interior knots have
        --     multiplicity Degree
        --  otherwise the surface is non uniform in the V direction.
        --  The tolerance criterion is Resolution from package gp.


  VKnots (me; Kv : out Array1OfReal from TColStd)
       ---Purpose : Returns the knots in the V direction.
     raises DimensionError;
       ---Purpose :
       --  Raised if the length of Kv is not equal to the number of 
       --  knots in the V direction.
  VKnots (me)
  returns Array1OfReal from TColStd
       ---Purpose : Returns the knots in the V direction.
       ---C++ : return const &
  is static;


  VKnotSequence (me; Kv : out Array1OfReal from TColStd)
        ---Purpose : Returns the vknots sequence.
        --  In this sequence the knots with a multiplicity greater than 1
        --  are repeated. 
        --- Example :
        --  Kv = {k1, k1, k1, k2, k3, k3, k4, k4, k4}
     raises DimensionError;
        ---Purpose :
        --  Raised if the length of Kv is not equal to NbVPoles + VDegree + 1
  VKnotSequence (me)
  returns Array1OfReal from TColStd
        ---Purpose : Returns the vknots sequence.
        --  In this sequence the knots with a multiplicity greater than 1
        --  are repeated.
        --- Example :
        --  Ku = {k1, k1, k1, k2, k3, k3, k4, k4, k4}
        ---C++ : return const &
  is static;


  VMultiplicity (me; VIndex : Integer)   returns Integer
        ---Purpose :
        --  Returns the multiplicity value of knot of range VIndex in 
        --  the v direction.
     raises OutOfRange;
        ---Purpose : Raised if VIndex < 1 or VIndex > NbVKnots

  
  VMultiplicities (me; Mv : out Array1OfInteger from TColStd)
       ---Purpose :
       --  Returns the multiplicities of the knots in the V direction.
     raises DimensionError;
       ---Purpose :
       --  Raised if the length of Mv is not equal to the number of 
       --  knots in the V direction.
  VMultiplicities (me)
  returns Array1OfInteger from TColStd
       ---Purpose : Returns the multiplicities of the knots in the V direction.
       ---C++ : return const &
  is static;


  Weight (me; UIndex, VIndex : Integer)   returns Real
        ---Purpose : Returns the weight value of range UIndex, VIndex.
     raises OutOfRange;
        ---Purpose : 
        --  Raised if UIndex < 1 or UIndex > NbUPoles or VIndex < 1
        --  or VIndex > NbVPoles.

  
  Weights (me; W : out Array2OfReal from TColStd)
        ---Purpose : Returns the weights of the B-spline surface.
     raises DimensionError;
        ---Purpose :
        --  Raised if the length of W in the U and V direction is 
        --  not equal to NbUPoles and NbVPoles.
  Weights (me)
  returns Array2OfReal from TColStd
        ---Purpose : Returns the weights of the B-spline surface.
        ---C++ : return const &
  is static;






        ---Purpose : value and derivatives computation

  D0 (me; U, V : Real; P : out Pnt);


  D1 (me; U, V : Real; P : out Pnt; D1U, D1V : out Vec)
     raises UndefinedDerivative;
        ---Purpose : Raised if the continuity of the surface is not C1.


  D2 (me; U, V : Real; P : out Pnt; D1U, D1V, D2U, D2V, D2UV : out Vec)
     raises UndefinedDerivative;
        ---Purpose : Raised if the continuity of the surface is not C2.


  D3 (me; U, V : Real; P : out Pnt; D1U, D1V, D2U, D2V, D2UV, D3U, D3V, D3UUV,
      D3UVV : out Vec)
     raises UndefinedDerivative;
        ---Purpose : Raised if the continuity of the surface is not C3.


  DN (me; U, V : Real; Nu, Nv : Integer)   returns Vec
        ---Purpose :
        --  Nu is the order of derivation in the U parametric direction and
        --  Nv is the order of derivation in the V parametric direction.
     raises UndefinedDerivative,
        ---Purpose :
        --  Raised if the continuity of the surface is not CNu in the U
        --  direction and CNv in the V direction.
            RangeError;
        ---Purpose :
        --  Raised if Nu + Nv < 1 or Nu < 0 or Nv < 0.






        ---Purpose  :
        --  The following functions computes the point for the
        --  parametric values (U, V) and the derivatives at 
        --  this point on the B-spline surface patch delimited
        --  with the knots FromUK1, FromVK1 and the knots ToUK2,
        --  ToVK2.  (U, V) can be out of these parametric bounds
        --  but for the computation we only use the definition
        --  of the surface between these knots. This method is 
        --  useful to compute local derivative, if the order of
        --  continuity of the whole surface is not greater enough.
        --  Inside the parametric knot's domain previously defined
        --  the evaluations are the same as if we consider the whole
        --  definition of the surface. Of course the evaluations are
        --  different outside this parametric domain.


  LocalD0 (me; U, V : Real; FromUK1, ToUK2, FromVK1, ToVK2 : Integer;
    	       P : out Pnt)
     raises DomainError,
	---Purpose : Raised if FromUK1 = ToUK2 or FromVK1 = ToVK2.
            OutOfRange;
	---Purpose :
	--  Raised if FromUK1, ToUK2 are not in the range [FirstUKnotIndex,
	--  LastUKnotIndex] or if FromVK1, ToVK2 are not in the range
	--  [FirstVKnotIndex, LastVKnotIndex]


  LocalD1 (me; U, V : Real;  FromUK1, ToUK2, FromVK1, ToVK2 : Integer;
          P : out Pnt; D1U, D1V : out Vec)
     raises UndefinedDerivative,
        ---Purpose :
        --  Raised if the local continuity of the surface is not C1 
        --  between the knots FromUK1, ToUK2 and FromVK1, ToVK2. 
            DomainError,
	---Purpose : Raised if FromUK1 = ToUK2 or FromVK1 = ToVK2.
            OutOfRange;
	---Purpose :
	--  Raised if FromUK1, ToUK2 are not in the range [FirstUKnotIndex,
	--  LastUKnotIndex] or if FromVK1, ToVK2 are not in the range
	--  [FirstVKnotIndex, LastVKnotIndex]


  LocalD2 (me; U, V : Real; FromUK1, ToUK2, FromVK1, ToVK2 : Integer;
           P : out Pnt; D1U, D1V, D2U, D2V, D2UV : out Vec)
     raises UndefinedDerivative,
        ---Purpose :
        --  Raised if the local continuity of the surface is not C2 
        --  between the knots FromUK1, ToUK2 and FromVK1, ToVK2. 
            DomainError,
	---Purpose : Raised if FromUK1 = ToUK2 or FromVK1 = ToVK2.
            OutOfRange;
	---Purpose :
	--  Raised if FromUK1, ToUK2 are not in the range [FirstUKnotIndex,
	--  LastUKnotIndex] or if FromVK1, ToVK2 are not in the range
	--  [FirstVKnotIndex, LastVKnotIndex]


  LocalD3 (me; U, V : Real; FromUK1, ToUK2, FromVK1, ToVK2 : Integer;
           P : out Pnt; D1U, D1V, D2U, D2V, D2UV, D3U, D3V, D3UUV, D3UVV :
           out Vec)
     raises UndefinedDerivative,
        ---Purpose :
        --  Raised if the local continuity of the surface is not C3
        --  between the knots FromUK1, ToUK2 and FromVK1, ToVK2. 
            DomainError,
	---Purpose : Raised if FromUK1 = ToUK2 or FromVK1 = ToVK2.
            OutOfRange;
	---Purpose :
	--  Raised if FromUK1, ToUK2 are not in the range [FirstUKnotIndex,
	--  LastUKnotIndex] or if FromVK1, ToVK2 are not in the range
	--  [FirstVKnotIndex, LastVKnotIndex]


  LocalDN (me; U, V : Real; FromUK1, ToUK2, FromVK1, ToVK2 : Integer; 
           Nu, Nv : Integer)
     returns Vec
     raises UndefinedDerivative,
        ---Purpose :
        --  Raised if the local continuity of the surface is not CNu 
        --  between the knots FromUK1, ToUK2 and CNv between the knots
        --  FromVK1, ToVK2. 
            DomainError,
	---Purpose : Raised if FromUK1 = ToUK2 or FromVK1 = ToVK2.
             RangeError,
        --  Raised if Nu + Nv < 1 or Nu < 0 or Nv < 0.
             OutOfRange;
	---Purpose :
	--  Raised if FromUK1, ToUK2 are not in the range [FirstUKnotIndex,
	--  LastUKnotIndex] or if FromVK1, ToVK2 are not in the range
	--  [FirstVKnotIndex, LastVKnotIndex]

  LocalValue(me; U, V : Real;  FromUK1, ToUK2, FromVK1, ToVK2 : Integer)
        ---Purpose  :
        --  Computes the point of parameter U, V on the BSpline surface patch 
        --  defines between the knots UK1 UK2, VK1, VK2. U can be out of the
        --  bounds [Knot UK1, Knot UK2] and V can be outof the bounds 
        --  [Knot VK1, Knot VK2]  but for the computation we only use the 
        --  definition of the surface between these knot values.
     returns Pnt
     raises DomainError,
	---Purpose : Raises if FromUK1 = ToUK2 or FromVK1 = ToVK2.
            OutOfRange;
	---Purpose :
	--  Raises if FromUK1, ToUK2 are not in the range [FirstUKnotIndex,
	--  LastUKnotIndex] or if FromVK1, ToVK2 are not in the range
	--  [FirstVKnotIndex, LastVKnotIndex]



  UIso (me; U : Real) returns Curve;
        ---Purpose :
        --  Computes the U isoparametric curve. 
        --  A B-spline curve is returned.


  VIso (me; V : Real)  returns Curve;
        ---Purpose :
        --  Computes the V isoparametric curve. 
        --  A B-spline curve is returned.


  UIso (me; U : Real; CheckRational : Boolean) returns Curve;
        ---Purpose :
        --  Computes the U isoparametric curve.  
	--  If CheckRational=False, no try to make it non-rational.
        --  A B-spline curve is returned.


  VIso (me; V : Real; CheckRational : Boolean) returns Curve;
        ---Purpose :
        --  Computes the V isoparametric curve. 
	--  If CheckRational=False, no try to make it non-rational.
        --  A B-spline curve is returned.




 
        ---Purpose : transformations

  Transform (me : mutable; T : Trsf) ;

    	--- Purpose: Applies the transformation T to this BSpline surface.

  MaxDegree (myclass)   returns Integer;
        ---Purpose :
        --  Returns the value of the maximum degree of the normalized 
        --  B-spline basis functions in the u and v directions.


  Resolution(me          : mutable; 
    	     Tolerance3D :     Real ;
    	     UTolerance  : out Real ;
	     VTolerance  : out Real) 
    	---Purpose: Computes two tolerance values for this BSpline
    	-- surface, based on the given tolerance in 3D space
    	-- Tolerance3D. The tolerances computed are:
    	-- - UTolerance in the u parametric direction, and
    	-- - VTolerance in the v parametric direction.
    	-- If f(u,v) is the equation of this BSpline surface,
    	-- UTolerance and VTolerance guarantee that :
      	--          | u1 - u0 | < UTolerance and 
      	--          | v1 - v0 | < VTolerance 
      	--          ====> |f (u1,v1) - f (u0,v0)| < Tolerance3D
  ;
  
  Copy (me)  returns like me;

    	---Purpose: Creates a new object which is a copy of this BSpline surface.

  UpdateUKnots(me : mutable)
        ---Purpose: Recompute  the  flatknots,  the knotsdistribution, the
    	--          continuity for U.
  is static private;

  UpdateVKnots(me : mutable)
    	---Purpose: Recompute  the  flatknots,  the knotsdistribution, the
	--          continuity for V.
  is static private;

  
  InvalidateCache(me : mutable)
    	---Purpose : Invalidates the cache. This has to be private this has to be private
      is static private;
      
  ValidateCache(me : mutable ; UParameter : Real; 
    	    	    	       VParameter : Real) 
  
    is static private;
    	---Purpose : updates the cache and validates it

  
fields
	     
   urational : Boolean;
   vrational : Boolean;
   uperiodic : Boolean;
   vperiodic : Boolean;
   uknotSet  : BSplKnotDistribution from GeomAbs; 
   vknotSet  : BSplKnotDistribution from GeomAbs; 
   Usmooth   : Shape from GeomAbs;
   Vsmooth   : Shape from GeomAbs;
   udeg      : Integer;
   vdeg      : Integer;
   poles     : HArray2OfPnt     from TColgp;
   weights   : HArray2OfReal    from TColStd;
   ufknots   : HArray1OfReal    from TColStd;
   vfknots   : HArray1OfReal    from TColStd;
   uknots    : HArray1OfReal    from TColStd;
   vknots    : HArray1OfReal    from TColStd;
   umults    : HArray1OfInteger from TColStd;
   vmults    : HArray1OfInteger from TColStd;
  -- Inplementation of the cache on surfaces
   cachepoles : HArray2OfPnt     from TColgp;
  -- Taylor expansion of the poles function, in homogeneous
  -- form if the curve is rational. The taylor expansion
  -- is normalized so that the span corresponds to
  -- [0 1]x[0 1]. The Taylor expension of lower degree
  -- is stored as consecutive Pnt in the array that is
  -- if udeg <= vdeg than the array stores the following
  -- 
  --                                  (2,0)           (3,0) 
  --               (1,0)             f     (u0,v0)   f     (u0,v0)
  --  f  (u0,v0)  f     (u0,v0)      -------------   -----------
  --                                      2             3!
  --                                
  --                                   (2,1)           (3,1) 
  --   (0,1)          (1,1)         f     (u0,v0)   f     (u0,v0)
  --  f     (u0,v0)  f     (u0,v0)  -------------   -----------
  --                                     2              3!
  --   
  -- Otherwise it is stored in the following fashion
  -- 
  --  
  --                                  (0,2)           (0,3) 
  --               (0,1)             f     (u0,v0)   f     (u0,v0)
  --  f  (u0,v0)  f     (u0,v0)      -------------   -----------
  --                                      2             3!
  --                                
  --                                 (1,2)           (1,3) 
  --   (1,0)          (1,1)         f     (u0,v0)   f     (u0,v0)
  --  f     (u0,v0)  f     (u0,v0)  -------------   -----------
  --                                     2              3!
  --   
  --   The size of the array is (1,Max degree) (1, Min degree) 
  -- 
    cacheweights   : HArray2OfReal    from TColStd;
  -- Taylor expansion of the poles function, in homogeneous
  -- form if the curve is rational. The taylor expansion
  -- is normalized so that the span corresponds to
  -- [0 1]x[0 1]. The Taylor expension of lower degree
  -- is stored as consecutive Real in the array as explained above
    ucacheparameter : Real ;
    vcacheparameter : Real ;
  -- Parameters at which the Taylor expension is stored in 
  -- the cache  
    ucachespanlenght : Real ;
    vcachespanlenght : Real ;
      -- Since the Taylor expansion is normalized in the 
  -- cache to evaluate the cache one has to use
  -- (UParameter - uparametercache) / ucachespanlenght
  -- (VParameter - vparametercache) / vcachespanlenght
    ucachespanindex : Integer ;
    vcachespanindex : Integer ;
  -- the span for which the cache is valid if 
  -- validcache is 1 
    validcache : Integer ;
    
  -- usefull to evaluate the parametric resolutions
    umaxderivinv  : Real from Standard;
    vmaxderivinv  : Real from Standard;
    maxderivinvok : Boolean from Standard;

    myMutex       : Mutex from Standard;
    -- protected bsplinesurface-cache

end;
