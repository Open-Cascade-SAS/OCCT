-- Created on: 1994-01-17
-- Created by: Modelistation
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PlaneAspect from Prs3d inherits BasicAspect from Prs3d
    	---Purpose: A framework to define the display of planes.
uses

    LineAspect from Prs3d,
    Length from Quantity,
    PlaneAngle from Quantity
    
is

    Create returns mutable PlaneAspect from Prs3d;
    	---Purpose: Constructs an empty framework for the display of planes.    
    EdgesAspect(me) returns mutable LineAspect from Prs3d;
    
    	---Purpose: Returns the attributes of displayed edges involved in the presentation of planes.    
    
    IsoAspect(me) returns mutable LineAspect from Prs3d;
    	---Purpose: Returns the attributes of displayed isoparameters involved in the presentation of planes.
        
    ArrowAspect(me) returns mutable LineAspect from Prs3d;
    	---Purpose: Returns the settings for displaying an arrow.    
    SetArrowsLength(me:mutable; L : Length from Quantity);
    
    
    ArrowsLength(me) returns Length from Quantity;
    	--- Purpose: Returns the length of the arrow shaft used in the display of arrows.   

    SetArrowsSize(me:mutable; L : Length from Quantity);
    	---Purpose: Sets the angle of the arrowhead used in the display of planes.    
    
    ArrowsSize(me) returns Length from Quantity;
    	---Purpose: Returns the size of arrows used in the display of planes.    
  
    SetArrowsAngle(me:mutable; ang : PlaneAngle from Quantity);
    	---Purpose: Sets the angle of the arrowhead used in the display
    	-- of arrows involved in the presentation of planes.    
    
    ArrowsAngle(me) returns PlaneAngle from Quantity;
    	---Purpose: Returns the angle of the arrowhead used in the
    	-- display of arrows involved in the presentation of planes.    
    
    SetDisplayCenterArrow(me:mutable ; draw: Boolean from Standard);
    	---Purpose: Sets the display attributes defined in DisplayCenterArrow to active.
    
    DisplayCenterArrow(me) returns Boolean from Standard;
    	---Purpose: Returns true if the display of center arrows is allowed.       
    SetDisplayEdgesArrows(me:mutable ; draw: Boolean from Standard);
    	---Purpose: Sets the display attributes defined in DisplayEdgesArrows to active. 
    
    DisplayEdgesArrows(me) returns Boolean from Standard;
 
    	--- Purpose: Returns true if the display of edge arrows is allowed.   
    SetDisplayEdges(me:mutable ; draw: Boolean from Standard);
    DisplayEdges(me) returns Boolean from Standard;
    
    SetDisplayIso(me:mutable ; draw: Boolean from Standard);
    	 ---Purpose: Sets the display attributes defined in DisplayIso to active.   
    
    DisplayIso(me) returns Boolean from Standard;
    	--- Purpose: Returns true if the display of isoparameters is allowed.   
    SetPlaneLength(me:mutable; LX,LY: Length from Quantity);
    PlaneXLength(me) returns Length from Quantity;
    	--- Purpose: Returns the length of the x axis used in the display of planes.   
    
    PlaneYLength(me) returns Length from Quantity;
    	---Purpose: Returns the length of the y axis used in the display of planes.    
    SetIsoDistance(me:mutable; L: Length from Quantity);
    	---Purpose: Sets the distance L between isoparameters used in the display of planes.  
    IsoDistance(me) returns Length from Quantity;
    	---Purpose: Returns the distance between isoparameters used in the display of planes.
        
fields

    myEdgesAspect: LineAspect from Prs3d;
    myIsoAspect: LineAspect from Prs3d;
    myArrowAspect: LineAspect from Prs3d;
    myArrowsLength: Length from Quantity;
    myArrowsSize: Length from Quantity;
    myArrowsAngle: PlaneAngle from Quantity;
    myDrawCenterArrow: Boolean from Standard;
    myDrawEdgesArrows: Boolean from Standard;
    myDrawEdges: Boolean from Standard;
    myDrawIso: Boolean from Standard;
    myPlaneXLength : Length from Quantity;    
    myPlaneYLength : Length from Quantity;    
    myIsoDistance: Length from Quantity;    

end PlaneAspect from Prs3d;

