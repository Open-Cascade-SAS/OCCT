-- Created on: 2000-05-10
-- Created by: Andrey BETENEV
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1

class AppliedExternalIdentificationAssignment from StepAP214
inherits ExternalIdentificationAssignment from StepBasic

    ---Purpose: Representation of STEP entity AppliedExternalIdentificationAssignment

uses
    HAsciiString from TCollection,
    IdentificationRole from StepBasic,
    ExternalSource from StepBasic,
    HArray1OfExternalIdentificationItem from StepAP214

is
    Create returns AppliedExternalIdentificationAssignment from StepAP214;
	---Purpose: Empty constructor

    Init (me: mutable; aIdentificationAssignment_AssignedId: HAsciiString from TCollection;
                       aIdentificationAssignment_Role: IdentificationRole from StepBasic;
                       aExternalIdentificationAssignment_Source: ExternalSource from StepBasic;
                       aItems: HArray1OfExternalIdentificationItem from StepAP214);
	---Purpose: Initialize all fields (own and inherited)

    Items (me) returns HArray1OfExternalIdentificationItem from StepAP214;
	---Purpose: Returns field Items
    SetItems (me: mutable; Items: HArray1OfExternalIdentificationItem from StepAP214);
	---Purpose: Set field Items

fields
    theItems: HArray1OfExternalIdentificationItem from StepAP214;

end AppliedExternalIdentificationAssignment;
