-- Created on: 1993-02-22
-- Created by: Modelistation
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class CurveOnSurface from Adaptor3d inherits Curve from Adaptor3d

	---Purpose: An interface between the services provided by a curve
    	-- lying on a surface from the package Geom and those
    	-- required of the curve by algorithms which use it. The
    	-- curve is defined as a 2D curve from the Geom2d
    	-- package, in the parametric space of the surface.


uses 
     Array1OfReal         from TColStd,
     Pnt                  from gp,
     Vec                  from gp,
     Circ                 from gp,
     Elips                from gp,
     Hypr                 from gp,
     Parab                from gp,
     Lin                  from gp,
     CurveType            from GeomAbs,
     Shape                from GeomAbs,
     BezierCurve          from Geom,
     BSplineCurve         from Geom,
     BSplineSurface       from Geom,   
     HCurve               from Adaptor3d,
     HCurve2d             from Adaptor2d,
     HSurface             from Adaptor3d,
     HSequenceOfReal      from TColStd,
     Pnt2d                from gp,
     Vec2d                from gp

raises NoSuchObject from Standard,
       DomainError  from Standard,
       OutOfRange   from Standard

is

    Create returns CurveOnSurface;
    
    Create(S : HSurface from Adaptor3d) returns CurveOnSurface;
    
    Create (C : HCurve2d from Adaptor2d; S : HSurface from Adaptor3d)
    returns CurveOnSurface;
	---Purpose: Creates a CurveOnSurface from the 2d curve <C> and
	--          the surface <S>.
   
    Load(me : in out;S : HSurface from Adaptor3d)
	---Purpose: Changes the surface.
    is static;
    
    Load(me : in out; C : HCurve2d from Adaptor2d)
	---Purpose: Changes the 2d curve.
    is static;

    GetCurve(me) returns HCurve2d from Adaptor2d
       ---C++: return const &
    is static;

    GetSurface(me) returns HSurface from Adaptor3d
       ---C++: return const &
    is static;

    ChangeCurve(me : in out) returns HCurve2d from Adaptor2d
       ---C++: return &
    is static;

    ChangeSurface(me : in out) returns HSurface from Adaptor3d
       ---C++: return &
    is static;

    --
    --      Implementation of Curve from Adaptor3d methods
    --      

    --
    --     Global methods - Apply to the whole curve.
    --     
    
    FirstParameter(me) returns Real
    is redefined static;

    LastParameter(me) returns Real
    is redefined static;
    
    Continuity(me) returns Shape from GeomAbs
    is redefined static;
    
    NbIntervals(me; S : Shape from GeomAbs) returns Integer
	---Purpose: Returns  the number  of  intervals for  continuity
	--          <S>. May be one if Continuity(me) >= <S>
    is redefined static;
    
    Intervals(me; T : in out Array1OfReal from TColStd; 
    	          S : Shape from GeomAbs)
	---Purpose: Stores in <T> the  parameters bounding the intervals
	--          of continuity <S>.
	--          
	--          The array must provide  enough room to  accomodate
	--          for the parameters. i.e. T.Length() > NbIntervals()
    raises
    	OutOfRange from Standard 
    is redefined static;
    
    Trim(me; First, Last, Tol : Real) returns HCurve from Adaptor3d
	---Purpose: Returns    a  curve equivalent   of  <me>  between
	--          parameters <First>  and <Last>. <Tol>  is used  to
	--          test for 3d points confusion.
    raises
    	OutOfRange from Standard
	---Purpose: If <First> >= <Last> 
    is redefined static;

    IsClosed(me) returns Boolean
    is redefined static;
     
    IsPeriodic(me) returns Boolean
    is redefined static;
    
    Period(me) returns Real
    raises
    	DomainError from Standard -- if the curve is not periodic
    is redefined static;
     
    Value(me; U : Real) returns Pnt from gp
         --- Purpose : Computes the point of parameter U on the curve.
    is redefined static;
    
    D0 (me; U : Real; P : out Pnt from gp)
         --- Purpose : Computes the point of parameter U on the curve.
    is redefined static;
    
    D1 (me; U : Real; P : out Pnt from gp ; V : out Vec from gp)
         --- Purpose : Computes the point of parameter U on the curve with its
         --  first derivative.
     raises 
    	DomainError from Standard
        --- Purpose : Raised if the continuity of the current interval
        --  is not C1.
    is redefined static;
    
    D2 (me; U : Real; P : out Pnt from gp; V1, V2 : out Vec from gp)
        --- Purpose :
        --  Returns the point P of parameter U, the first and second
        --  derivatives V1 and V2.
     raises 
    	DomainError from Standard
        --- Purpose : Raised if the continuity of the current interval
        --  is not C2.
     is redefined static;

    D3 (me; U : Real; P : out Pnt from gp; V1, V2, V3 : out Vec from gp)
        --- Purpose :
        --  Returns the point P of parameter U, the first, the second 
        --  and the third derivative.
     raises 
    	DomainError from Standard
        --- Purpose : Raised if the continuity of the current interval
        --  is not C3.
     is redefined static;
        
    DN (me; U : Real; N : Integer)   returns Vec from gp
        --- Purpose :
        --  The returned vector gives the value of the derivative for the 
        --  order of derivation N.
     raises  
    	DomainError from Standard,
        --- Purpose : Raised if the continuity of the current interval
        --  is not CN.
        OutOfRange from Standard
        --- Purpose : Raised if N < 1.            
     is redefined static;

    Resolution(me; R3d : Real) returns Real
         ---Purpose :  Returns the parametric  resolution corresponding
         --         to the real space resolution <R3d>.
    is redefined static;   
        
    GetType(me) returns CurveType from GeomAbs
	---Purpose: Returns  the  type of the   curve  in the  current
	--          interval :   Line,   Circle,   Ellipse, Hyperbola,
	--          Parabola, BezierCurve, BSplineCurve, OtherCurve.
    is redefined static;

    --
    --     The following methods must  be called when GetType returned
    --     the corresponding type.
    --     

     Line(me) returns Lin from gp
     raises 
    	NoSuchObject from Standard
     is redefined static;
     
     Circle(me) returns Circ from gp
     raises 
    	NoSuchObject from Standard
     is redefined static;
     
     Ellipse(me) returns Elips from gp
     raises 
    	NoSuchObject from Standard
     is redefined static;
     
     Hyperbola(me) returns  Hypr from gp
     raises 
    	NoSuchObject from Standard
     is redefined static;
     
     Parabola(me) returns Parab from gp
     raises 
    	NoSuchObject from Standard
     is redefined static;
     
     Degree(me) returns Integer
     raises 
    	NoSuchObject from Standard
     is redefined static;

     
     IsRational(me) returns Boolean
     raises 
    	NoSuchObject from Standard
     is redefined static;
     
     NbPoles(me) returns Integer
     raises 
    	NoSuchObject from Standard
     is redefined static;

  
     NbKnots(me) returns Integer
     raises 
    	NoSuchObject from Standard
     is redefined static;   
     ---Warning:  will raize if this asked on a curve
     --           that is not planar

     Bezier(me) returns BezierCurve from Geom
     raises 
    	NoSuchObject from Standard
     is redefined static;
    
     BSpline(me) returns BSplineCurve from Geom
     raises 
    	NoSuchObject from Standard
     is redefined static;
    
     EvalKPart(me : in out)
     is static private;
       
     EvalFirstLastSurf(me :  in  out) 
     	---Purpose:  Evaluates  myFirstSurf and myLastSurf 
        --	  for trimming the curve on surface.          
     is  static  private; 


        ---Purpose: Following  methods  output left-bottom and right-top points 
	--  of located part on surface  
	--  for trimming the curve on surface.      		
    
     LocatePart(me; UV : Pnt2d  from  gp; DUV : Vec2d from gp; 
    	S  :  HSurface  from  Adaptor3d; 
      LeftBot, RightTop : out Pnt2d from gp)  
     is  static  private;  

     LocatePart_RevExt(me; UV : Pnt2d  from  gp; DUV : Vec2d from gp; 
    	S  :  HSurface  from  Adaptor3d; 
      LeftBot, RightTop : out Pnt2d from gp) 
     returns  Boolean       
     is  static  private;  

     LocatePart_Offset(me; UV : Pnt2d  from  gp; DUV : Vec2d from gp; 
    	S  :  HSurface  from  Adaptor3d; 
      LeftBot, RightTop : out Pnt2d from gp)  
     returns  Boolean       
     is  static  private;  

     FindBounds(me;  Arr  :  Array1OfReal  from  TColStd; 
    	    	  XYComp : Real  from  Standard; 
    	    	 DUVComp : Real  from  Standard;  
    	            Bnd1 :  out  Integer from  Standard; 
		    Bnd2 :  out  Integer from  Standard; 
	       DerIsNull :  out  Boolean  from  Standard) 
        ---Purpose: Extracts the numbers of knots which equal 
	--  the point and checks derivative components 
	--  by  zero equivalence.   		     
     is  static  private;  
      
    

fields

  mySurface  : HSurface  from Adaptor3d;
  myCurve    : HCurve2d  from Adaptor2d;
    
  myType     : CurveType from GeomAbs;
  myCirc     : Circ      from gp;
  myLin      : Lin       from gp;

  myFirstSurf  :  HSurface  from  Adaptor3d; 
  myLastSurf   :  HSurface  from  Adaptor3d;  
  
  myIntervals  : HSequenceOfReal from TColStd;
  myIntCont    : Shape from GeomAbs;

end CurveOnSurface;




