-- Created on: 1993-03-02
-- Created by: Philippe DAUTRY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class OffsetSurface from PGeom inherits Surface from PGeom

        ---Purpose : This class implements  the basis services for  an
        --         offset surface in 3D space.
        --         

uses Surface from PGeom

is


  Create returns OffsetSurface from PGeom;
    ---Purpose: Creates an OffsetSurface with default values.
    	---Level: Internal 


  Create (
    	    aBasisSurface : Surface from PGeom;
    	    aOffsetValue : Real from Standard)
     returns OffsetSurface from PGeom;
        ---Purpose :  <aBasisSurface>    is  the   basis      surface,
        --         <aOffsetValue> is the distance between <me> and the
        --         basis  surface at any  point.    <aOffsetDirection>
        --         defines  the  fixed  reference  direction   (offset
        --         direction).
    	---Level: Internal 


  BasisSurface (me : mutable; aBasisSurface : Surface from PGeom);
	---Purpose: Set the field basisSurface with <aBasisSurface>.
    	---Level: Internal 
      

  BasisSurface (me) returns Surface from PGeom;
        ---Purpose : The basis surface can be an offset surface.
    	---Level: Internal 


  OffsetValue (me : mutable; aOffsetValue : Real from Standard);
        ---Purpose : Set the field offsetValue with <aOffsetValue>.
    	---Level: Internal 


  OffsetValue (me) returns Real from Standard;
        ---Purpose : Returns the value of the field offsetValue.
    	---Level: Internal 


fields

  basisSurface : Surface from PGeom;
  offsetValue  : Real from Standard;

end;
