-- Created on: 1998-06-30
-- Created by: Christian CAILLET
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class RepresentationRelationshipWithTransformation  from StepRepr
    inherits ShapeRepresentationRelationship

    -- in principle, inherits RepresentationRelationship
    -- But <Shape>... only adds a constraint on a field, this allows to
    -- simplify the multiple inheritance between ShapeRR and RRWithTransf...

uses
     HAsciiString from TCollection,
     Representation from StepRepr,
     Transformation from StepRepr

is

    Create returns RepresentationRelationshipWithTransformation;

    Init (me : mutable;
              aName : HAsciiString from TCollection;
              aDescription : HAsciiString from TCollection;
              aRep1 : Representation from StepRepr;
              aRep2 : Representation from StepRepr;
	      aTransf : Transformation);

    TransformationOperator (me) returns Transformation;
    SetTransformationOperator (me : mutable; aTrans : Transformation);

fields

    theTrans : Transformation;

end RepresentationRelationshipWithTransformation;
