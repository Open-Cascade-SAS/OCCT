-- Created on: 1991-01-10
-- Created by: Arnaud BOUZY
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class PolyExpression from Expr

inherits GeneralExpression from Expr

uses SequenceOfGeneralExpression from Expr,
    NamedUnknown from Expr

raises OutOfRange from Standard, 
    NumericError from Standard,
    InvalidOperand from Expr

is

    Initialize;
    ---Purpose: initialize an empty list of operands.
    
    NbOperands(me)
    ---Purpose: returns the number of operands contained in <me>
    ---Level : Internal
    returns Integer
    is static;

    Operand(me; index : Integer)
    ---Purpose: Returns the <index>-th operand used in <me>.
    --          An exception is raised if index is out of range
    ---C++: inline
    ---C++: return const &
    ---Level : Internal
    returns any GeneralExpression
    raises OutOfRange
    is static;

    SetOperand(me : mutable; exp : GeneralExpression; index : Integer)
    ---Purpose: Sets the <index>-th operand used in <me>.
    --          An exception is raised if <index> is out of range
    --          Raises InvalidOperand if <exp> contains <me>.
    ---Level : Internal
    raises OutOfRange,InvalidOperand
    is static;

    AddOperand(me : mutable; exp : GeneralExpression)
    ---Purpose: Adds an operand to the list of <me>.
    ---Level : Internal
    is static protected;

    RemoveOperand(me : mutable; index : Integer)
    ---Purpose: Remove the operand denoted by <index> from the list of 
    --          <me>. 
    --          Raises exception if <index> is out of range or if 
    --          removing operand intend to leave only one or no 
    --          operand. 
    ---Level : Internal
    raises OutOfRange
    is static protected;

    NbSubExpressions(me)
    ---Purpose: returns the number of sub-expressions contained
    --          in <me> ( >= 2)
    returns Integer
    is static;

    SubExpression(me; I : Integer)
    ---Purpose: Returns the sub-expression denoted by <I> in <me>
    --          Raises OutOfRange if <I> > NbSubExpressions(me)
    ---C++: return const &
    returns any GeneralExpression
    raises OutOfRange
    is static;

    ContainsUnknowns(me) 
    ---Purpose: Does <me> contains NamedUnknown ?
    returns Boolean
    is static;

    Contains(me; exp : GeneralExpression)
    ---Purpose: Tests if <exp> is contained in <me>.
    returns Boolean
    is static;

    Replace(me : mutable ; var : NamedUnknown ; with : GeneralExpression)
    ---Purpose: Replaces all occurences of <var> with <with> in <me>
    --          Raises InvalidOperand if <with> contains <me>.
    raises InvalidOperand
    is static;
    
    Simplified(me) 
    ---Purpose: Returns a GeneralExpression after replacement of
    --          NamedUnknowns by an associated expression and after
    --          values computation.
    returns any GeneralExpression
    raises NumericError;
    
fields

    myOperands  : SequenceOfGeneralExpression;

end PolyExpression;
