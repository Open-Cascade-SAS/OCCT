-- Created on: 1993-02-22
-- Created by: Philippe DAUTRY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Axis1Placement from PGeom inherits AxisPlacement from PGeom

	---Purpose : This class describes an axis  one placement built
	--         with a point and a direction.
	--          

uses Ax1 from gp

is


  Create returns mutable Axis1Placement from PGeom;
        --- Purpose : Creates an Axis1Placement with Ax1 default value.
    	---Level: Internal 

  Create (aAxis : Ax1 from gp) returns mutable Axis1Placement from PGeom;
        --- Purpose : Creates an Axis1Placement with <aAxis>.
    	---Level: Internal 


end;


