-- Created on: 2000-03-01
-- Created by: Denis PASCAL
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class DrawDocument from DDocStd inherits Data from DDF

	---Purpose: draw variable for TDocStd_Document.
	--          ==================================

uses Document    from TDocStd,
     Drawable3D  from Draw,
     Interpretor from Draw,
     Display     from Draw

is 


    Find (myclass; Doc : Document from TDocStd)
    returns DrawDocument from DDocStd;

    Create (Doc : Document from TDocStd)
    returns mutable DrawDocument from DDocStd;

    GetDocument(me) returns Document from TDocStd;

    DrawOn (me; dis : in out Display from Draw);
    
    Copy (me) 
    returns mutable Drawable3D from Draw
    is redefined;
	
    Dump (me; S : in out OStream) 
    is redefined;
    
    Whatis (me; I : in out Interpretor from Draw)
    is redefined;

fields

    myDocument : Document from TDocStd;

end DrawDocument;
