-- Created on: 1994-11-07
-- Created by: Christian CAILLET
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class CheckCounter  from IFSelect  inherits SignatureList

    ---Purpose : A CheckCounter allows to see a CheckList (i.e. CheckIterator)
    --           not per entity, its messages, but per message, the entities
    --           attached (count and list). Because many messages can be
    --           repeated if they are due to systematic errors

uses CheckIterator, InterfaceModel, SignText from MoniTool

is

    Create (withlist : Boolean = Standard_False) returns mutable CheckCounter;
    ---Purpose : Creates a CheckCounter, empty ready to work

    SetSignature (me : mutable; sign : SignText);
    ---Purpose : Sets a specific signature
    --           Else, the current SignType (in the model) is used

    Signature    (me) returns SignText;
    ---Purpose : Returns the Signature;
 
    Analyse (me : mutable;
    	 list  : CheckIterator;
    	 model : InterfaceModel;
	 original  : Boolean = Standard_False;
	 failsonly : Boolean = Standard_False);
    ---Purpose : Analyses a CheckIterator according a Model (which detains the
    --           entities for which the CheckIterator has messages), i.e.
    --           counts messages for entities
    --           If <original> is True, does not consider final messages but
    --             those before interpretation (such as inserting variables :
    --             integers, reals, strings)
    --           If <failsonly> is True, only Fails are considered
    --           Remark : global messages are recorded with a Null entity

fields

    thesign : SignText;  -- optional

end CheckCounter;
