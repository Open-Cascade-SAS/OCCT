-- Created on: 1997-07-28
-- Created by: Pierre CHALAMET
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

class Texture2Dmanual from Graphic3d

inherits Texture2D from Graphic3d

  ---Purpose: This class defined a manual texture 2D
  -- facets MUST define texture coordinate
  -- if you want to see somethings on.

uses

  NameOfTexture2D from Graphic3d,
  AsciiString     from TCollection

is

  Create (theFileName : AsciiString from TCollection) returns mutable Texture2Dmanual from Graphic3d;
  ---Purpose: Creates a texture from a file

  Create (theNOT : NameOfTexture2D from Graphic3d) returns mutable Texture2Dmanual from Graphic3d;
  ---Purpose: Creates a texture from a predefined texture name set.

end Texture2Dmanual;
