-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class OrientedEdge from StepShape 

inherits Edge from StepShape 

uses

	Boolean from Standard, 
	Vertex from StepShape, 
	HAsciiString from TCollection
is

	Create returns mutable OrientedEdge;
	---Purpose: Returns a OrientedEdge
	

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aEdgeElement : mutable Edge from StepShape;
	      aOrientation : Boolean from Standard) is virtual;

	-- Specific Methods for Field Data Access --

	SetEdgeElement(me : mutable; aEdgeElement : mutable Edge);
	EdgeElement (me) returns mutable Edge;
	SetOrientation(me : mutable; aOrientation : Boolean);
	Orientation (me) returns Boolean;
	SetEdgeStart(me : mutable; aEdgeStart : mutable Vertex) is redefined;
	EdgeStart (me) returns mutable Vertex is redefined;
	SetEdgeEnd(me : mutable; aEdgeEnd : mutable Vertex) is redefined;
	EdgeEnd (me) returns mutable Vertex is redefined;

fields

	edgeElement : Edge from StepShape;
	orientation : Boolean from Standard;

 -- 
 -- NB : field <edge_start> inherited from classe <edge> is redeclared.
 --      it shall appears in a physical file as a *.
 --

 -- 
 -- NB : field <edge_end> inherited from classe <edge> is redeclared.
 --      it shall appears in a physical file as a *.
 --

end OrientedEdge;
