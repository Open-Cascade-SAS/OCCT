-- Created on: 1996-07-01
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

private class HBuilder from LocOpe 

	---Purpose: 

inherits HBuilder from TopOpeBRepBuild

uses BuildTool from TopOpeBRepDS

is

    Create(BT: BuildTool from TopOpeBRepDS)
    
	---C++: inline
    	returns mutable HBuilder from LocOpe;
    

    Classify(me)
    
	---C++: inline
    	returns Boolean from Standard
	is static;
    

    Classify(me: mutable; B: Boolean from Standard)
    
	---C++: inline
    	is static;


end HBuilder;
