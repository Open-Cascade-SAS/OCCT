-- Created on: 1994-03-30
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class SITopolTool from IntStart 

	---Purpose: template class for a topological tool.
	--          This tool is linked with the surface on which
	--          the classification has to be made.


inherits TShared from MMgt

uses State from TopAbs,
     Pnt2d from gp


is

    Classify(me: mutable; P: Pnt2d from gp; Tol: Real from Standard)
    
    	returns State from TopAbs
	is deferred;


end SITopolTool;
