-- Created on: 1999-12-20
-- Created by: data exchange team
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class MakeTriangulation from ShapeConstruct  inherits MakeShape from BRepBuilderAPI

	---Purpose: 

uses

    Array1OfPnt from TColgp,
    Wire from TopoDS

is

    Create (pnts : Array1OfPnt from TColgp; prec : Real = 0.0)
    returns MakeTriangulation from ShapeConstruct;

    Create (wire : Wire from TopoDS; prec : Real = 0.0)
    returns MakeTriangulation from ShapeConstruct;

    Build (me : in out) is redefined;

    IsDone (me) returns Boolean is redefined;

    Triangulate (me : in out; wire : Wire from TopoDS) is private;

    AddFacet (me : in out; wire : Wire from TopoDS) is private;

fields

    myPrecision : Real from Standard;
    myWire      : Wire from TopoDS;

end MakeTriangulation;
