
-- File:	Graphic2d_Circle.cdl
-- Created:	Tue Jun 22 16:36:51 1993
-- Author:	Jean Louis FRENKEL, Gerard GRAS
--		<jlf@stylox>
-- Modified: TCL G002, 07-08-00, new inquire methods Center, Radius, FirstAngle, SecondAngle
--                               new methods SetRadius, SetCenter, SetAngles

---Copyright:	 Matra Datavision 1993

class Circle from Graphic2d inherits Line from Graphic2d

	---Purpose: Constructs a primitive Circle

	
uses
	Drawer		from Graphic2d,
	GraphicObject	from Graphic2d,
	Length		from Quantity,
	PlaneAngle	from Quantity,
	FStream		from Aspect,
	IFStream	from Aspect

raises
	CircleDefinitionError	from Graphic2d

is
	-------------------------
	-- Category: Constructors
	-------------------------

	Create (aGraphicObject: GraphicObject from Graphic2d;
		X, Y: Length from Quantity;
		Radius: Length from Quantity)
	returns mutable Circle from Graphic2d
	---Level: Public
	---Purpose: Creates a complete circle.
	--	    The center is <X>, <Y>.
	--	    The radius is <Radius>.
	--  Warning: Raises CircleDefinitionError if the
	--          radius is null.
	raises CircleDefinitionError from Graphic2d;

	Create (aGraphicObject: GraphicObject from Graphic2d;
		X, Y: Length from Quantity;
		Radius: Length from Quantity;
		Alpha, Beta: PlaneAngle from Quantity)
	returns mutable Circle from Graphic2d
	---Level: Public
	---Purpose: Creates an arc.
	--	    The center is <X>, <Y>.
	--	    The radius is <Radius>.
	--	    Angles are measured counterclockwise with 0 radian
	--	    at 3 o'clock.
	--  Warning: Raises CircleDefinitionError if the
	--          radius is null.
	raises CircleDefinitionError from Graphic2d;

	----------------------------
	-- Category: Inquire methods
	----------------------------

	Center( me; X, Y: out Length from Quantity );  
	---Level: Public
	---Purpose: returns the coordinates of center of the circle
	
	Radius( me ) returns Length from Quantity;
	---Level: Public
	---Purpose: returns the radius of this circle
	
	FirstAngle( me ) returns PlaneAngle from Quantity;
	---Level: Public
	---Purpose: returns the first angle of the arc
	
	SecondAngle( me ) returns PlaneAngle from Quantity;
	---Level: Public
	---Purpose: returns the second angle of the arc
	

	--------------------------------------------------------
	-- Category: Methods for the definition of the circle's properties
	--------------------------------------------------------

	SetCenter( me: mutable; X, Y: Length from Quantity );  
	---Level: Public
	---Purpose: defines the coordinates of center of the circle
	
	SetRadius( me: mutable; theR: Length from Quantity );
	---Level: Public
	---Purpose: defines the radius of this circle
	
	SetAngles( me: mutable; Alpha, Beta: PlaneAngle from Quantity );
	---Level: Public
	---Purpose: defines the angles of the arc

	--------------------------
	-- Category: Draw and Pick
	--------------------------

	Draw (me : mutable; aDrawer: Drawer from Graphic2d)
	is static protected;
	---Level: Internal
	---Purpose: Draws the circle <me>.

	DrawElement( me : mutable; aDrawer: Drawer from Graphic2d;
		 anIndex: Integer from Standard)
	is redefined protected;
	---Level: Internal
	---Purpose: Draws element <anIndex> of the circle <me>.

	DrawVertex( me : mutable; aDrawer: Drawer from Graphic2d;
		anIndex: Integer from Standard)
	is redefined protected;
	---Level: Internal
	---Purpose: Draws vertex <anIndex> of the circle <me>.

	Pick (me : mutable; X, Y: ShortReal from Standard;
		aPrecision: ShortReal from Standard;
		aDrawer: Drawer from Graphic2d)
	returns Boolean from Standard is static protected;
	---Level: Internal
	---Purpose: Returns Standard_True if the circle <me> is picked,
	--	    Standard_False if not.

	DoMinMax( me: mutable ) is private;

	----------------------------------------------------------------------

	Save( me; aFStream: in out FStream from Aspect ) is virtual;
	Retrieve( myclass; anIFStream: in out IFStream from Aspect;
		aGraphicObject: GraphicObject from Graphic2d );

fields

	myX:		ShortReal from Standard;
	myY:		ShortReal from Standard;
	myRadius:	ShortReal from Standard;
	myFirstAngle:	ShortReal from Standard;
	mySecondAngle:	ShortReal from Standard;
	myisArc:	Boolean from Standard;

end Circle from Graphic2d;
