-- Created on: 1992-12-02
-- Created by: Isabelle GRIGNON
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class VelGProps from GProp  inherits GProps

        --- Purpose :
        --  Computes the global properties of a geometric solid 
        --  (3D closed region of space) 
        --  The solid can be elementary(definition in the gp package) 


uses   	Cone     from gp,
	Cylinder from gp,
        Pnt      from gp,
	Sphere   from gp,
	Torus    from gp


is


  Create returns VelGProps;

  
  Create (S : Cylinder; Alpha1, Alpha2, Z1, Z2 : Real; VLocation : Pnt)   
     returns VelGProps;


  Create (S : Cone; Alpha1, Alpha2, Z1, Z2 : Real; VLocation : Pnt) 
     returns VelGProps;


  Create (S : Sphere; Teta1, Teta2, Alpha1, Alpha2 : Real; VLocation : Pnt)
     returns VelGProps;


  Create (S : Torus; Teta1, Teta2, Alpha1, Alpha2 : Real; VLocation : Pnt)
     returns VelGProps;


  SetLocation(me : in out ;VLocation :Pnt);
  
  Perform(me : in out;S : Cylinder; Alpha1, Alpha2, Z1, Z2 : Real);

  Perform(me : in out;S : Cone; Alpha1, Alpha2, Z1, Z2 : Real);

  Perform(me : in out;S : Sphere; Teta1, Teta2, Alpha1, Alpha2 : Real);

  Perform(me : in out;S : Torus; Teta1, Teta2, Alpha1, Alpha2 : Real);

end VelGProps;

