-- File:        BSplineCurveWithKnotsAndRationalBSplineCurve.cdl
-- Created:     Mon Dec  4 12:02:33 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWBSplineCurveWithKnotsAndRationalBSplineCurve from RWStepGeom

	---Purpose : Read & Write Module for BSplineCurveWithKnotsAndRationalBSplineCurve
	--           Check added by CKY , 7-OCT-1996

uses Check from Interface, ShareTool from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     BSplineCurveWithKnotsAndRationalBSplineCurve from StepGeom,
     EntityIterator from Interface

is

	Create returns RWBSplineCurveWithKnotsAndRationalBSplineCurve;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable BSplineCurveWithKnotsAndRationalBSplineCurve from StepGeom);

	WriteStep (me; SW : in out StepWriter; ent : BSplineCurveWithKnotsAndRationalBSplineCurve from StepGeom);

	Share(me; ent : BSplineCurveWithKnotsAndRationalBSplineCurve from StepGeom; iter : in out EntityIterator);

    	Check(me; ent : BSplineCurveWithKnotsAndRationalBSplineCurve from StepGeom; shares : ShareTool; ach : in out Check);

end RWBSplineCurveWithKnotsAndRationalBSplineCurve;
