-- Created on: 2000-10-31
-- Created by: Vladislav ROMASHKO
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

class Limitation from QANewBRepNaming inherits BooleanOperationFeat from QANewBRepNaming

uses

    Label from TDF, 
    MakeShape from BRepBuilderAPI,
    Limitation from QANewModTopOpe

is
 
    Create returns Limitation from QANewBRepNaming;

    Create(ResultLabel : Label from TDF) 
    returns Limitation from QANewBRepNaming;

    Load (me; MakeShape : in out Limitation from QANewModTopOpe); 
     
    LoadContent(me; MakeShape : in out Limitation from QANewModTopOpe)
    ---Purpose: Loads the content of the result.
    is protected;

    LoadResult(me; MakeShape : in out Limitation from QANewModTopOpe)
    ---Purpose: Loads the result.
    is protected;

    LoadDegenerated(me; MakeShape : in out Limitation from QANewModTopOpe)
    ---Purpose: Loads the deletion of the degenerated edges.
    is protected;    


    LoadWire(me; MakeShape : in out Limitation from QANewModTopOpe)
    ---Purpose: A default implementation for naming of a wire as an object of
    --          a boolean operation.
    is protected;

    LoadShell(me; MakeShape : in out Limitation from QANewModTopOpe)
    ---Purpose: A default implementation for naming of a shell as an object of
    --          a boolean operation.
    is protected;

end Limitation;
