-- Created on: 1998-06-03
-- Created by: data exchange team
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Surface from ShapeCustom 

    ---Purpose: Converts a surface to the analitical form with given 
    --          precision. Conversion is done only the surface is bspline
    --          of bezier and this can be approximed by some analytical
    --          surface with that precision.

uses
    Surface from Geom

is

    Create returns Surface from ShapeCustom;
    
    Create (S: Surface from Geom) returns Surface from ShapeCustom;

    Init (me: in out; S: Surface from Geom);

    Gap (me) returns Real;
    ---C++: inline
    	---Purpose: Returns maximal deviation of converted surface from the original 
	--          one computed by last call to ConvertToAnalytical

    ConvertToAnalytical (me: in out; tol: Real;
    	    	    	    	     substitute: Boolean)
    returns Surface from Geom;
    	---Purpose: Tries to convert the Surface to an Analytic form
    	--          Returns the result
    	--          Works only if the Surface is BSpline or Bezier.
    	--          Else, or in case of failure, returns a Null Handle
    	--
    	--          If <substitute> is True, the new surface replaces the actual
    	--          one in <me>
    	--
    	--          It works by analysing the case which can apply, creating the
    	--          corresponding analytic surface, then checking coincidence
    	--  Warning: Parameter laws are not kept, hence PCurves should be redone
	
    ConvertToPeriodic (me: in out; substitute: Boolean; preci: Real = -1)
    returns Surface from Geom;
        ---Purpose: Tries to convert the Surface to the Periodic form
    	--          Returns the resulting surface
    	--          Works only if the Surface is BSpline and is closed with 
        --          Precision::Confusion()
    	--          Else, or in case of failure, returns a Null Handle
fields

    mySurf: Surface from Geom;
    myGap : Real; -- maximal deviation of converted surface from original one

end Surface;
