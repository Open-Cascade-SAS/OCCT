-- Created by: Tanya COOL
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class AspectFramedText from Prs2d inherits AspectRoot from Prs2d

---Purpose: defines the attributes when drawing a framed text Presentation.

uses 
    
	 NameOfColor from Quantity,
	 WidthOfLine from Aspect,
	 TypeOfFont from Aspect

is
 
    Create(  ColorInd:        NameOfColor from Quantity;
             FrameColorInd:   NameOfColor from Quantity;
             FrameWidthInd:   WidthOfLine from Aspect;
             FontInd:         TypeOfFont from Aspect;
             aSlant:          ShortReal from Standard;
             aHScale,aWScale: ShortReal from Standard;
             isUnderlined:    Boolean from Standard )
	 	   returns mutable AspectFramedText from Prs2d;

    SetColorOfText( me: mutable;  aColor:        NameOfColor from Quantity); 
    SetFrameColor ( me: mutable;  aFrameColor:   NameOfColor from Quantity);  
    SetFrameWidth ( me: mutable;  aFrameWidth:   WidthOfLine from Aspect); 
    SetFontOfText ( me: mutable;  aFont:         TypeOfFont from Aspect);  
    SetSlant      ( me: mutable;  aSlant:        ShortReal  from  Standard); 
    SetHScale     ( me: mutable;  aHScale:       ShortReal  from  Standard); 
    SetWScale     ( me: mutable;  aWScale:       ShortReal  from  Standard);  
    SetUnderlined ( me: mutable;  anIsUnderlined:Boolean from  Standard); 

    Values( me;
	      aColorInd:        out NameOfColor from Quantity;
            aFrameColorInd:   out NameOfColor from Quantity;
            aFrameWidthInd:   out WidthOfLine from Aspect;
            aFontInd:         out TypeOfFont from Aspect;
            aSlant:           out ShortReal from Standard;
            aHScale,aWScale:  out ShortReal from Standard;
            isUnderlined:     out Boolean from Standard );
    
fields

    myColor	          : NameOfColor from Quantity;
    myFrameColor      : NameOfColor from Quantity;
    myFont	          : TypeOfFont from Aspect;
    myFrameWidth      : WidthOfLine from Aspect;
    mySlant           : ShortReal from Standard;
    myHScale          : ShortReal from Standard;
    myWScale          : ShortReal from Standard;
    myIsUnderlined    : Boolean from Standard;
 
end AspectFramedText from Prs2d;
