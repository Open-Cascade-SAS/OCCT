-- Created on: 2004-03-05
-- Created by: Mikhail KUZMITCHEV
-- Copyright (c) 2004-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package QANCollection

uses
    Draw,
    TCollection, 
    TColStd,
    gp

is
    class  ListOfPnt   instantiates  List  from  TCollection    (Pnt  from  gp);
    class  StackOfPnt  instantiates  Stack from  TCollection    (Pnt  from  gp);
    class  SListOfPnt  instantiates  SList from  TCollection    (Pnt  from  gp);
    class  DataMapOfRealPnt instantiates DataMap from TCollection  
                                        (Real from Standard, 
                                         Pnt from gp, 
                                         MapRealHasher from TColStd);
    class  IndexedDataMapOfRealPnt instantiates IndexedDataMap from TCollection
                                        (Real from Standard, 
                                         Pnt from gp, 
                                         MapRealHasher from TColStd);
    class  DoubleMapOfRealInteger instantiates DoubleMap from TCollection  
                                        (Real from Standard, 
                                         Integer from Standard, 
                                         MapRealHasher from TColStd, 
                                         MapIntegerHasher from TColStd);


---    HashCode (thePnt   : Pnt from gp;
---              theUpper : Integer from Standard)
---    returns Integer from Standard;
    
---    IsEqual (thePnt1   : Pnt from gp;
---             thePnt2   : Pnt from gp)
---    returns Boolean from Standard;
    
    Commands(DI : in out Interpretor from Draw);
    Commands1(DI : in out Interpretor from Draw);
    Commands2(DI : in out Interpretor from Draw);
    Commands3(DI : in out Interpretor from Draw);
    Commands4(DI : in out Interpretor from Draw);

end;
