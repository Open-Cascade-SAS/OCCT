-- Created on: 1992-09-29
-- Created by: Didier PIFFAULT
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



generic class InterferencePolygon3d from Intf 
    (Polygon3d1 as any;
     ToolPolygon3d1 as any;         -- as ToolPolygon(Pnt,Polygon3d1,Box)
     Polygon3d2 as any;
     ToolPolygon3d2 as any)         -- as ToolPolygon(Pnt,Polygon3d2,Box)
    inherits Interference from Intf
    	
	---Purpose: Computes the  interference between two polygons  or the
	--          self interference of a polygon in 3 dimensions .  In 3
	--          dimensions the result can be  a common perpendicular ,
	--          an  orthogonal  projection or  a  real  intersections.
	--          There  are two  different  instantiation arguments  to
	--          authorize an interference  between two  polygons  from
	--          differents origin.  Ex :  to intersect a curve polygon
	--          with an  algorithmic   curve   from numerical  walking
	--          between two surfaces.

uses    Pnt from gp,
    	SectionPoint      from Intf,
    	SeqOfSectionPoint from Intf,
    	SectionLine       from Intf,
    	SeqOfSectionLine  from Intf

raises  OutOfRange from Standard


is
-- Interface :

    Create          returns InterferencePolygon3d from Intf;
    ---Purpose: Constructs an empty interference of 3d Polygon.


    Create         (Obje1 : in Polygon3d1 ;Obje2 : in Polygon3d2) 
    	            returns InterferencePolygon3d from Intf;
    ---Purpose: Constructs and computes an interference between two Polygons.


    Create         (Obje : in Polygon3d1) 
    	            returns InterferencePolygon3d from Intf;
    ---Purpose: Constructs and computes the self interference of a Polygon.


    Perform        (me   : in out;
    	    	    Obje1 : in Polygon3d1 ;Obje2 : in Polygon3d2);
    ---Purpose: Computes an interference between two Polygons.


    Perform        (me   : in out;
    	    	    Obje : in Polygon3d1);
    ---Purpose: Computes the auto interference of a Polygon.


    NbResults      (me)
    	    	    returns Integer is static;
    ---Purpose: Gives  the number  of common  Perpendiculars or orthogonal
    --          projections between the two polygons.

    ResultLine     (me;
    	    	    Index      : in Integer)
    	    	    returns SectionLine from Intf
    	    	    raises OutOfRange from Standard
    	    	    is static;
    ---Purpose: Gives the  segment of address  <Index> in the interference
    --          representing    the     perpendicular  or the   orthogonal
    --          projection .
    --          
    ---C++: return const &


    ResultValue    (me;
    	    	    Index      : in Integer)
    	    	    returns Real from Standard
    	    	    raises OutOfRange from Standard
    	    	    is static;
    ---Purpose: Gives the distance between the two polygons 


    MinimalDistance(me)
    	    	    returns Real from Standard
    	    	    is static;
    ---Purpose: Gives   the distance  between  the  two  polygon3d at  the
    --          perpendicular or projection of minimal length.


    MinimalResult  (me)
    	    	    returns Integer from Standard
    	    	    is static;
    ---Purpose: Give the  perpendicular or projection  of minimal  length.
    --          WARNING : if there  are points of intersection the minimal
    --          result is one of them and this function is unusuable.


-- Implementation :

    Interference   (me         : in out;
    	    	    Obje1      : in Polygon3d1;
     	    	    Obje2      : in Polygon3d2)
    	    	    is private;

    Interference   (me         : in out;
    	    	    Obje       : in Polygon3d1)
    	    	    is private;

    CommonPerpen   (me         : in out;
		    BegO : in Pnt from gp;
		    EndO : in Pnt from gp;
		    BegT : in Pnt from gp;
		    EndT : in Pnt from gp)
    	    	    is private;
    ---Purpose: Computes   the common  perpendicular   between the two
    --          segments <BegO><EndO> and <BegT><EndT>.

    Projections    (me         : in out;
		    BegO : in Pnt from gp;
		    EndO : in Pnt from gp;
		    BegT : in Pnt from gp;
		    EndT : in Pnt from gp)
    	    	    is private;
    ---Purpose: Computes  the    different  orthogonal projections  between
    --          segment <BegO><EndO> and  points <BegT>,<EndT> and segment
    --          <BegT><EndT> and points <BegO>,<EndO>.


fields  IndexMin             : Integer from Standard;
    	MinimalDist          : Real from Standard;
        iObje1, iObje2       : Integer from Standard;
        beginOfNotClosedFirst: Boolean from Standard;
        beginOfNotClosedSecon: Boolean from Standard;


end InterferencePolygon3d;
