-- Created on: 1994-06-01
-- Created by: Christian CAILLET
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class FloatFormat  from StepSelect    inherits FileModifier  from StepSelect

    ---Purpose : This class gives control out format for floatting values :
    --           ZeroSuppress or no, Main Format, Format in Range (for values
    --           around 1.), as StepWriter allows to manage it.
    --           Formats are given under C-printf form

uses CString, AsciiString from TCollection, HSequenceOfInteger from TColStd,
     CheckIterator, StepWriter , ContextWrite

is

    Create returns mutable FloatFormat;
    ---Purpose : Creates a new FloatFormat, with standard options :
    --           ZeroSuppress, Main Format = %E,
    --           Format between 0.001 and 1000. = %f

    SetDefault (me : mutable; digits : Integer = 0);
    ---Purpose : Sets FloatFormat to default value (see Create) but if <digits>
    --           is given positive, it commands Formats (main and range) to
    --           ensure <digits> significant digits to be displayed

    SetZeroSuppress (me : mutable; mode : Boolean);
    ---Purpose : Sets ZeroSuppress mode to a new value

    SetFormat (me : mutable; format : CString = "%E");
    ---Purpose : Sets Main Format to a new value
    --           Remark : SetFormat, SetZeroSuppress and SetFormatForRange are
    --           independant

    SetFormatForRange (me : mutable; format : CString = "%f";
    	    	       Rmin : Real = 0.1; Rmax : Real = 1000.0);
    ---Purpose : Sets Format for Range to a new value with its range of
    --           application.
    --           To cancel it, give format as "" (empty string)
    --           Remark that if the condition (0. < Rmin < Rmax)  is not
    --           verified, this secondary format will be ignored.
    --           Moreover, this secondary format is intended to be used in a
    --           range around 1.


    Format (me; zerosup  : out Boolean;
    	    	mainform : out AsciiString from TCollection;
		hasrange : out Boolean;
		forminrange : out AsciiString from TCollection;
		rangemin, rangemax : out Real);
    ---Purpose : Returns all recorded parameters :
    --           zerosup  : ZeroSuppress status
    --           mainform : Main Format (which applies out of the range, or
    --                       for every real if no range is set)
    --           hasrange : True if a FormatInRange is set, False else
    --                      (following parameters do not apply if it is False)
    --           forminrange : Secondary Format (it applies inside the range)
    --           rangemin, rangemax : the range in which the secondary format
    --                                applies


    Perform (me; ctx : in out ContextWrite;
    	     writer  : in out StepWriter);
    ---Purpose : Sets the Floatting Formats of StepWriter to the recorded
    --           parameters

    Label (me) returns AsciiString from TCollection;
    ---Purpose : Returns specific Label : for instance,
    --           "Float Format [ZeroSuppress] %E [, in range R1-R2 %f]"

fields

    thezerosup   : Boolean;
    themainform  : AsciiString from TCollection;
    theformrange : AsciiString from TCollection;
    therangemin  : Real;
    therangemax  : Real;

end FloatFormat;

