-- Created on: 1992-02-18
-- Created by: Christophe MARION
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class PolyAlgo from HLRAlgo inherits TShared from MMgt

	---Purpose: to remove Hidden lines on Triangulations.

uses
    Address                    from Standard,
    Boolean                    from Standard,
    Integer                    from Standard,
    Real                       from Standard,
    HArray1OfTransient         from TColStd,
    Array1OfTransient          from TColStd,
    ListIteratorOfListOfBPoint from HLRAlgo,
    EdgeStatus                 from HLRAlgo
    
is
    Create
    returns mutable PolyAlgo from HLRAlgo;
    
    Init(me : mutable; HShell : HArray1OfTransient from TColStd)
    is static;

    PolyShell(me) returns Array1OfTransient from TColStd
	---C++: return &
	---C++: inline
    is static;
    
    Clear(me : mutable)
    is static;
    
    Update(me : mutable)
	---Purpose: Prepare all the data to process the algo.
    is static;
    
    InitHide(me : mutable)
	---C++: inline
    is static;

    MoreHide(me) returns Boolean from Standard
	---C++: inline
    is static;

    NextHide(me : mutable)
    is static;

    Hide(me : mutable; Coordinates : out Address    from Standard;
                       status      : out EdgeStatus from HLRAlgo;
		       Index       : out Integer    from Standard;
                       reg1,regn   : out Boolean    from Standard;
                       outl,intl   : out Boolean    from Standard)
	---Purpose: process hiding between <Pt1> and <Pt2>.
    is static;
    
    InitShow(me : mutable)
	---C++: inline
    is static;

    MoreShow(me) returns Boolean from Standard
	---C++: inline
    is static;

    NextShow(me : mutable)
    is static;

    Show(me : mutable; Coordinates : out Address from Standard;
		       Index       : out Integer from Standard;
                       reg1,regn   : out Boolean from Standard;
                       outl,intl   : out Boolean from Standard)
	---Purpose: process hiding between <Pt1> and <Pt2>.
    is static;
    
fields
    myHShell    : HArray1OfTransient         from TColStd;
    myRealPtr   : Real                       from Standard[10];
    mySegListIt : ListIteratorOfListOfBPoint from HLRAlgo;
    myNbrShell  : Integer                    from Standard;
    myCurShell  : Integer                    from Standard;
    myFound     : Boolean                    from Standard;

end PolyAlgo;
