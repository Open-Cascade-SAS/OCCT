-- Created on: 1991-05-14
-- Created by: Laurent PAINNOT
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class Jacobi from math
    	---Purpose:
      	-- This class implements the Jacobi method to find the eigenvalues and
      	-- the eigenvectors of a real symmetric square matrix.
      	-- A sort of eigenvalues is done.

uses Vector from math, 
     Matrix from math,
     OStream from Standard

raises NotDone from StdFail

is

      Create(A: Matrix)
      	---Purpose:
      	-- Given a Real n X n matrix A, this constructor computes all its
      	-- eigenvalues and eigenvectors using the Jacobi method.
      	-- The exception NotSquare is raised if the matrix is not square.
      	-- No verification that the matrix A is really symmetric is done.
      
      returns Jacobi;
      

    IsDone(me)
    	---Purpose: Returns true if the computations are successful, otherwise returns false.
        ---C++: inline
    returns Boolean
    is static;
    

    Values(me)
    	---Purpose: Returns the eigenvalues vector.
        -- Exception NotDone is raised if calculation is not done successfully.
    	---C++: inline
    	---C++: return const&
    returns Vector
    raises NotDone
    is static;
    
    
    Value(me; Num: Integer)
    	---Purpose: returns the eigenvalue number Num.
        -- Eigenvalues are in the range (1..n).
        -- Exception NotDone is raised if calculation is not done successfully.
        ---C++: inline
    returns Real
    raises NotDone
    is static;
    
    
    Vectors(me)
    	---Purpose: returns the eigenvectors matrix.
        -- Exception NotDone is raised if calculation is not done successfully.
    	---C++: inline
    	---C++: return const&
    returns Matrix
    raises NotDone
    is static;
    
    
    Vector(me; Num: Integer; V : out Vector)
    	---Purpose: Returns the eigenvector V of number Num.
        -- Eigenvectors are in the range (1..n).    
        -- Exception NotDone is raised if calculation is not done successfully.
    	---C++: inline
    raises NotDone
    is static;



    Dump(me; o: in out OStream)
    	---Purpose: Prints information on the current state of the object.
    	--          Is used to redefine the operator <<.

    is static;


fields

Done:         Boolean;
AA:           Matrix;
NbRotations:  Integer;
EigenValues:  Vector;
EigenVectors: Matrix;

end Jacobi;
