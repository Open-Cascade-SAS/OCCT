-- File:	ShapeFix_Shell.cdl
-- Created:	Wed Aug 12 10:26:46 1998
-- Author:	Galina KULIKOVA
--		<gka@nnov.matra-dtv.fr>
---Copyright:	 Matra Datavision 1998


class Shell from ShapeFix inherits Root from ShapeFix

	---Purpose: Fixing orientation of faces in shell

uses

    Compound            from TopoDS,
    Shell               from TopoDS,
    Shape               from TopoDS,
    Status              from ShapeExtend,
    BasicMsgRegistrator from ShapeExtend,
    Face                from ShapeFix,
    ProgressIndicator   from Message
    
is

    Create returns Shell from ShapeFix;
    	---Purpose: Empty constructor

    Create (shape: Shell from TopoDS)
    returns Shell from ShapeFix;
    	---Purpose: Initializes by shell.

    Init (me: mutable; shell: Shell from TopoDS);
    	---Purpose: Initializes by shell.

    Perform (me: mutable;
             theProgress : ProgressIndicator from Message = 0) returns Boolean;
        ---Purpose: Iterates on subshapes and performs fixes
        --          (for each face calls ShapeFix_Face::Perform and
        --          then calls FixFaceOrientation). The passed progress
        --          indicator allows user to consult the current progress
        --          stage and abort algorithm if needed.

    FixFaceOrientation (me : mutable; shell : Shell from TopoDS;
    	    	    	isAccountMultiConex : Boolean = Standard_True;
    	    	    	NonManifold : Boolean = Standard_False ) returns Boolean;
      ---Purpose: Fixes orientation of faces in shell.
      --          Changes orientation of face in the shell, if it is oriented opposite
      --          to neigbouring faces. If it is not possible to orient all faces in the
      --          shell (like in case of mebious band), this method orients only subset
      --          of faces. Other faces are stored in Error compound.
      --          Modes : 
      --    	    isAccountMultiConex - mode for account cases of multiconnexity.
      --          If this mode is equal to Standard_True, separate shells will be created 
      --          in the cases of multiconnexity. If this mode is equal to Standard_False,
      --          one shell will be created without account of multiconnexity.By defautt - Standard_True;
      --          NonManifold - mode for creation of non-manifold shells.
      --          If this mode is equal to Standard_True one non-manifold will be created from shell
      --          contains multishared edges. Else if this mode is equal to Standard_False only 
      --          manifold shells will be created. By default - Standard_False.
      --          
      ---Returns: If resulting shell is ok returns TRUE, else returns FALSE.
      ---Status : OK   - faces in shall were oriented correcty.
      --          DONE - faces in shell oriented succesfully
      --          FAIL - faces orientation process has been failed
	
    Shell(me : mutable) returns Shell from TopoDS;
    	---Purpose: Returns fixed shell (or subset of oriented faces).
	
    Shape(me : mutable) returns Shape from TopoDS;
    	---Purpose: In case of multiconnexity returns compound of fixed shells
    	--          else returns one shell..
    NbShells(me) returns Integer;
    	---Purpose: Returns Number of obtainrd shells;
	
    ErrorFaces(me) returns Compound from TopoDS;
    	---Purpose: Returns not oriented subset of faces.

    Status (me; status : Status from  ShapeExtend) returns Boolean;
    	---Purpose: Returns the status of the last Fix.

    FixFaceTool (me:mutable) returns Face from ShapeFix;
    	---Purpose: Returns tool for fixing faces.
      ---C++:inline

    SetMsgRegistrator (me: mutable; msgreg: BasicMsgRegistrator from ShapeExtend) is redefined;
      ---Purpose: Sets message registrator

    SetPrecision (me: mutable; preci: Real) is redefined;
    	---Purpose: Sets basic precision value (also to FixWireTool)

    SetMinTolerance (me: mutable; mintol: Real) is redefined;
    	---Purpose: Sets minimal allowed tolerance (also to FixWireTool)

    SetMaxTolerance (me: mutable; maxtol: Real) is redefined;
    	---Purpose: Sets maximal allowed tolerance (also to FixWireTool)

    FixFaceMode (me: mutable) returns Integer;
    	---C++: return &
      ---C++: inline
      ---Purpose: Returns (modifiable) the mode for applying fixes of 
      --          ShapeFix_Face, by default True.

    FixOrientationMode (me: mutable) returns Integer;
    	---C++: return &
      ---C++: inline
      ---Purpose: Returns (modifiable) the mode for applying 
      --          FixFaceOrientation, by default True.
    
fields

    myShell              : Shell from TopoDS is protected;
    myErrFaces           : Compound from TopoDS is protected;
    myStatus             : Integer is protected;
    myFixFace            : Face from ShapeFix is protected;
    myFixFaceMode        : Integer is protected;   
    myFixOrientationMode : Integer is protected; 
    myNbShells           : Integer is protected; 

end Shell;
