-- Created on: 1993-01-09
-- Created by: CKY / Contract Toubro-Larsen ( TCD )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class LineFontPredefined from IGESGraph  inherits IGESEntity

        ---Purpose: defines IGESLineFontPredefined, Type <406> Form <19>
        --          in package IGESGraph
        --
        --          Provides the ability to specify a line font pattern
        --          from a predefined list rather than from
        --          Directory Entry Field 4

uses  Integer  -- no one specific type


is

        Create returns mutable LineFontPredefined;

        -- Specific Methods pertaining to the class

        Init (me                   : mutable;
              nbProps              : Integer;
              aLineFontPatternCode : Integer);
        ---Purpose : This method is used to set the fields of the class
        --           LineFontPredefined
        --       - nbProps              : Number of property values (NP = 1)
        --       - aLineFontPatternCode : Line Font Pattern Code

        -- Specific Access Methods : According to each type of Entity

        NbPropertyValues (me) returns Integer;
        ---Purpose : returns the number of property values in <me>

        LineFontPatternCode (me) returns Integer;
        ---Purpose : returns the Line Font Pattern Code of <me>

fields

--
-- Class    : IGESGraph_LineFontPredefined
--
-- Purpose  : Declaration of the variables specific to a
--            LineFontPredefined property.
--
-- Reminder : A LineFontPredefined property is defined by :
--                  - Number of property values
--                  - Line Font Pattern Code
--

        theNbPropertyValues    : Integer;

        theLineFontPatternCode : Integer;

end LineFontPredefined;
