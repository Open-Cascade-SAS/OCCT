-- File:	StepToGeom_MakeParabola.cdl
-- Created:	Thu Sep  8 09:00:04 1994
-- Author:	Frederic MAUPAS
---Copyright:	 Matra Datavision 1994

class MakeParabola from StepToGeom

    ---Purpose: This class implements the mapping between classes 
    --          Parabola from StepGeom which describes a Parabola from
    --          Prostep and Parabola from Geom.

uses 
     Parabola from Geom,
     Parabola from StepGeom

is 

    Convert ( myclass; SC : Parabola from StepGeom;
                       CC : out Parabola from Geom )
    returns Boolean from Standard;

end MakeParabola;
