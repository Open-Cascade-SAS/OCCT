-- Created on: 1990-12-11
-- Created by: Remi Lequette
-- Copyright (c) 1990-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package TopoDS 

    ---Purpose: Provides methods to cast objects of class
-- TopoDS_Shape to be onjects of more specialized
-- sub-classes. Types are verified, thus in the example
-- below, the first two blocks are correct but the third is
-- rejected by the compiler.

uses
    MMgt,
    TCollection,
    TopAbs,      -- basic enumerations : ShapeEnum, Orientation
    TopLoc       -- the Location (Local Coordinate System)

is

    -- exceptions

    exception FrozenShape inherits DomainError;
	---Purpose: An  attempt was  made to   modify  a Shape  already
	--          shared or protected.

    exception LockedShape inherits DomainError;
	---Purpose: An attempt was made to modify a geometry of Shape already
	--          shared or protected.
	
    exception UnCompatibleShapes inherits DomainError;
	---Purpose: An incorrect insertion was attempted.
	
    -- classes

    class Shape;

    class HShape;

    class ListOfShape instantiates List from TCollection (Shape from TopoDS);
	---Purpose: Used to implement the TShape.

    deferred class TShape;

    deferred class TVertex;

    class Vertex;

    deferred class TEdge;

    class Edge;

    class TWire;

    class Wire;

    class TFace;

    class Face;

    class TShell;

    class Shell;

    class TSolid;

    class Solid;

    class TCompSolid;

    class CompSolid;

    class TCompound;

    class Compound;

    class Builder;

    class Iterator;
	---Purpose: Basic tool to access the data structure.

    Vertex(S : Shape from TopoDS) returns Vertex from TopoDS
	---C++: inline
	---C++: return const &
	---C++: alias "inline static TopoDS_Vertex& Vertex(TopoDS_Shape&);"
    ---Purpose: Casts shape S to the more specialized return type, Vertex.
    -- Exceptions
    -- Standard_TypeMismatch if S cannot be cast to this return type.
    raises TypeMismatch from Standard;

    Edge(S : Shape from TopoDS) returns Edge from TopoDS
	---C++: inline
	---C++: return const &
	---C++: alias "inline static TopoDS_Edge& Edge(TopoDS_Shape&);"
    ---Purpose: Casts shape S to the more specialized return type, Edge
    -- Exceptions
    -- Standard_TypeMismatch if S cannot be cast to this return type.
    raises TypeMismatch from Standard;

    Wire(S : Shape from TopoDS) returns Wire from TopoDS
	---C++: inline
	---C++: return const &
	---C++: alias "inline static TopoDS_Wire& Wire(TopoDS_Shape&);"
    ---Purpose: Casts shape S to the more specialized return type, Wire.
    -- Exceptions
    -- Standard_TypeMismatch if S cannot be cast to this return type.
    raises TypeMismatch from Standard;

    Face(S : Shape from TopoDS) returns Face from TopoDS
	---C++: inline
	---C++: return const &
	---C++: alias "inline static TopoDS_Face& Face(TopoDS_Shape&);"
    ---Purpose: Casts shape S to the more specialized return type, Face.
    -- Exceptions
    -- Standard_TypeMismatch if S cannot be cast to this return type.
    raises TypeMismatch from Standard;

    Shell(S : Shape from TopoDS) returns Shell from TopoDS
	---C++: inline
	---C++: return const &
	---C++: alias "inline static TopoDS_Shell& Shell(TopoDS_Shape&);"
    ---Purpose: Casts shape S to the more specialized return type, Shell.
    -- Exceptions
    -- Standard_TypeMismatch if S cannot be cast to this return type.
    raises TypeMismatch from Standard;

    Solid(S : Shape from TopoDS) returns Solid from TopoDS
	---C++: inline
	---C++: return const &
	---C++: alias "inline static TopoDS_Solid& Solid(TopoDS_Shape&);"
    ---Purpose: Casts shape S to the more specialized return type, Solid.
    -- Exceptions
    -- Standard_TypeMismatch if S cannot be cast to this return type.
    raises TypeMismatch from Standard;

    CompSolid(S : Shape from TopoDS) returns CompSolid from TopoDS
	---C++: inline
	---C++: return const &
	---C++: alias "inline static TopoDS_CompSolid& CompSolid(TopoDS_Shape&);"
    ---Purpose: Casts shape S to the more specialized return type, CompSolid.
    -- Exceptions
    -- Standard_TypeMismatch if S cannot be cast to this return type.
    raises TypeMismatch from Standard;

    Compound(S : Shape from TopoDS) returns Compound from TopoDS
	---C++: inline
	---C++: return const &
	---C++: alias "inline static TopoDS_Compound& Compound(TopoDS_Shape&);"
    ---Purpose: Casts shape S to the more specialized return type, Compound.
    -- Exceptions
    -- Standard_TypeMismatch if S cannot be cast to this return type.
    raises TypeMismatch from Standard;

end TopoDS;
