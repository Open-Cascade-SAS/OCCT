-- Created on: 1995-02-07
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class LineConstructor from IntTools

        ---Purpose: Splits given Line.

uses Line           from IntPatch,
     TopolTool      from Adaptor3d,
     HSurface       from GeomAdaptor,
     SequenceOfReal from TColStd


raises NotDone    from StdFail,
       OutOfRange from Standard

is

    Create
    	returns LineConstructor from IntTools;
	---C++: inline
	---Purpose: 
	--- Empty constructor
	---

    Load(me: in out; D1,D2: TopolTool from Adaptor3d;
                     S1,S2: HSurface  from GeomAdaptor)
    	is static;
	---C++: inline
	---Purpose:
	--- Initializes me by two surfaces and corresponding
	--- tools which represent boundaries of surfaces
	---

    Perform(me: in out; L: Line from IntPatch)
    	is static;
	---Purpose:
	--- Splits line
	---

    IsDone(me)
    	returns Boolean from Standard
	is static;
	---C++: inline
	---Purpose:
	--- Returns True if splitting was successful
	---

    NbParts(me)
    	returns Integer from Standard
	raises NotDone from StdFail
	is static;
	---C++: inline
	---Purpose:
	--- Returns number of splits
	---

    Part(me; I: Integer from Standard; WFirst,WLast: out Real from Standard) 
    	raises NotDone    from StdFail,
               OutOfRange from Standard
	is static;
	---C++: inline
	---Purpose:
	--- Return first and last parameters 
    	--- for given index of split
	---

    ---PeriodicLine(me; L: Line from IntPatch)
    ---	is protected;
 
    TreatCircle(me:out; 
    	    aLine : Line from IntPatch; 
    	    aTol: Real from Standard)
    	is protected; 
	
fields
    
    done  : Boolean        from Standard;
    seqp  : SequenceOfReal from TColStd;
    myDom1: TopolTool      from Adaptor3d;
    myDom2: TopolTool      from Adaptor3d;
    myHS1 : HSurface       from GeomAdaptor;
    myHS2 : HSurface       from GeomAdaptor;    

end LineConstructor;
