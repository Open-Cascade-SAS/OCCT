-- Created on: 2008-08-15
-- Created by: Sergey ZARITCHNY <szy@opencascade.com>
-- Copyright (c) 2008-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Naming_1 from PNaming inherits Attribute from PDF

	---Purpose: 
uses 
    Name_1 from PNaming
			    
is
    Create
    returns mutable Naming_1 from PNaming;
    
    SetName(me : mutable ; aName : Name_1 from PNaming);

    GetName(me) returns Name_1 from PNaming;

fields

    myName :  Name_1 from PNaming;


end Naming_1;
