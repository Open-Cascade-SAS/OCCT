-- File:        StepAP214_AppliedDateAndTimeAssignment.cdl
-- Created:     Tue Mar 9 11:11:13 1999
-- Author:      data exchange team
--		<det@androx.nnov.matra-dtv.fr>
-- Copyright:   Matra-Datavision 1999


class AppliedDateAndTimeAssignment from StepAP214 

inherits DateAndTimeAssignment from StepBasic 

uses

	HArray1OfDateAndTimeItem from StepAP214, 
	DateAndTimeItem from StepAP214, 
	DateAndTime from StepBasic, 
	DateTimeRole from StepBasic
is

	Create returns mutable AppliedDateAndTimeAssignment;
	---Purpose: Returns a AppliedDateAndTimeAssignment


	Init (me : mutable;
	      aAssignedDateAndTime : mutable DateAndTime from StepBasic;
	      aRole : mutable DateTimeRole from StepBasic) is redefined;

	Init (me : mutable;
	      aAssignedDateAndTime : mutable DateAndTime from StepBasic;
	      aRole : mutable DateTimeRole from StepBasic;
	      aItems : mutable HArray1OfDateAndTimeItem from StepAP214) is virtual;

	-- Specific Methods for Field Data Access --

	SetItems(me : mutable; aItems : mutable HArray1OfDateAndTimeItem);
	Items (me) returns mutable HArray1OfDateAndTimeItem;
	ItemsValue (me; num : Integer) returns DateAndTimeItem;
	NbItems (me) returns Integer;

fields

	items : HArray1OfDateAndTimeItem from StepAP214; -- a SelectType

end AppliedDateAndTimeAssignment;
