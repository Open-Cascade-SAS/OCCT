-- Created on: 1995-05-17
-- Created by: Mister rmi
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

private class ListOfTransient from V3d inherits ListOfTransient from TColStd

is

    Create returns ListOfTransient from V3d;
    
    Contains(me; aTransient: Transient from Standard)
    returns Boolean from Standard
    is static;
    
    Remove(me: in out; aTransient: Transient from Standard)
    is static;
    
    
end ListOfTransient from V3d;
