-- Created on: 2007-01-25
-- Created by: Sergey KOCHETKOV
-- Copyright (c) 2007-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class SensitiveMesh from MeshVS inherits SensitiveEntity from Select3D

	---Purpose: This class provides custom mesh sensitive entity used in advanced mesh selection.  
    	---It provides detection of mesh entities accordingly to activated selection mode 

uses
  EntityOwner from SelectBasics,
  Array1OfPnt2d from TColgp, 
  Box from Bnd, 
  Box2d from Bnd, 
  Location from TopLoc, 
  Lin from gp, 
  ListOfBox2d from SelectBasics,
  PickArgs from SelectBasics,
  Projector from Select3D      
is

  Create ( theOwner    : EntityOwner from SelectBasics; 
           theMode     : Integer = 0 )
    returns mutable SensitiveMesh from MeshVS; 
      
  GetMode( me ) returns Integer from Standard;     
     
  GetConnected( me: mutable;  aLocation  :  Location from TopLoc )
    returns SensitiveEntity from Select3D is redefined; 

  Matches (me : mutable;
           thePickArgs : PickArgs from SelectBasics;
           theMatchDMin, theMatchDepth : out Real from Standard)
    returns Boolean is redefined;

  Matches  ( me: mutable;   XMin, YMin, XMax, YMax  : Real;
             	    	    aTol                    : Real ) returns Boolean  
    is redefined;

  Matches  ( me: mutable;   Polyline  :  Array1OfPnt2d from TColgp;
                            aBox      :  Box2d;  
    	    	    	    aTol      :  Real ) returns Boolean  
    is redefined; 
      
  Project ( me:mutable; aProjector : Projector from Select3D ) is redefined static;
     
  Areas   ( me: mutable ; boxes : in out ListOfBox2d from SelectBasics ) is redefined static;  
   
  ProjectOneCorner( me: mutable; aProjector : Projector from Select3D; 
    	    	    	    	 X,Y,Z      : Real from Standard ) is private;     
 
fields 
   
  myMode  : Integer from Standard;          
  mybox   : Box    from Bnd; 
  mybox2d : Box2d  from Bnd;   
 
end SensitiveMesh;
