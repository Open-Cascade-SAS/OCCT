-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SurfaceStyleFillArea from StepVisual 

inherits TShared from MMgt

uses

	FillAreaStyle from StepVisual
is

	Create returns mutable SurfaceStyleFillArea;
	---Purpose: Returns a SurfaceStyleFillArea

	Init (me : mutable;
	      aFillArea : mutable FillAreaStyle from StepVisual) is virtual;

	-- Specific Methods for Field Data Access --

	SetFillArea(me : mutable; aFillArea : mutable FillAreaStyle);
	FillArea (me) returns mutable FillAreaStyle;

fields

	fillArea : FillAreaStyle from StepVisual;

end SurfaceStyleFillArea;
