-- Created on: 1995-10-17
-- Created by: Andre LIEUTIER
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


package Plate

uses
     TCollection,  TColStd,
     math, gp, TColgp
is

    class Plate; 
    
-- Basic  Constraints Class
    class PinpointConstraint;
    class LinearScalarConstraint;
    class LinearXYZConstraint;
--
-- geometric Constraints Class
--
    class GlobalTranslationConstraint;  
--    
    class PlaneConstraint; 
    class LineConstraint;  
--  
    class SampledCurveConstraint;
--   
--  class LinearizedHighlightConstraint;
--  
--  class DirectionalPressureConstraint;
--  
--  
--  Geometric contact of order k Constraint 
    class GtoCConstraint;
    class FreeGtoCConstraint;


-- utilities and internal Classes
    class D1;
    class D2;
    class D3;
    class SequenceOfPinpointConstraint instantiates Sequence from TCollection  
                                       (PinpointConstraint from Plate);
    class SequenceOfLinearXYZConstraint instantiates Sequence from TCollection  
                                       (LinearXYZConstraint from Plate);
    class SequenceOfLinearScalarConstraint instantiates Sequence from TCollection  
                                       (LinearScalarConstraint from Plate);
    class Array1OfPinpointConstraint instantiates Array1 from TCollection
                                       (PinpointConstraint from Plate);    
    class HArray1OfPinpointConstraint instantiates HArray1 from TCollection
                                       (PinpointConstraint         from Plate,
                                        Array1OfPinpointConstraint from Plate);    
end Plate;
