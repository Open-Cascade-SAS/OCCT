-- Created on: 2003-06-04
-- Created by: Galina KULIKOVA
-- Copyright (c) 2003-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class GeometricTolerance from StepDimTol
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity GeometricTolerance

uses
    HAsciiString from TCollection,
    MeasureWithUnit from StepBasic,
    ShapeAspect from StepRepr

is
    Create returns GeometricTolerance from StepDimTol;
	---Purpose: Empty constructor

    Init (me: mutable; aName: HAsciiString from TCollection;
                       aDescription: HAsciiString from TCollection;
                       aMagnitude: MeasureWithUnit from StepBasic;
                       aTolerancedShapeAspect: ShapeAspect from StepRepr);
	---Purpose: Initialize all fields (own and inherited)

    Name (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Name
    SetName (me: mutable; Name: HAsciiString from TCollection);
	---Purpose: Set field Name

    Description (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Description
    SetDescription (me: mutable; Description: HAsciiString from TCollection);
	---Purpose: Set field Description

    Magnitude (me) returns MeasureWithUnit from StepBasic;
	---Purpose: Returns field Magnitude
    SetMagnitude (me: mutable; Magnitude: MeasureWithUnit from StepBasic);
	---Purpose: Set field Magnitude

    TolerancedShapeAspect (me) returns ShapeAspect from StepRepr;
	---Purpose: Returns field TolerancedShapeAspect
    SetTolerancedShapeAspect (me: mutable; TolerancedShapeAspect: ShapeAspect from StepRepr);
	---Purpose: Set field TolerancedShapeAspect

fields
    theName: HAsciiString from TCollection;
    theDescription: HAsciiString from TCollection;
    theMagnitude: MeasureWithUnit from StepBasic;
    theTolerancedShapeAspect: ShapeAspect from StepRepr;

end GeometricTolerance;
