-- File:	StepData_SelectNamed.cdl
-- Created:	Mon Dec 16 16:44:07 1996
-- Author:	Christian CAILLET
--		<cky@heliox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1996


class SelectNamed  from StepData    inherits SelectMember

    ---Purpose : This select member can be of any kind, and be named
    --           But its takes more memory than some specialised ones
    --           This class allows one name for the instance

uses CString, Logical, AsciiString from TCollection,  Field from StepData

is

    Create  returns mutable SelectNamed;

    HasName (me) returns Boolean  is redefined;

    Name (me) returns CString  is redefined;

    SetName (me : mutable; name : CString)  returns Boolean  is redefined;
    -- redefined to accept any name

    Field (me) returns Field;
    ---C++ : return const &

    CField (me : mutable) returns Field;
    ---C++ : return &


    Kind (me) returns Integer  is redefined;
    --  see Field for Kind (same codes)

    SetKind  (me : mutable; kind : Integer)  is redefined;
    --  called by various Set*

    Int (me) returns Integer  is redefined;
    ---Purpose : This internal method gives access to a value implemented by an
    --           Integer (to read it)

    SetInt (me : mutable; val : Integer)  is redefined;
    ---Purpose : This internal method gives access to a value implemented by an
    --           Integer (to set it)

    Real (me) returns Real  is redefined;

    SetReal (me : mutable; val : Real)  is redefined;

    String (me) returns CString  is redefined;

    SetString (me : mutable; val : CString)  is redefined;

fields

    thename : AsciiString;
    theval  : Field from StepData;

end SelectNamed;
