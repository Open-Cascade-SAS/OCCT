-- File:	SelectMgr_Filter.cdl
-- Created:	Wed Mar  5 13:51:25 1997
-- Author:	Robert COUBLANC
--		<rob@robox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1997


deferred class Filter from SelectMgr inherits TShared from MMgt

	---Purpose: The root class to define filter objects for selection.
    	-- Advance handling of objects requires the services of
    	-- filters. These only allow dynamic detection and
    	-- selection of objects which correspond to the criteria defined in each.
    	-- Eight standard filters inheriting SelectMgr_Filter are
    	-- defined in Open CASCADE.
    	--  You can create your own filters by defining new filter
    	-- classes inheriting this framework. You use these
    	-- filters by loading them into an AIS interactive context. 

uses
     EntityOwner from SelectMgr,
     ShapeEnum from TopAbs
is
    IsOk(me; anObj : EntityOwner from SelectMgr)
    returns Boolean from Standard
    is deferred;
    	---Purpose: Indicates that the selected Interactive Object
    	-- passes the filter. The owner, anObj, can be either
    	-- direct or user. A direct owner is the corresponding
    	-- construction element, whereas a user is the
    	-- compound shape of which the entity forms a part.
    	-- When an object is detected by the mouse - in AIS,
    	-- this is done through a context selector - its owner
    	-- is passed to the filter as an argument.
    	-- If the object returns Standard_True, it is kept; if
    	-- not, it is rejected.
    	-- If you are creating a filter class inheriting this
    	-- framework, and the daughter class is to be used in
    	-- an AIS local context, you will need to implement the
    	-- virtual function ActsOn.
        
    ActsOn(me; aStandardMode : ShapeEnum from TopAbs)
    returns Boolean from Standard is virtual;
	---Purpose: Returns true in an AIS local context, if this filter
    	-- operates on a type of subshape defined in a filter
    	-- class inheriting this framework.
    	-- This function completes IsOk in an AIS local context.
    

end Filter;
