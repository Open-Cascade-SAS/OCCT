-- Created on: 1994-01-25
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

generic class Extremity from Blend 
    (TheVertex               as any;
     TheArc                  as any;
     ThePointOnRst           as any; -- as PointOnRst from Blend(TheArc)
     TheSequenceOfPointOnRst as any) -- as Iterator   from Blend(ThePointOnRst)



	---Purpose: 

uses Pnt from gp, 
     Vec from  gp,
     Transition from IntSurf


raises DomainError from Standard,
       OutOfRange  from Standard

is

    Create
    
    	returns Extremity from Blend;


    Create(P: Pnt from gp; 
           U,V,Param: Real from Standard; Tol: Real from Standard)
	---Purpose: Creates an extremity on a surface
    	returns Extremity from Blend;


    Create(P: Pnt from gp; 
           U,V,Param: Real from Standard; Tol: Real from Standard;
           Vtx: TheVertex)
	---Purpose: Creates an extremity on a surface. This extremity matches
	--          the vertex <Vtx>.

    	returns Extremity from Blend;


    Create(P: Pnt from gp; 
           W,  Param: Real from Standard; Tol: Real from Standard)
	---Purpose: Creates an extremity on a curve
    	returns Extremity from Blend;


    SetValue(me: in out; P: Pnt from gp; 
    	    	    	 U,V,Param : Real from Standard;
                         Tol: Real from Standard)
	---Purpose: Set the values for an extremity on a surface.
    	is static;


    SetValue(me: in out; P: Pnt from gp; 
                         U,V,Param: Real from Standard;
                         Tol: Real from Standard; Vtx: TheVertex)
	---Purpose: Set the values for an extremity on a surface.This
	--          extremity matches the vertex <Vtx>.
    	is static;


    SetValue(me: in out; P: Pnt from gp;
                         W,Param: Real from Standard;
                         Tol: Real from Standard)
	---Purpose: Set the values for an extremity on curve.
    	is static;


    Value(me)
    
	---Purpose: This method returns the value of the point in 3d space.
    
    	returns Pnt from gp
	---C++: inline
	---C++: return const&
	
	is static; 
	 
    SetTangent(me: in out; Tangent  : Vec from gp) 
	---Purpose:   Set the tangent   vector  for an extremity on  a
	--          surface.
	---C++: inline
    	is static;	
 
     HasTangent(me)

	---Purpose: Returns TRUE if the Tangent is  stored.

    	returns Boolean from Standard
	---C++: inline
	
	is static;      
   
    Tangent(me) 
    
    	---Purpose: This  method returns the   value of tangent  in 3d
    	--          space.
    
    	returns Vec from gp
	---C++: inline
	---C++: return const&
	
    	is static; 

    Tolerance(me)
    
	---Purpose: This method returns the fuzziness on the point
	--          in 3d space.
    
    	returns Real from Standard
	---C++: inline
	
	is static;



-- methods for an extremity on a surface

    SetVertex(me: in out; V: TheVertex)
	---Purpose: Set the values for an extremity on a curve.
    	is static;


    AddArc(me: in out; A: TheArc; Param: Real from Standard;
                       TLine, TArc: Transition from IntSurf)

	---Purpose: Sets the values of a point which is on the arc
	--          A, at parameter Param.


    	is static;


    Parameters(me; U,V: out Real from Standard)
    
	---Purpose: This method returns the parameters of the point
	--          on the concerned surface.
    
	---C++: inline
	is static;


    IsVertex(me)
    
	---Purpose: Returns Standard_True when the point coincide with
	--          an existing vertex.
    
    	returns Boolean from Standard
	---C++: inline

	is static;


    Vertex(me)
    
	---Purpose: Returns the vertex when IsVertex returns Standard_True.
    
    	returns any TheVertex
	---C++: inline
	---C++: return const&

    	raises DomainError from Standard
	--- The exception is raised when IsVertex returns Standard_False
    	is static;


    NbPointOnRst(me)
    
	---Purpose: Returns the number of arc containing the extremity.
	--          If the method returns 0, the point is inside the
	--          surface.
	--          Otherwise, the extremity lies on at least 1 arc,
	--          and all the information (arc, parameter, transitions)
	--          are given by the point on restriction (PointOnRst)
	--          returned by the next method.
    
    	returns Integer from Standard
	---C++: inline
	
	is static;


    PointOnRst(me; Index: Integer from Standard)
    
	---Purpose: 
    
    	returns any ThePointOnRst
	---C++: inline
	---C++: return const&

	raises OutOfRange from Standard
	--- The exception is raised when Index <=0 or Index > NbPointOnRst
	is static;


-- method for an extremity on a curve

    Parameter(me)
    
    	returns Real from Standard
	---C++: inline
	is static; 
	 
-- method for the parameter on the guide
   ParameterOnGuide(me) 
    
    	returns Real from Standard
	---C++: inline
	is static;  

fields
    vtx    : TheVertex;
    seqpt  : TheSequenceOfPointOnRst;
    pt     : Pnt     from gp;   
    tang   : Vec     from gp;
    param  : Real    from Standard;
    u      : Real    from Standard;
    v      : Real    from Standard;
    tol    : Real    from Standard;
    isvtx  : Boolean from Standard;
    hastang: Boolean from Standard;

end Extremity;


