-- File:	StepToGeom_MakeDirection2d.cdl
-- Created:	Wed Aug  4 11:49:16 1993
-- Author:	Martine LANGLOIS
---Copyright:	 Matra Datavision 1993

class MakeDirection2d from StepToGeom

    ---Purpose: This class implements the mapping between classes 
    --          Direction from StepGeom which describes a direction
    --          from Prostep and Direction from Geom2d.

uses 
     Direction from Geom2d,
     Direction from StepGeom

is 

    Convert ( myclass; SD : Direction from StepGeom;
                       CD : out Direction from Geom2d )
    returns Boolean from Standard;

end MakeDirection2d;
