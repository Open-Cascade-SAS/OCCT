-- Created on: 1998-05-06
-- Created by: Andre LIEUTIER
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class SampledCurveConstraint from Plate
---Purpose: define m PinPointConstraint driven by m unknown
--          
--          
--          
--                   
uses 
 SequenceOfPinpointConstraint from Plate, 
 LinearXYZConstraint from Plate
raises
    DimensionMismatch from Standard

is
    Create(SOPPC  :  SequenceOfPinpointConstraint; 
    	    n  :  Integer) 
    	    returns SampledCurveConstraint
	    raises DimensionMismatch from Standard;
    --  n have to be less than the length of SOPPC
    --  

     -- Accessors :
    LXYZC(me) returns LinearXYZConstraint;
    ---C++: inline 
    ---C++: return const &

fields
    myLXYZC : LinearXYZConstraint;
    
end;


