-- Created on: 1992-02-14
-- Created by: Jean Claude VAUTHIER
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.







class PGProps

from GProp

inherits GProps
---Purpose: A framework for computing the global properties of a
-- set of points.
-- A point mass is attached to each point. The global
-- mass of the system is the sum of each individual
-- mass. By default, the point mass is equal to 1 and the
-- mass of a system composed of N points is equal to N.
-- Warning
-- A framework of this sort provides functions to handle
-- sets of points easily. But, like any GProp_GProps
-- object, by using the Add function, it can theoretically
-- bring together the computed global properties and
-- those of a system more complex than a set of points .
-- The mass of each point and the density of each
-- component of the composed system must be
-- coherent. Note that this coherence cannot be checked.
-- Nonetheless, you are advised to restrict your use of a
-- GProp_PGProps object to a set of points and to
-- create a GProp_GProps object in order to bring
-- together global properties of different systems.
        
uses Pnt          from gp,
     Array1OfPnt  from TColgp,
     Array2OfPnt  from TColgp,
     Array1OfReal from TColStd,
     Array2OfReal from TColStd

     
raises DimensionError from Standard,
       DomainError    from Standard
     
is

  Create   returns PGProps;
        --- Purpose : Initializes a framework to compute global properties
-- on a set of points.
-- The point relative to which the inertia of the system is
-- computed will be the origin (0, 0, 0) of the
-- absolute Cartesian coordinate system.
-- At initialization, the framework is empty, i.e. it retains
-- no dimensional information such as mass and inertia.
-- It is, however, now able to keep global properties of a
-- set of points while new points are added using the
-- AddPoint function.
-- The set of points whose global properties are brought
-- together by this framework will then be referred to as
-- the current system. The current system is, however,
-- not kept by this framework, which only keeps that
-- system's global properties. Note that the current
-- system may be more complex than a set of points.
       

  AddPoint (me : in out; P : Pnt)
        --- Purpose : Brings together the global properties already
-- retained by this framework with those induced by
-- the point Pnt. Pnt may be the first point of the current system.
-- A point mass is attached to the point Pnt, it is either
-- equal to 1. or to Density.
            is static;


  AddPoint (me : in out; P : Pnt; Density : Real)
        --- Purpose :
        --  Adds a new point P with its density in the system of points
   -- Exceptions
-- Standard_DomainError if the mass value Density
-- is less than gp::Resolution().
      raises DomainError
     is static;
     
     
  Create (Pnts : Array1OfPnt) returns PGProps;
        --- Purpose :
        --  computes the global properties of the system of points Pnts.
        --  The density of the points are defaulted to all being 1


  Create (Pnts : Array2OfPnt) returns PGProps;
        --- Purpose :
        --  computes the global properties of the system of points Pnts.
        --  The density of the points are defaulted to all being 1


  Create (Pnts : Array1OfPnt; Density : Array1OfReal) returns PGProps
        --- Purpose :
        --  computes the global properties of the system of points Pnts.
        --  A density is associated with each point.
     raises DomainError,
        --- Purpose : 
        --  raises if a density is lower or equal to Resolution from package
        --  gp.
            DimensionError;
        --- Purpose : 
        --  raises if the length of Pnts and the length of Density
        --  is not the same.



  Create (Pnts : Array2OfPnt; Density : Array2OfReal) returns PGProps
        --- Purpose :
        --  computes the global properties of the system of points Pnts.
        --  A density is associated with each point.
     raises DomainError,
        --- Purpose : 
        --  Raised if a density is lower or equal to Resolution from package
        --  gp.
            DimensionError;
        --- Purpose : 
        --  Raised if the length of Pnts and the length of Density
        --  is not the same.




  Barycentre (myclass; Pnts : Array1OfPnt from TColgp)  returns Pnt;
        --- Purpose : 
        --  Computes the barycentre of a set of points. The density of the
        --  points is defaulted to 1.


  Barycentre (myclass; Pnts : Array2OfPnt from TColgp)   returns Pnt;
        --- Purpose : 
        --  Computes the barycentre of a set of points. The density of the
        --  points is defaulted to 1.


  Barycentre (myclass; Pnts : Array1OfPnt from TColgp; 
              Density : Array1OfReal from TColStd;
              Mass : out Real; G : out Pnt)
        --- Purpose : 
        --  Computes the barycentre of a set of points. A density is associated
        --  with each point.
     raises DomainError,
        --- Purpose : 
        --  raises if a density is lower or equal to Resolution from package
        --  gp.
            DimensionError;
        --- Purpose : 
        --  Raised if the length of Pnts and the length of Density
        --  is not the same.


  Barycentre (myclass; Pnts : Array2OfPnt from TColgp; 
              Density : Array2OfReal from TColStd;
              Mass : out Real; G : out Pnt)
        --- Purpose : 
        --  Computes the barycentre of a set of points. A density is associated
        --  with each point.
     raises DomainError,
        --- Purpose : 
        --  Raised if a density is lower or equal to Resolution from package
        --  gp.
            DimensionError;
        --- Purpose : 
        --  Raised if the length of Pnts and the length of Density
        --  is not the same.


end PGProps;



