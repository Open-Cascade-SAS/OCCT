-- File:	StepToGeom_MakeEllipse.cdl
-- Created:	Thu Sep  1 13:46:53 1994
-- Author:	Frederic MAUPAS
---Copyright:	 Matra Datavision 1994

class MakeEllipse from StepToGeom

    ---Purpose: This class implements the mapping between classes 
    --          Ellipse from StepGeom which describes a Ellipse from
    --          Prostep and Ellipse from Geom.
  
uses 
     Ellipse from Geom,
     Ellipse from StepGeom

is 

    Convert ( myclass; SC : Ellipse from StepGeom;
                       CC : out Ellipse from Geom )
    returns Boolean from Standard;

end MakeEllipse;
