-- Created on: 2001-09-11
-- Created by: Julia DOROVSKIKH
-- Copyright (c) 2001-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



package XmlXCAFDrivers 

        ---Purpose: 

uses
    TCollection,
    CDM,
    XmlDrivers,
    XmlMDF
    
is
    class DocumentRetrievalDriver;
    
    class DocumentStorageDriver;

    ---Category: Factory methods
    --           ==============================================================

    Factory (aGUID: GUID from Standard)
    returns Transient from Standard;
        ---Purpose: Depending from the  ID, returns a list of  storage
        --          or retrieval attribute drivers. Used for plugin.
        --          
        --          Standard data model drivers
        --          ===========================
        --          47b0b826-d931-11d1-b5da-00a0c9064368 Transient-Persistent 
        --          47b0b827-d931-11d1-b5da-00a0c9064368 Persistent-Transient
        --          
        --          XCAF data model drivers
        --          =================================
        --          ed8793f8-3142-11d4-b9b5-0060b0ee281b Transient-Persistent 
        --          ed8793f9-3142-11d4-b9b5-0060b0ee281b Persistent-Transient
        --          ed8793fa-3142-11d4-b9b5-0060b0ee281b XCAFSchema


end XmlXCAFDrivers;
