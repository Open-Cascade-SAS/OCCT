-- File:        DateTimeSelect.cdl
-- Created:     Fri Dec  1 11:11:11 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993



class DateTimeSelect from StepBasic inherits SelectType from StepData

	-- <DateTimeSelect> is an EXPRESS Select Type construct translation.
	-- it gathers : Date, LocalTime, DateAndTime

uses

	Date,
	LocalTime,
	DateAndTime
is

	Create returns DateTimeSelect;
	---Purpose : Returns a DateTimeSelect SelectType

	CaseNum (me; ent : Transient) returns Integer;
	---Purpose: Recognizes a DateTimeSelect Kind Entity that is :
	--        1 -> Date
	--        2 -> LocalTime
	--        3 -> DateAndTime
	--        0 else

	Date (me) returns any Date;
	---Purpose : returns Value as a Date (Null if another type)

	LocalTime (me) returns any LocalTime;
	---Purpose : returns Value as a LocalTime (Null if another type)

	DateAndTime (me) returns any DateAndTime;
	---Purpose : returns Value as a DateAndTime (Null if another type)


end DateTimeSelect;

