-- Created on: 2010-08-27
-- Created by: Paul SUPRYATKIN
-- Copyright (c) 2010-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Localizer from OSD 

	---Purpose:  Define the locale.

is
 Create ( Category : Integer from Standard;
          Locale   : CString from Standard);
    ---Purpose: Set locale
    ---Level: Public

 Restore( me: in out );
    ---Purpose: Restore previously locale
    ---Level: Public     

 SetLocale( me: in out;
            Category : Integer from Standard;
            Locale   : CString from Standard);
    ---Purpose: Set locale
    ---Level: Public
 
 Locale( me ) 
   returns CString from Standard;
    ---Purpose: Get locale
    ---Level: Public


 Category( me ) 
   returns Integer from Standard;
    ---Purpose: Get Gategory
    ---Level: Public


fields

   myLocale        : CString from Standard; 
   myCategory      : Integer from Standard;    

end Localizer from OSD;


