-- Created on: 1993-01-09
-- Created by: CKY / Contract Toubro-Larsen ( Anand NATRAJAN )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class ExternalReferenceFile from IGESBasic  inherits IGESEntity

        ---Purpose: defines ExternalReferenceFile, Type <406> Form <12>
        --          in package IGESBasic
        --          References definitions residing in another file

uses

        HAsciiString from TCollection,
        HArray1OfHAsciiString from Interface

raises OutOfRange

is

        Create returns mutable ExternalReferenceFile;

        -- Specific Methods pertaining to the class

        Init (me : mutable; aNameArray : HArray1OfHAsciiString);
        ---Purpose : This method is used to set the fields of the class
        --           ExternalReferenceFile
        --       - aNameArray : External Reference File Names

        NbListEntries (me) returns Integer;
        ---Purpose : returns number of External Reference File Names

        Name (me; Index : Integer) returns HAsciiString from TCollection
        raises OutOfRange;
        ---Purpose : returns External Reference File Name
        -- raises exception if Index <= 0 or Index > NbListEntries()

fields

--
-- Class    : IGESBasic_ExternalReferenceFile
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class ExternalReferenceFile.
--
-- Reminder : A ExternalReferenceFile instance is defined by :
--            - External Reference File Names

        theNames : HArray1OfHAsciiString;

end ExternalReferenceFile;
