-- Created on: 1993-01-28
-- Created by: Laurent BUCHARD
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class  PrmPrmIntersection_T3Bits from IntPatch

uses Integer from Standard

is 
     
    Create (size : Integer from Standard);

    Destroy(me : in out);
    ---C++: alias ~
	 
    Add (me : in out; t : Integer from Standard);
    ---C++: inline

    Val (me ; t : Integer from Standard) returns Integer from Standard;
    ---C++: inline
   	
    Raz (me : in out; t : Integer from Standard);
    ---C++: inline

    ResetAnd (me : in  out);

    And (me : in out;
         Oth             : in out PrmPrmIntersection_T3Bits from IntPatch;
		 indiceprecedent : in out Integer from Standard)
    returns Integer from Standard;

fields
    -- ind   : Integer from Standard;
    p     : Address from Standard;
    Isize : Integer from Standard;

end PrmPrmIntersection_T3Bits;
