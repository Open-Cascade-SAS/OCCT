-- Created on: 1995-10-24
-- Created by: Mister rmi
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package PPoly 

	---Purpose: This  package  provides  persistent classes  to
	--          handle :
	--          
	--          * 3D triangular polyhedrons.
	--          
	--          * 3D polygons.
	--          
	--          * 2D polygon.

uses    PCollection,
        PColStd,
   	PColgp

is

    class Triangle;

    class Triangulation;

    class Polygon3D;

    class Polygon2D;

    class PolygonOnTriangulation;

    class HArray1OfTriangle
    instantiates HArray1 from PCollection(Triangle from PPoly);

end PPoly;
