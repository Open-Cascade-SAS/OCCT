-- Created on: 1996-01-09
-- Created by: Denis PASCAL
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



deferred class PlanarDimension from DrawDim inherits Dimension from DrawDim

	---Purpose: 

uses Face from TopoDS

is

    SetPlane (me : mutable; plane : Face from TopoDS);
    
    GetPlane (me)
    returns Face from TopoDS;


--    Point (myclass; s : Shape from TopoDS; p : in out Pnt from gp)

--    returns Boolean from Standard;    


--    Line (myclass; s : Shape from TopoDS; l : in out Lin from gp)

--    returns Boolean from Standard;    


--    Circle (myclass; s : Shape from TopoDS; c : in out Circ from gp)

--    returns Boolean from Standard;    


--    Ellipse (myclass; s : Shape from TopoDS; c : in out Elips from gp)

--    returns Boolean from Standard;


fields

    myPlane : Face from TopoDS  is protected;
    
end PlanarDimension;
