-- File:        FileName.cdl
-- Created:     Thu Jun 16 18:05:55 1994
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWFileName from RWHeaderSection

	---Purpose : Read & Write Module for FileName

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     FileName from HeaderSection

is

	Create returns RWFileName;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable FileName from HeaderSection);

	WriteStep (me; SW : in out StepWriter; ent : FileName from HeaderSection);

end RWFileName;
