-- Created on: 1993-10-29
-- Created by: Christophe MARION
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class PolyShellData from HLRAlgo inherits TShared from MMgt

uses
    Address            from Standard,
    Boolean            from Standard,
    Integer            from Standard,
    Array1OfTransient  from TColStd,
    HArray1OfTransient from TColStd,
    ListOfBPoint       from HLRAlgo

is
    Create(nbFace : Integer from Standard)
    returns mutable PolyShellData from HLRAlgo;

    UpdateGlobalMinMax(me        : mutable;
                       TotMinMax : Address from Standard)
    is static;
    
    UpdateHiding(me       : mutable;
  	         nbHiding : Integer from Standard)
    is static;

    Hiding(me) returns Boolean from Standard
	---C++: inline
    is static;

    PolyData(me : mutable) 
	---C++: return &
	---C++: inline
    returns Array1OfTransient from TColStd
    is static;

    HidingPolyData(me : mutable) 
	---C++: return &
	---C++: inline
    returns Array1OfTransient from TColStd
    is static;

    Edges(me : mutable) 
	---C++: return &
	---C++: inline
    returns ListOfBPoint from HLRAlgo
    is static;

    Indices(me : mutable) returns Address from Standard
    	---C++: inline
    is static;

fields
    myMinMax    : Integer            from Standard[2];
    myPolyg     : Array1OfTransient  from TColStd;
    myHPolHi    : HArray1OfTransient from TColStd;
    mySegList   : ListOfBPoint       from HLRAlgo;

end PolyShellData;
