-- Created on: 2003-06-04
-- Created by: Galina KULIKOVA
-- Copyright (c) 2003-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class DatumTarget from StepDimTol
inherits ShapeAspect from StepRepr

    ---Purpose: Representation of STEP entity DatumTarget

uses
    HAsciiString from TCollection,
    ProductDefinitionShape from StepRepr,
    Logical from StepData

is
    Create returns DatumTarget from StepDimTol;
	---Purpose: Empty constructor

    Init (me: mutable; aShapeAspect_Name: HAsciiString from TCollection;
                       aShapeAspect_Description: HAsciiString from TCollection;
                       aShapeAspect_OfShape: ProductDefinitionShape from StepRepr;
                       aShapeAspect_ProductDefinitional: Logical from StepData;
                       aTargetId: HAsciiString from TCollection);
	---Purpose: Initialize all fields (own and inherited)

    TargetId (me) returns HAsciiString from TCollection;
	---Purpose: Returns field TargetId
    SetTargetId (me: mutable; TargetId: HAsciiString from TCollection);
	---Purpose: Set field TargetId

fields
    theTargetId: HAsciiString from TCollection;

end DatumTarget;
