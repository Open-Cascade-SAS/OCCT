-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class ViewVolume from StepVisual 

inherits TShared from MMgt

uses

	CentralOrParallel from StepVisual, 
	CartesianPoint from StepGeom, 
	Real from Standard, 
	Boolean from Standard, 
	PlanarBox from StepVisual
is

	Create returns mutable ViewVolume;
	---Purpose: Returns a ViewVolume

	Init (me : mutable;
	      aProjectionType : CentralOrParallel from StepVisual;
	      aProjectionPoint : mutable CartesianPoint from StepGeom;
	      aViewPlaneDistance : Real from Standard;
	      aFrontPlaneDistance : Real from Standard;
	      aFrontPlaneClipping : Boolean from Standard;
	      aBackPlaneDistance : Real from Standard;
	      aBackPlaneClipping : Boolean from Standard;
	      aViewVolumeSidesClipping : Boolean from Standard;
	      aViewWindow : mutable PlanarBox from StepVisual) is virtual;

	-- Specific Methods for Field Data Access --

	SetProjectionType(me : mutable; aProjectionType : CentralOrParallel);
	ProjectionType (me) returns CentralOrParallel;
	SetProjectionPoint(me : mutable; aProjectionPoint : mutable CartesianPoint);
	ProjectionPoint (me) returns mutable CartesianPoint;
	SetViewPlaneDistance(me : mutable; aViewPlaneDistance : Real);
	ViewPlaneDistance (me) returns Real;
	SetFrontPlaneDistance(me : mutable; aFrontPlaneDistance : Real);
	FrontPlaneDistance (me) returns Real;
	SetFrontPlaneClipping(me : mutable; aFrontPlaneClipping : Boolean);
	FrontPlaneClipping (me) returns Boolean;
	SetBackPlaneDistance(me : mutable; aBackPlaneDistance : Real);
	BackPlaneDistance (me) returns Real;
	SetBackPlaneClipping(me : mutable; aBackPlaneClipping : Boolean);
	BackPlaneClipping (me) returns Boolean;
	SetViewVolumeSidesClipping(me : mutable; aViewVolumeSidesClipping : Boolean);
	ViewVolumeSidesClipping (me) returns Boolean;
	SetViewWindow(me : mutable; aViewWindow : mutable PlanarBox);
	ViewWindow (me) returns mutable PlanarBox;

fields

	projectionType : CentralOrParallel from StepVisual; -- an Enumeration
	projectionPoint : CartesianPoint from StepGeom;
	viewPlaneDistance : Real from Standard;
	frontPlaneDistance : Real from Standard;
	frontPlaneClipping : Boolean from Standard;
	backPlaneDistance : Real from Standard;
	backPlaneClipping : Boolean from Standard;
	viewVolumeSidesClipping : Boolean from Standard;
	viewWindow : PlanarBox from StepVisual;

end ViewVolume;
