-- File:	StepToGeom_MakeVectorWithMagnitude2d.cdl
-- Created:	Wed Aug  4 11:43:33 1993
-- Author:	Martine LANGLOIS
---Copyright:	 Matra Datavision 1993

class MakeVectorWithMagnitude2d from StepToGeom

    ---Purpose: This class implements the mapping between classes 
    --          Vector from StepGeom which describes a VectorWithMagnitude 
    --          from Prostep and VectorWithMagnitude from Geom2d.
  
uses 
     VectorWithMagnitude from Geom2d,
     Vector from StepGeom

is 

    Convert ( myclass; SV : Vector from StepGeom;
                       CV : out VectorWithMagnitude from Geom2d )
    returns Boolean from Standard;

end MakeVectorWithMagnitude2d;
