-- File:	Sweep_Tool.cdl
-- Created:	Wed May 26 11:50:51 1993
-- Author:	Laurent BOURESCHE
--		<lbo@phylox>
---Copyright:	 Matra Datavision 1993


deferred generic class Tool from Sweep (TheShape as any)

    ---Purpose: This  is a signature  class  describing the indexation
    --          and type analysis  services required by  the Directing
    --          and Generating Shapes of Swept Primitives.
    --          

uses

    ShapeEnum from TopAbs,
    Orientation from TopAbs

raises 

    OutOfRange from Standard

is

    Initialize(aShape: TheShape);
	---Purpose: Initialize the tool  with <aShape>.  The IndexTool
	--          must prepare an indexation for  all  the subshapes
	--          of this shape.

    NbShapes(me) returns Integer
	---Purpose: Returns the number of subshapes in the shape.
    is deferred;

    Index(me; aShape : TheShape) returns Integer
	---Purpose: Returns the index of <aShape>.
    is deferred;
    
    Shape(me; anIndex : Integer from Standard) returns TheShape
	---Purpose: Returns the Shape of index anIndex
    is deferred;
    
    Type(me; aShape : TheShape) returns ShapeEnum from TopAbs
	---Purpose: Returns the type of <aShape>.
    is deferred;
    
    Orientation(me; aShape : TheShape) returns Orientation from TopAbs
	---Purpose: Returns the Orientation of <aShape>.
    is deferred;
    
    SetOrientation(me; aShape : in out TheShape; Or : Orientation from TopAbs) 
	---Purpose: Set the Orientation of <aShape> with Or.
    is deferred;

------------------------------------------
--- Methods used for Directing Shapes only
------------------------------------------

    HasFirstVertex(me) returns Boolean from Standard
	---Purpose: Returns true if there is a First Vertex in the Shape.
    is deferred;

    HasLastVertex(me) returns Boolean from Standard
	---Purpose: Returns true if there is a Last Vertex in the Shape.
    is deferred;

    FirstVertex(me) returns TheShape
	---Purpose: Returns the first vertex.
    is deferred;

    LastVertex(me) returns TheShape
	---Purpose: Returns the last vertex.
    is deferred;

end Tool from Sweep;
