-- Created on: 1993-03-23
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class LoopSet from TopOpeBRepBuild

uses

    Loop                     from TopOpeBRepBuild,
    ListOfLoop               from TopOpeBRepBuild,
    ListIteratorOfListOfLoop from TopOpeBRepBuild

is
    
    Create returns LoopSet;
    
    Delete(me:out) is virtual;
    ---C++: alias "Standard_EXPORT virtual ~TopOpeBRepBuild_LoopSet(){Delete() ; }"
    
    -- filling : append loops (shapes,blocks) in list
    ChangeListOfLoop(me : in out) returns ListOfLoop is static;
    ---C++: return &

    -- exploration of the loops
    InitLoop(me : in out) is virtual;
    MoreLoop(me) returns Boolean is virtual;
    NextLoop(me : in out) is virtual;
    Loop(me) returns Loop from TopOpeBRepBuild is virtual;
    ---C++: return const &
    
fields

    myListOfLoop : ListOfLoop;
    myLoopIterator : ListIteratorOfListOfLoop;
    myLoopIndex : Integer from Standard;
    myNbLoop : Integer from Standard;
    
end LoopSet from TopOpeBRepBuild;
