-- Created on: 1998-08-26
-- Created by: Julia GERASIMOVA
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MakeFilling from BRepOffsetAPI inherits MakeShape from BRepBuilderAPI

	---Purpose: N-Side Filling
	--  This algorithm avoids to build a face from:
	--  * a set of edges defining the bounds of the face and some
	--    constraints the surface of the face has to satisfy
	--  * a set of edges and points defining some constraints
	--    the support surface has to satisfy
	--  * an initial surface to deform for satisfying the constraints
	--  * a set of parameters to control the constraints.
	--
	--  The support surface of the face is computed by deformation
	--  of the initial surface in order to satisfy the given constraints.
	--  The set of bounding edges defines the wire of the face.
	--
	--  If no initial surface is given, the algorithm computes it
	--  automatically.
	--  If the set of edges is not connected (Free constraint)
	--  missing edges are automatically computed.
	--
	--  Limitations:
	--  * If some constraints are not compatible
	--    The algorithm does not take them into account.
	--    So the constraints will not be satisfyed in an area containing
	--    the incompatibilitries.
	--  * The constraints defining the bound of the face have to be
	--    entered in order to have a continuous wire.
	--
	--  Other Applications:
	--  * Deformation of a face to satisfy internal constraints
	--  * Deformation of a face to improve Gi continuity with
	--    connected faces
	
	---Level: Advanced

uses
    Shape from TopoDS,
    Edge  from TopoDS,
    Face  from TopoDS,
    Pnt   from gp,
    Shape from GeomAbs,
    ListOfShape from TopTools,
    Filling from BRepFill

raises
    NotDone,
    OutOfRange,
    ConstructionError

is
    Create( Degree      : Integer from Standard = 3;
    	    NbPtsOnCur  : Integer from Standard = 15;
	    NbIter      : Integer from Standard = 2;
	    Anisotropie : Boolean from Standard = Standard_False;
	    Tol2d       : Real    from Standard = 0.00001;
	    Tol3d       : Real    from Standard = 0.0001;
	    TolAng      : Real    from Standard = 0.01;
	    TolCurv     : Real    from Standard = 0.1;
	    MaxDeg      : Integer from Standard = 8;
	    MaxSegments : Integer from Standard = 9 )
    	---Purpose: Constructs a wire filling object defined by
    	-- - the energy minimizing criterion Degree
    	-- - the number of points on the curve NbPntsOnCur
    	-- - the number of iterations NbIter
    	-- - the Boolean Anisotropie
    	-- - the 2D tolerance Tol2d
    	-- - the 3D tolerance Tol3d
    	-- - the angular tolerance TolAng
    	-- - the tolerance for curvature TolCur
    	-- - the highest polynomial degree MaxDeg
    	-- - the greatest number of segments MaxSeg.
    	-- If the Boolean Anistropie is true, the algorithm's
    	-- performance is better in cases where the ratio of the
    	-- length U and the length V indicate a great difference
    	-- between the two. In other words, when the surface is, for
    	-- example, extremely long.
         returns MakeFilling from BRepOffsetAPI;
    
    
    SetConstrParam( me : in out; Tol2d   : Real    from Standard = 0.00001;
    	    	    	    	 Tol3d   : Real    from Standard = 0.0001;
				 TolAng  : Real    from Standard = 0.01;
				 TolCurv : Real    from Standard = 0.1 );
    	---Purpose: Sets the values of Tolerances used to control the constraint.
    	--	Tol2d:
    	--	Tol3d:   it is the maximum distance allowed between the support surface
    	--	         and the constraints
    	--	TolAng:  it is the maximum angle allowed between the normal of the surface
    	--	         and the constraints
    	--	TolCurv: it is the maximum difference of curvature allowed between
    	--	         the surface and the constraint
    
    SetResolParam( me : in out; Degree      : Integer from Standard = 3;
    	    	    	    	NbPtsOnCur  : Integer from Standard = 15;
				NbIter      : Integer from Standard = 2;
				Anisotropie : Boolean from Standard = Standard_False );
    	---Purpose: Sets the parameters used for resolution.
    	--	The default values of these parameters have been chosen for a good
    	--	ratio quality/performance.
    	--	Degree:      it is the order of energy criterion to minimize for computing
    	--	             the deformation of the surface.
    	--	             The default value is 3
    	--	             The recommanded value is i+2 where i is the maximum order of the
    	--	             constraints.
    	--	NbPtsOnCur:  it is the average number of points for discretisation
    	--	             of the edges.
    	--	NbIter:      it is the maximum number of iterations of the process.
    	--	             For each iteration the number of discretisation points is
    	--	             increased.
    	--	Anisotropie: 
    
    SetApproxParam( me : in out; MaxDeg      : Integer from Standard = 8;
				 MaxSegments : Integer from Standard = 9 );
    	---Purpose: Sets the parameters used to approximate the filling
    	-- surface. These include:
    	-- - MaxDeg - the highest degree which the polynomial
    	--   defining the filling surface can have
    	-- - MaxSegments - the greatest number of segments
    	--   which the filling surface can have.
    
    
    LoadInitSurface( me : in out; Surf : Face from TopoDS );
    	---Purpose: Loads the initial surface Surf to
    	-- begin the construction of the surface.
    	-- This optional function is useful if the surface resulting from
    	-- construction for the algorithm is likely to be complex.
    	-- The support surface of the face under construction is computed by a
    	-- deformation of Surf which satisfies the given constraints.
    	-- The set of bounding edges defines the wire of the face.
    	-- If no initial surface is given, the algorithm computes it
    	-- automatically. If the set of edges is not connected (Free constraint),
    	-- missing edges are automatically computed.
    
    
    Add( me : in out; Constr : Edge from TopoDS;
    	    	      Order  : Shape from GeomAbs;
		      IsBound : Boolean from Standard = Standard_True )
    returns Integer from Standard
    	---Purpose: Adds a new constraint which also defines an edge of the wire
    	--	        of the face
    	--	Order: Order of the constraint:
    	--	       GeomAbs_C0 : the surface has to pass by 3D representation
    	--	                    of the edge
    	--	       GeomAbs_G1 : the surface has to pass by 3D representation
    	--	                    of the edge and to respect tangency with the first
    	--	                    face of the edge
    	--	       GeomAbs_G2 : the surface has to pass by 3D representation
    	--	                    of the edge and to respect tangency and curvature
    	--	                    with the first face of the edge.
    	--  Raises ConstructionError if the edge has no representation on a face and Order is
    	-- GeomAbs_G1 or GeomAbs_G2.
    raises ConstructionError from Standard;
   
    
    Add( me : in out; Constr  : Edge from TopoDS;
    	    	      Support : Face from TopoDS;
		      Order   : Shape from GeomAbs;
		      IsBound : Boolean from Standard = Standard_True )
    returns Integer from Standard
    	---Purpose: Adds a new constraint which also defines an edge of the wire
    	--	        of the face
    	--	Order: Order of the constraint:
    	--	       GeomAbs_C0 : the surface has to pass by 3D representation
    	--	                    of the edge
    	--	       GeomAbs_G1 : the surface has to pass by 3D representation
    	--	                    of the edge and to respect tangency with the
    	--	                    given face
    	--	       GeomAbs_G2 : the surface has to pass by 3D representation
    	--	                    of the edge and to respect tangency and curvature
    	--                    with the given face.
	-- Raises ConstructionError if the edge has no 2d representation on the given face
    raises ConstructionError from Standard;
    
    Add( me : in out; Support : Face from TopoDS;
		      Order   : Shape from GeomAbs )
    returns Integer from Standard;
    	---Purpose: Adds a free constraint on a face. The corresponding edge has to
    	--	be automatically recomputed. It is always a bound.
    
    Add( me : in out; Point : Pnt from gp )
    returns Integer from Standard;
    	---Purpose: Adds a punctual constraint.
    
    Add( me : in out; U, V    : Real from Standard;
    	    	      Support : Face from TopoDS;
		      Order   : Shape from GeomAbs )
    returns Integer from Standard;
    	---Purpose: Adds a punctual constraint.
    

    Build( me : in out )
    	---Purpose: Builds the resulting faces
    is redefined;
    
    IsDone(me) returns Boolean from Standard
    is redefined;
    	--- Purpose: Tests whether computation of the filling plate has been completed.
    
    Generated (me: in out; S : Shape from TopoDS)
    	---Purpose: Returns the list of shapes generated from the
    	--          shape <S>. 
        ---C++: return const & 
        ---Level: Public
    returns ListOfShape from TopTools
    is redefined;     
   
    G0Error(me) returns Real from Standard;
    	--- Purpose: Returns the maximum distance between the result and
    	-- the constraints. This is set at construction time.
    
    G1Error(me) returns Real from Standard;
    	---Purpose: Returns the maximum angle between the result and the
    	-- constraints. This is set at construction time. 
    
    G2Error(me) returns Real from Standard;
    	---Purpose: Returns the maximum angle between the result and the
    	-- constraints. This is set at construction time. 
    
    G0Error( me : in out; Index : Integer from Standard ) returns Real from Standard;
    	---Purpose: Returns the maximum distance attained between the
    	-- result and the constraint Index. This is set at construction time.
    
    G1Error( me : in out; Index : Integer from Standard ) returns Real from Standard;
    	---Purpose: Returns the maximum angle between the result and the
    	-- constraints. This is set at construction time. 
    
    G2Error( me : in out; Index : Integer from Standard ) returns Real from Standard;
    	---Purpose: Returns the greatest difference in curvature found
    	-- between the result and the constraint Index.
    
fields

    myFilling : Filling from BRepFill;

end MakeFilling;
