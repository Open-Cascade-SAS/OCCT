-- Created on: 1992-11-18
-- Created by: Christian CAILLET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class SelectEntityNumber  from IFSelect  inherits SelectBase

    ---Purpose : A SelectEntityNumber gets in an InterfaceModel (through a
    --           Graph), the Entity which has a specified Number (its rank of
    --           adding into the Model) : there can be zero (if none) or one.
    --           The Number is not directly defined as an Integer, but as a
    --           Parameter, which can be externally controled

uses AsciiString from TCollection, EntityIterator, Graph, IntParam

is

    Create  returns mutable SelectEntityNumber;
    ---Purpose : Creates a SelectEntityNumber, initially with no specified Number

    SetNumber (me : mutable; num : mutable IntParam);
    ---Purpose : Sets Entity Number to be taken (initially, none is set : 0)

    Number (me) returns mutable IntParam;
    ---Purpose : Returns specified Number (as a Parameter)

    RootResult (me; G : Graph) returns EntityIterator;
    ---Purpose : Returns the list of selected entities : the Entity having the
    --           specified Number (this result assures naturally uniqueness)

    Label (me) returns AsciiString from TCollection;
    ---Purpose : Returns a text defining the criterium : "Entity Number ..."

fields

    thenum : IntParam;

end SelectEntityNumber;
