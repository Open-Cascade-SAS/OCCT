-- File:	GeomToStep_MakeSweptSurface.cdl
-- Created:	Tue Jun 22 14:40:20 1993
-- Author:	Martine LANGLOIS
--		<mla@mastox>
---Copyright:	 Matra Datavision 1993

class MakeSweptSurface from GeomToStep inherits Root from GeomToStep

    ---Purpose: This class implements the mapping between classes 
    --          SweptSurface from Geom and the class SweptSurface from 
    --          StepGeom which describes a SweptSurface from prostep.
    --          As SweptSurface is an abstract SweptSurface this class 
    --          is an access to the sub-class required.
  
uses SweptSurface from Geom,
     SweptSurface from StepGeom
     
raises NotDone from StdFail
     
is 

Create ( S : SweptSurface from Geom ) returns MakeSweptSurface;

Value (me) returns SweptSurface from StepGeom
    raises NotDone
    is static;
    ---C++: return const&

fields

    theSweptSurface : SweptSurface from StepGeom;
    	-- The solution from StepGeom
    	
end MakeSweptSurface;



