-- Created on: 1994-09-15
-- Created by: Bruno DUMORTIER
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class ProjectOnSurface from ProjLib 

uses

    HCurve       from Adaptor3d,
    HSurface     from Adaptor3d,
    BSplineCurve from Geom

is

    Create 
    	---Purpose:  Create an empty projector.
    returns ProjectOnSurface from ProjLib;
    

    Create( S  : HSurface from Adaptor3d)
    	---Purpose: Create a projector normaly to the surface <S>.
    returns ProjectOnSurface from ProjLib;

    Delete(me:out) is virtual;
    ---C++: alias "Standard_EXPORT virtual ~ProjLib_ProjectOnSurface(){Delete() ; }"
    
    Load(me : in out; S : HSurface from Adaptor3d)
	---Purpose: Set the Surface to <S>.
	--          To compute the projection, you have to Load the Curve.
    is static;
    
    Load(me : in out; C : HCurve from Adaptor3d; Tolerance : Real)
	---Purpose: Compute the projection of the curve <C> on the Surface.
    is static;

    IsDone(me) returns Boolean ;
    
    BSpline(me) returns BSplineCurve from Geom  
    is static ;

fields

    myCurve      : HCurve   from Adaptor3d ;
    mySurface    : HSurface from Adaptor3d ;
    myTolerance  : Real ;
    myIsDone     : Boolean ;
    myResult     : BSplineCurve from Geom ;

end ProjectOnSurface;
