-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SecurityClassification from StepBasic 

inherits TShared from MMgt

uses

	HAsciiString from TCollection, 
	SecurityClassificationLevel from StepBasic
is

	Create returns mutable SecurityClassification;
	---Purpose: Returns a SecurityClassification

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aPurpose : mutable HAsciiString from TCollection;
	      aSecurityLevel : mutable SecurityClassificationLevel from StepBasic) is virtual;

	-- Specific Methods for Field Data Access --

	SetName(me : mutable; aName : mutable HAsciiString);
	Name (me) returns mutable HAsciiString;
	SetPurpose(me : mutable; aPurpose : mutable HAsciiString);
	Purpose (me) returns mutable HAsciiString;
	SetSecurityLevel(me : mutable; aSecurityLevel : mutable SecurityClassificationLevel);
	SecurityLevel (me) returns mutable SecurityClassificationLevel;

fields

	name : HAsciiString from TCollection;
	purpose : HAsciiString from TCollection;
	securityLevel : SecurityClassificationLevel from StepBasic;

end SecurityClassification;
