-- Created on: 1993-03-10
-- Created by: Philippe DAUTRY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package TColgp  


        ---Purpose :   This package  provides  standard and frequently
    	-- used instantiations of generic classes from the
    	-- TCollection package with geometric objects from the gp package.     

uses TCollection, TColStd, gp

is



    -- Array1 of 2D objects.

  imported Array1OfCirc2d;
  imported Array1OfDir2d;
  imported Array1OfLin2d;
  imported Array1OfPnt2d;
  imported Array1OfVec2d;
  imported Array1OfXY;


    -- Array1 of 3D objects.

  imported Array1OfDir;
  imported Array1OfPnt;
  imported Array1OfVec;
  imported Array1OfXYZ;


    -- Array2 of 2D objects.

  imported Array2OfCirc2d;
  imported Array2OfDir2d;
  imported Array2OfLin2d;
  imported Array2OfPnt2d;
  imported Array2OfVec2d;
  imported Array2OfXY;


    -- Array2 of 3D objects.

  imported Array2OfDir;
  imported Array2OfPnt;
  imported Array2OfVec;
  imported Array2OfXYZ;


    -- HArray1 of 2D objects.

  imported transient class HArray1OfCirc2d;
  imported transient class HArray1OfDir2d;
  imported transient class HArray1OfLin2d;
  imported transient class HArray1OfPnt2d;
  imported transient class HArray1OfVec2d;
  imported transient class HArray1OfXY;


    -- HArray1 of 3D objects.

  imported transient class HArray1OfDir;
  imported transient class HArray1OfPnt;
  imported transient class HArray1OfVec;
  imported transient class HArray1OfXYZ;


    -- HArray2 of 2D objects.

  imported transient class HArray2OfCirc2d;
  imported transient class HArray2OfDir2d;
  imported transient class HArray2OfLin2d;
  imported transient class HArray2OfPnt2d;
  imported transient class HArray2OfVec2d;
  imported transient class HArray2OfXY;


    -- HArray2 of 3D objects.

  imported transient class HArray2OfDir;
  imported transient class HArray2OfPnt;
  imported transient class HArray2OfVec;
  imported transient class HArray2OfXYZ;


    -- Sequences of 3D objects.

  imported SequenceOfDir;
  imported SequenceOfPnt;
  imported SequenceOfVec;
  imported SequenceOfXYZ;
  imported SequenceOfAx1;


    -- HSequences of 3D objects.

  imported transient class HSequenceOfDir;
  imported transient class HSequenceOfPnt;

  imported transient class HSequenceOfVec;

  imported transient class HSequenceOfXYZ;


    -- Sequences of 2D objects.

  imported SequenceOfDir2d;
  imported SequenceOfPnt2d;
  imported SequenceOfVec2d;
  imported SequenceOfXY;
  imported SequenceOfArray1OfPnt2d;


    -- HSequences of 2D objects.

  imported transient class HSequenceOfDir2d;
  imported transient class HSequenceOfPnt2d;
  imported transient class HSequenceOfVec2d;
  imported transient class HSequenceOfXY;

end TColgp;
