-- Created on: 1997-04-29
-- Created by: Stagiaire Francois DUMONT
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class CompCurveToBSplineCurve from Geom2dConvert 

	    ---Purpose: This algorithm converts and concat several curve in an BSplineCurve

uses
 ParameterisationType from Convert,
 BoundedCurve from Geom2d,
 BSplineCurve from Geom2d

--raises

is

    Create(Parameterisation : ParameterisationType from Convert = Convert_TgtThetaOver2);
    ---Purpose: Initialize the algorithme
    --        - Parameterisation is used to convert

    Create (BasisCurve : BoundedCurve from Geom2d; 
     	    Parameterisation : ParameterisationType from Convert 
    	    	       =  Convert_TgtThetaOver2)
	    ---Purpose: Initialize the algorithme with one curve
	    --        - Parameterisation is used to convert 
    returns CompCurveToBSplineCurve;

    Add (me : in out; 
         NewCurve :  BoundedCurve from Geom2d;
         Tolerance:  Real from Standard;
         After      : Boolean from Standard = Standard_False)
	    ---Purpose: Append a curve in the BSpline
	    --          Return False if the curve is not G0 with the BSplineCurve.
	    --          Tolerance is used to check continuity and decrease 
	    --          Multiplicty at the common Knot 
	    --          After is usefull if BasisCurve is a closed curve .
    returns Boolean;
       
    
    Add (me : in out; 
         FirstCurve : in out BSplineCurve from Geom2d;
    	 SecondCurve: in out BSplineCurve from Geom2d;
         After      : Boolean from Standard)
	    ---Purpose: Concat two BSplineCurves.
    	is private;    
    
    BSplineCurve(me) returns BSplineCurve from Geom2d;

    Clear(me : in out);
    ---Purpose: Clear result curve

fields
 myCurve :  BSplineCurve from Geom2d;
 myTol   :  Real;
 myType  :  ParameterisationType from Convert;

end CompCurveToBSplineCurve;
