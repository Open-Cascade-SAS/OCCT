-- File:	QAAlcatel.cdl
-- Created:	Tue May 21 19:15:02 2002
-- Author:	QA Admin
--		<qa@russox>
---Copyright:	 Matra Datavision 2002

package QAAlcatel
     uses Draw
is
    Commands(DI : in out Interpretor from Draw);
end;
