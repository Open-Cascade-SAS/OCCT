-- File:	BinMNaming_NamingDriver.cdl
-- Created:	Thu May 13 16:51:27 2004
-- Author:	Sergey ZARITCHNY <szy@opencascade.com>
-- Copyright:	Open CasCade S.A. 2004

class NamingDriver from BinMNaming inherits ADriver from BinMDF

	---Purpose: Naming  Attribute Driver.

uses
    SRelocationTable from BinObjMgt,
    RRelocationTable from BinObjMgt,
    Persistent       from BinObjMgt,
    MessageDriver    from CDM,
    Attribute        from TDF


is
    Create (theMessageDriver:MessageDriver from CDM)
        returns mutable NamingDriver from BinMNaming;

    NewEmpty (me)  returns mutable Attribute from TDF;

    Paste(me; Source     : Persistent from BinObjMgt;
              Target     : mutable Attribute from TDF;
              RelocTable : out RRelocationTable from BinObjMgt)
        returns Boolean from Standard;

    Paste(me; Source     : Attribute from TDF;
              Target     : in out Persistent from BinObjMgt;
              RelocTable : out SRelocationTable from BinObjMgt);
    

end NamedShapeDriver;

