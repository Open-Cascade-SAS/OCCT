-- File:	BRepPrimAPI_MakeCylinder.cdl
-- Created:	Wed Jul 21 16:07:20 1993
-- Author:	Remi LEQUETTE
--		<rle@nonox>
---Copyright:	 Matra Datavision 1993


class MakeCylinder from BRepPrimAPI  inherits MakeOneAxis from BRepPrimAPI

	---Purpose: Describes functions to build cylinders or portions of  cylinders.
    	-- A MakeCylinder object provides a framework for:
    	-- -   defining the construction of a cylinder,
    	-- -   implementing the construction algorithm, and
    	-- -   consulting the result.

uses
    Ax2      from gp,
    Cylinder from BRepPrim,
    OneAxis  from BRepPrim

raises
    DomainError from Standard
    
is

    Create(R, H : Real)
    returns MakeCylinder from BRepPrimAPI
	---Purpose: Make a cylinder of radius R and length H.
	---Level: Public
    raises
    	DomainError from Standard; -- if R or H <= Precision::Confusion()

    Create(R, H, Angle : Real)
    returns MakeCylinder from BRepPrimAPI
	---Purpose: Make a cylinder   of  radius R  and  length H with
	--          angle  H.
	---Level: Public
    raises
    	DomainError from Standard; -- if R or H <= Precision::Confusion()

    Create(Axes : Ax2 from gp; R, H : Real)
    returns MakeCylinder from BRepPrimAPI
	---Purpose: Make a cylinder of radius R and length H.
	---Level: Public
    raises
    	DomainError from Standard; -- if R or H <= Precision::Confusion()

    Create(Axes : Ax2 from gp; R, H, Angle : Real)
    returns MakeCylinder from BRepPrimAPI
	---Purpose: Make a cylinder   of  radius R  and  length H with
	--          angle  H.
	---Level: Public
    raises
    	DomainError from Standard; -- if R or H <= Precision::Confusion()

    	---Purpose: Constructs
    	-- -   a cylinder of radius R and height H, or
    	-- -   a portion of cylinder of radius R and height H, and of
    	--   the angle Angle defining the missing portion of the cylinder.    
    	-- The cylinder is constructed about the "Z Axis" of either:
    	-- -   the global coordinate system, or
    	-- -   the local coordinate system Axes.
    	-- It is limited in this coordinate system as follows:
    	-- -   in the v parametric direction (the Z axis), by the two
    	--   parameter values 0 and H,
    	-- -   and in the u parametric direction (the rotation angle
    	--   around the Z Axis), in the case of a portion of a
    	--   cylinder, by the two parameter values 0 and Angle.
    	--   Angle is given in radians.
    	-- The resulting shape is composed of:
    	-- -   a lateral cylindrical face,
    	-- -   two planar faces in the planes z = 0 and z = H
    	--   (in the case of a complete cylinder, these faces are circles), and
    	-- -   in case of a portion of a cylinder, two additional
    	--   planar faces to close the shape.(two rectangles in the
    	--   planes u = 0 and u = Angle).
    	-- Exceptions Standard_DomainError if:
    	-- -   R is less than or equal to Precision::Confusion(), or
    	-- -   H is less than or equal to Precision::Confusion().
        
    OneAxis(me : in out) returns Address;
	---Purpose: Returns the algorithm.
	---Level: Advanced

    Cylinder(me : in out) returns Cylinder from BRepPrim
	---Purpose: Returns the algorithm.
	--          
	---C++: return &
	---Level: Public 
    is static;

fields

    myCylinder : Cylinder from BRepPrim;

end MakeCylinder;
