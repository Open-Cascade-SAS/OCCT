-- Created by: Peter KURNEV
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package BOPTools 

        ---Purpose: 

uses
    gp,  
    Bnd,
    TopAbs, 
    Geom,   
    Geom2d,
    GeomAPI, 
    BRepClass3d,
    TopoDS, 
    TopTools, 
    IntTools,   
    ProjLib,
    --                 
    BOPCol, 
    BOPInt 
is 

    -- 
    -- classes
    -- 
    class ShapeSet; 
    class EdgeSet; 
    class AlgoTools; 
    class Set; 
    class SetMapHasher;  
    class AlgoTools2D; 
    class AlgoTools3D;
    -- 
    imported MapOfSet;
    imported DataMapOfShapeSet;
    --
    -- primitives
    --
    imported ListOfShapeSet from BOPTools;
    imported ListOfEdgeSet from BOPTools;
    imported ConnexityBlock from BOPTools;
    imported ListOfConnexityBlock from BOPTools;
    imported CoupleOfShape from BOPTools;
    imported ListOfCoupleOfShape from BOPTools;
    --
    --  static methods 
    -- 
    MapShapes(S : Shape from TopoDS;
                  M : in out MapOfShape from BOPCol); 
               
    MapShapes(S : Shape from TopoDS;
                  M : in out IndexedMapOfShape from BOPCol); 
              
    MapShapes(S : Shape from TopoDS;
                  T : ShapeEnum from TopAbs;
                  M : in out IndexedMapOfShape from BOPCol);
          

    MapShapesAndAncestors
            (S  : Shape from TopoDS;
             TS : ShapeEnum from TopAbs;
         TA : ShapeEnum from TopAbs;
         M  : in out IndexedDataMapOfShapeListOfShape from BOPCol);
    
end BOPTools;
