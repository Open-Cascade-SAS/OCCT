-- Created on: 1993-02-22
-- Created by: Philippe DAUTRY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package PGeom 

        ---Purpose :  This  package contains   the definition   of the
        --         geometric persistent objects such as point, vector,
        --         axis placement, curves, surfaces.
        --  
        --  All these entities are defined in 3D space.
        --  This package gives the possibility :
        --    . to create geometric objects with given or default field values,
        --    . to set field values,
        --    . to get field values.


uses PColStd, gp, PColgp, GeomAbs

is


  class Transformation from PGeom;


  deferred class Geometry from PGeom;


     deferred class Point from PGeom;
              class  CartesianPoint from PGeom;


     deferred class Vector from PGeom;
              class Direction from PGeom;
              class VectorWithMagnitude from PGeom;
     

     deferred class AxisPlacement from PGeom;
              class Axis1Placement from PGeom;
              class Axis2Placement from PGeom;


     deferred class Curve from PGeom;

              class Line from PGeom;

              deferred class Conic from PGeom;
                       class Circle from PGeom;
                       class Ellipse from PGeom;
                       class Hyperbola from PGeom;
                       class Parabola from PGeom;

              deferred class BoundedCurve from PGeom;
                       class BezierCurve from PGeom;
                       class BSplineCurve from PGeom;
                       class TrimmedCurve from PGeom;

              class  OffsetCurve from PGeom;


     deferred class Surface from PGeom;

              deferred class ElementarySurface from PGeom;
                       class Plane from PGeom;
                       class ConicalSurface from PGeom;
                       class CylindricalSurface from PGeom;
                       class SphericalSurface from PGeom;
                       class ToroidalSurface from PGeom;

              deferred class SweptSurface from PGeom;
                       class SurfaceOfLinearExtrusion from PGeom;
                       class SurfaceOfRevolution from PGeom;

              deferred class BoundedSurface from PGeom;
                       class BezierSurface from PGeom;
                       class BSplineSurface from PGeom;
                       class RectangularTrimmedSurface from PGeom;

              
              class OffsetSurface from PGeom;


end PGeom;
