-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ProductRelatedProductCategory from StepBasic 

inherits ProductCategory from StepBasic 

uses

	HArray1OfProduct from StepBasic, 
	Product from StepBasic, 
	HAsciiString from TCollection, 
	Boolean from Standard
is

	Create returns mutable ProductRelatedProductCategory;
	---Purpose: Returns a ProductRelatedProductCategory


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      hasAdescription : Boolean from Standard;
	      aDescription : mutable HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      hasAdescription : Boolean from Standard;
	      aDescription : mutable HAsciiString from TCollection;
	      aProducts : mutable HArray1OfProduct from StepBasic) is virtual;

	-- Specific Methods for Field Data Access --

	SetProducts(me : mutable; aProducts : mutable HArray1OfProduct);
	Products (me) returns mutable HArray1OfProduct;
	ProductsValue (me; num : Integer) returns mutable Product;
	NbProducts (me) returns Integer;

fields

	products : HArray1OfProduct from StepBasic;

end ProductRelatedProductCategory;
