-- File:        CartesianPoint.cdl
-- Created:     Fri Dec  1 11:11:16 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class CartesianPoint from StepGeom 

inherits Point from StepGeom 

uses

	HArray1OfReal from TColStd, 
	Real from Standard, 
	HAsciiString from TCollection
is

	Create returns mutable CartesianPoint;
	---Purpose: Returns a CartesianPoint


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aCoordinates : mutable HArray1OfReal from TColStd) is virtual;

    	Init2D (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      X,Y : Real);

    	Init3D (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      X,Y,Z : Real);

	-- Specific Methods for Field Data Access --

	SetCoordinates(me : mutable; aCoordinates : mutable HArray1OfReal);
	Coordinates (me) returns mutable HArray1OfReal;
	CoordinatesValue (me; num : Integer) returns Real;
	NbCoordinates (me) returns Integer;

fields

    nbcoord : Integer; -- optimised formula
    coords  : Real[3];
--	coordinates : HArray1OfReal from TColStd;

end CartesianPoint;
