-- Created on: 2001-03-07
-- Created by: Peter KURNEV
-- Copyright (c) 2001-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class PaveBlockIterator from BOPTools 

	---Purpose: 
        ---         class providing iterations for PaveSet to   
        ---         have the right order of paves along the edge           	 
	--- 
uses
    PaveSet from BOPTools, 
    CArray1OfPave from BOPTools, 
    PaveBlock from BOPTools 

is 
    Create 
    	returns PaveBlockIterator from BOPTools; 
    	---Purpose:  
    	--- Empty constructor 
    	---
    Create (aEdge   :  Integer from Standard; 
            aPaveSet:  PaveSet from BOPTools)
    	returns PaveBlockIterator from BOPTools; 
    	---Purpose:  
    	--- Constructor 
    	--- aEdge     -   DS-index of the edge	 
    	--- aPaveSet  -   a set of paves for the edge	  
    	---
    Initialize(me:out;aEdge   :  Integer from Standard; 
                      aPaveSet:  PaveSet from BOPTools); 
    	---Purpose:  
    	--- Resets the iterator on the PaveSet <aPaveSet> 
    	---
    More(me) 
    	returns  Boolean from Standard; 
    	---Purpose:  
    	--- Returns True if there is a current Pave in 
    	--- the iteration. 
    	---
    Next(me:out); 
    	---Purpose: 
    	--- Moves to the next Pave in the PaveSet 
    	---
    Value(me:out) 
    	returns PaveBlock from BOPTools; 
    	---C++:  return &	
    	---Purpose:  
    	--- Returns the current Pave 
    	---
fields 
    myEdge     : Integer from Standard; 
    myIndex    : Integer from Standard;   
    myPaveSet  : PaveSet from BOPTools; 
    myPaves    : CArray1OfPave from BOPTools;      
    myPaveBlock: PaveBlock from BOPTools;  
    
end PaveBlockIterator;
