-- File:	StepToGeom_MakeConic2d.cdl
-- Created:	Fri Aug 26 11:36:35 1994
-- Author:	Frederic MAUPAS
---Copyright:	 Matra Datavision 1994

class MakeConic2d from StepToGeom

    ---Purpose: This class implements the mapping between classes 
    --          Conic from StepGeom
    --          which describes a Conic from prostep and Conic from Geom2d.
    --          As Conic is an abstract class
    --          this class is an access to the sub-class required.
  
uses Conic from Geom2d,
     Conic from StepGeom
     
is 

    Convert ( myclass; SC : Conic from StepGeom;
                       CC : out Conic from Geom2d )
    returns Boolean from Standard;

end MakeConic2d;
