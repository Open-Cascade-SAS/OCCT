-- Created on: 1996-04-10
-- Created by: Joelle CHAUVET
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Modified:	Mon Dec  9 10:30:56 1996
--    by:	Joelle CHAUVET
--		G1135 : Empty constructor


class Network from AdvApp2Var

uses

    Boolean,Integer,Real from Standard,
    SequenceOfReal,HArray1OfReal from TColStd,
    IsoType from GeomAbs,
    Patch, SequenceOfPatch, Framework from AdvApp2Var

raises NoSuchObject from Standard 

is
    Create returns Network;
    Create(Net : SequenceOfPatch; TheU,TheV : SequenceOfReal) returns Network;
    FirstNotApprox(me; Index :  out Integer)
    ---Purpose: search the Index of the first Patch not approximated,
    --          if all Patches are approximated Standard_False is returned
    returns Boolean; 
    ChangePatch(me: in out; Index : Integer) 
    ---C++: alias operator()
    ---C++: return &
    ---C++: inline
    returns Patch;
    UpdateInU(me: in out; CuttingValue : Real);
    UpdateInV(me: in out; CuttingValue : Real);
    SameDegree(me : in out; iu, iv : Integer; ncfu, ncfv : out Integer);
    NbPatch(me) returns Integer;
    NbPatchInU(me) returns Integer;
    NbPatchInV(me) returns Integer;
    UParameter(me; Index : Integer) returns Real;
    VParameter(me; Index : Integer) returns Real;
    Patch(me; UIndex, VIndex : Integer) 
    ---C++: alias operator()
    ---C++: return const &
    ---C++: inline
    returns Patch;
    

fields

    myNet         : SequenceOfPatch;
    myUParameters : SequenceOfReal;
    myVParameters : SequenceOfReal;

end Network;

