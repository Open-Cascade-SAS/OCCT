-- Created on: 1998-09-22
-- Created by: Philippe MANGINGeomLib_PolyFunc.c
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



private  class PolyFunc from GeomLib inherits  FunctionWithDerivative from math

	---Purpose: Polynomial  Function        

uses 
  Vector  from  math

is 
 
    Create(Coeffs:Vector) returns  PolyFunc from GeomLib;  
    
    Value(me: in out; X: Real; F: out Real)
        ---Purpose: computes the value <F>of the function for the variable <X>.
    	--          Returns True if the calculation were successfully done, 
    	--          False otherwise.

    returns Boolean
    is redefined;
 
    Derivative(me: in out; X: Real; D: out Real)
         ---Purpose: computes the derivative <D> of the function 
         --          for the variable <X>.
    	--           Returns True if the calculation were successfully done, 
    	--           False otherwise.

    returns Boolean
    is redefined;    

    Values(me: in out; X: Real; F, D: out Real)
    	---Purpose: computes the value <F> and the derivative <D> of the 
    	--          function for the variable <X>.
    	--          Returns True if the calculation were successfully done,
    	--          False otherwise.

    returns Boolean
    is redefined; 
    
fields 
  myCoeffs  :  Vector;

end PolyFunc;
