-- Created on: 1993-04-13
-- Created by: Gerard GRAS
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class SetOfPolylines from Graphic2d inherits Line from Graphic2d

	---Version:

	---Purpose: The primitive SetOfPolylines
        --  Warning: This primitive must be use as possible for to insure 
	--	   that the sets is drawn correctly when the line type or
	--	   line width attrib is not SOLID and 1 pixel for the set.
        --         NOTE: than the method PickedIndex() permits to known
        --              the last picked polyline and segment in the set.
	---References:

uses
	Drawer			from Graphic2d,
	GraphicObject		from Graphic2d,
	Length			from Quantity,
	SequenceOfPolyline	from Graphic2d,
	FStream			from Aspect,
	IFStream		from Aspect



raises
	OutOfRange from Standard

is
	-------------------------
	-- Category: Constructors
	-------------------------

	Create (aGraphicObject: GraphicObject from Graphic2d)
	returns mutable SetOfPolylines from Graphic2d;
	---Level: Public
	---Purpose: Creates an empty set of polylines in the graphic 
	--         object <aGraphicObject>.
	---Category: Constructors

	Add(me : mutable; X, Y: Length from Quantity;
			  NewPolyline: Boolean from Standard = Standard_False);
	---Level: Public
	---Purpose: Add a point in the current polyline of the set 
	--	    or creates a new one when <NewPolyline> flag is TRUE.
	---Category: Update method

	Add(me : mutable; X1, Y1, X2, Y2: Length from Quantity);
	---Level: Public
	---Purpose: Add a segment in the set to one of polyline
	--	    which has the last point identical to one of the segment
	--	    or creates a new polyline in the sets with the 2 segment points.
	--	    The first point is <X1>, <Y1>.
	--	    The second point is <X2>, <Y2>.
	---Category: Update method

	Length(me) returns Integer from Standard;
	---Level: Public
	---Purpose: Returns the number of polylines in the set.
	---Category: Inquiry method

	Length(me; aPrank: Integer from Standard) 
		returns Integer from Standard
	---Level: Public
	---Purpose: Returns the number of points of the polylines
	--    of rank <aPrank>.
	--  Trigger: Raises OutOfRange if <aPrank> is <1 or >Length()
	raises OutOfRange from Standard;
	---Category: Inquiry method

	Values( me; aPrank : Integer from Standard;
	            aVrank : Integer from Standard;
		        X,Y    : out Length from Quantity)
	---Level: Public
	---Purpose: Returns the point of rank <aVrank>
	--	    from the polyline of rank <aPrank>.
	--  Trigger: Raises OutOfRange if <aPrank> is <1 or >Length()
	--	 or if <aVrank> is <1 or >Length(<aPrank>)
	raises OutOfRange from Standard;
	---Category: Inquiry method

	--------------------------
	-- Category: Draw and Pick
	--------------------------

	Draw (me : mutable; aDrawer: Drawer from Graphic2d)
	is static protected;
	---Level: Internal
	---Purpose: Draws the set of polylines <me>.

	Pick (me : mutable; X, Y: ShortReal from Standard;
		aPrecision: ShortReal from Standard;
		aDrawer: Drawer from Graphic2d)
	returns Boolean from Standard
	is static protected;
	---Level: Internal
        ---Purpose: Returns Standard_True if one point of the set <me> 
	--	    is picked, Standard_False if not.
	--  Warning: The PickIndex() method returns the rank of the picked
	--	    polyline point if any under the format :
	--	    (<aPrank> << 16) | <aVrank>.

	----------------------------------------------------------------------

	Save( me; aFStream: in out FStream from Aspect ) is virtual;
--	Retrieve( me; aIFStream: in out IFStream from AIS2D ) is virtual;

fields
	myPolylines:	SequenceOfPolyline from Graphic2d;

end SetOfPolylines from Graphic2d;
