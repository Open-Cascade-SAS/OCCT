-- Created on: 1992-08-21
-- Created by: Christophe MARION
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Intersection from HLRAlgo

	---Purpose: Describes  an intersection  on   an edge to  hide.
	--          Contains a parameter and   a state (ON =   on  the
	--          face, OUT = above the face, IN = under the Face)

uses
    Integer     from Standard,
    Real        from Standard,
    ShortReal   from Standard,
    Orientation from TopAbs,
    State       from TopAbs

is
    Create returns Intersection from HLRAlgo;

    Create(Ori    : Orientation from TopAbs;
           Lev    : Integer     from Standard;
           SegInd : Integer     from Standard;
           Ind    : Integer     from Standard;
           P      : Real        from Standard;
           Tol    : ShortReal   from Standard;
           S      : State       from TopAbs)
    returns Intersection from HLRAlgo;
    
    Orientation(me : in out; Ori : Orientation from TopAbs)
	---C++: inline
    is static;

    Orientation(me) returns Orientation from TopAbs
	---C++: inline
    is static;
    
    Level(me : in out; Lev : Integer from Standard)
	---C++: inline
    is static;

    Level(me) returns Integer from Standard
	---C++: inline
    is static;
    
    SegIndex(me : in out; SegInd : Integer from Standard)
	---C++: inline
    is static;

    SegIndex(me) returns Integer from Standard
	---C++: inline
    is static;
    
    Index(me : in out; Ind : Integer from Standard)
	---C++: inline
    is static;

    Index(me) returns Integer from Standard
	---C++: inline
    is static;
    
    Parameter(me : in out; P : Real from Standard)
	---C++: inline
    is static;

    Parameter(me) returns Real from Standard
	---C++: inline
    is static;
    
    Tolerance(me : in out; T : ShortReal from Standard)
	---C++: inline
    is static;
    
    Tolerance(me) returns ShortReal from Standard
	---C++: inline
    is static;
    
    State(me : in out; S : State from TopAbs)
	---C++: inline
    is static;

    State(me) returns State from TopAbs
	---C++: inline
    is static;

fields
    myOrien    : Orientation from TopAbs;
    mySegIndex : Integer     from Standard;
    myIndex    : Integer     from Standard;
    myLevel    : Integer     from Standard;
    myParam    : Real        from Standard;
    myToler    : ShortReal   from Standard;
    myState    : State       from TopAbs;

end Intersection;
