-- Created on: 1994-06-03
-- Created by: Christian CAILLET
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Activator  from IGESSelect  inherits Activator  from IFSelect

    ---Purpose : Performs Actions specific to IGESSelect, i.e. creation of
    --           IGES Selections and Dispatches, plus dumping specific to IGES

uses CString, SessionPilot, ReturnStatus

is

    Create returns mutable Activator from IGESSelect;


    Do   (me : mutable; number : Integer; pilot : mutable SessionPilot)
    	returns ReturnStatus;
    ---Purpose : Executes a Command Line for IGESSelect

    Help (me; number : Integer) returns CString;
    ---Purpose : Sends a short help message for IGESSelect commands

end Activator;
