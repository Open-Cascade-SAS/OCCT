-- Created on: 1993-01-20
-- Created by: Laurent PAINNOT
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.





class MyLineTool from AppDef

uses MultiLine     from AppDef,
     Pnt           from gp,
     Pnt2d         from gp,
     Vec           from gp,
     Vec2d         from gp,
     Array1OfPnt   from TColgp,
     Array1OfPnt2d from TColgp,
     Array1OfVec   from TColgp,
     Array1OfVec2d from TColgp,
     Status        from Approx

is
    
    
    FirstPoint(myclass; ML: MultiLine) returns Integer;
    	---Purpose: Returns the first index of multipoints of the MultiLine.


    LastPoint(myclass; ML: MultiLine) returns Integer;
    	---Purpose: Returns the last index of multipoints of the MultiLine.



    NbP2d(myclass; ML: MultiLine) returns Integer;
    	---Purpose: Returns the number of 2d points of a MultiLine.


    NbP3d(myclass; ML: MultiLine) returns Integer;
    	---Purpose: Returns the number of 3d points of a MultiLine.


    Value(myclass; ML: MultiLine; MPointIndex: Integer; 
          tabPt: out Array1OfPnt);
    	---Purpose: returns the 3d points of the multipoint <MPointIndex>
    	--          when only 3d points exist.


    Value(myclass; ML: MultiLine; MPointIndex: Integer; 
          tabPt2d: out Array1OfPnt2d);
    	---Purpose: returns the 2d points of the multipoint <MPointIndex>
    	--          when only 2d points exist.


    Value(myclass; ML: MultiLine; MPointIndex: Integer; 
          tabPt: out Array1OfPnt; tabPt2d: out Array1OfPnt2d);
    	---Purpose: returns the 3d and 2d points of the multipoint 
    	--          <MPointIndex>.


    Tangency(myclass; ML: MultiLine; MPointIndex: Integer; 
             tabV: out Array1OfVec) returns Boolean;
    	---Purpose: returns the 3d points of the multipoint <MPointIndex>
    	--          when only 3d points exist.


    Tangency(myclass; ML: MultiLine; MPointIndex: Integer; 
          tabV2d: out Array1OfVec2d) returns Boolean;
    	---Purpose: returns the 2d tangency points of the multipoint 
    	--          <MPointIndex> only when 2d points exist.


    Tangency(myclass; ML: MultiLine; MPointIndex: Integer; 
             tabV: out Array1OfVec; tabV2d: out Array1OfVec2d)
    returns Boolean;
    	---Purpose: returns the 3d and 2d points of the multipoint 
    	--          <MPointIndex>.


    Curvature(myclass; ML: MultiLine; MPointIndex: Integer; 
             tabV: out Array1OfVec) returns Boolean;
    	---Purpose: returns the 3d curvatures of the multipoint <MPointIndex>
    	--          when only 3d points exist.


    Curvature(myclass; ML: MultiLine; MPointIndex: Integer; 
          tabV2d: out Array1OfVec2d) returns Boolean;
    	---Purpose: returns the 2d curvatures of the multipoint 
    	--          <MPointIndex> only when 2d points exist.


    Curvature(myclass; ML: MultiLine; MPointIndex: Integer; 
             tabV: out Array1OfVec; tabV2d: out Array1OfVec2d)
    returns Boolean;
    	---Purpose: returns the 3d and 2d curvatures of the multipoint 
    	--          <MPointIndex>.



    WhatStatus(myclass; ML: MultiLine; I1, I2: Integer) 
    returns Status from Approx;
    	---Purpose:  returns NoPointsAdded
    
    MakeMLBetween(myclass; ML: MultiLine; I1, I2: Integer;
                  NbPMin: Integer) 
    returns MultiLine;
    	---Purpose: Is never called in the algorithms.
    	--          Nothing is done.
    	---C++: return &


end MyLineTool;
