-- Created on: 1992-09-22
-- Created by: Gilles DEBARBOUILLE
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


generic class Mat from MAT (Tool as any)

	---Purpose: this class contains the generic algoritm of 
	--          computation of the bisecting locus.

uses
    Side                     from MAT,
    Bisector                 from MAT,
    ListOfEdge              from MAT,
    ListOfBisector          from MAT,
    DataMapOfIntegerBisector from MAT,
    DataMapOfIntegerInteger  from TColStd
    
is

    Create
    ---Purpose: Empty construtor.
    returns Mat from MAT;
    
--- Category : Computation.    
    
    CreateMat(me : in out ; aTool : in out Tool)
       ---Purpose: Algoritm of computation of the bisecting locus.
    is static;
    
    IsDone(me) returns Boolean from Standard
       ---Purpose:  Returns <TRUE> if CreateMat has succeeded. 
    is static;

    LoadBisectorsToRemove(me                    : in out ; 
    	    	    	  noofbisectorstoremove : in out Integer;
    	    	          distance1             :        Real;
			  distance2             :        Real;
			  bisector1             :        Bisector from MAT;
			  bisector2             :        Bisector from MAT;
			  bisector3             :        Bisector from MAT;
			  bisector4             :        Bisector from MAT)
    is static private;


    Intersect( me                   : in out                   ;
    	       atool                : in out  Tool             ;
    	       aside                :         Integer          ;
    	       noofbisectorstoremove: in out  Integer           ;
	       bisector1            : mutable Bisector from MAT;
	       bisector2            : mutable Bisector from MAT)
    is static private;	       
  			       

--- Category : Querying.    
    
    Init(me : in out)
	--- Purpose : Initialize an iterator on the set of the roots
	--            of the trees of bisectors.
    is static;
    
    More(me) returns Boolean
	--- Purpose : Return False if there is no more roots.
    is static;
    
    Next(me : in out)
	--- Purpose : Move to the next root.
    is static;
    
    Bisector(me) returns any Bisector from MAT
	--- Purpose : Returns the current root.
    is static;

    SemiInfinite(me) returns Boolean from Standard
	--- Purpose : Returns True if there are semi_infinite bisectors.
	--            So there is a tree for each semi_infinte bisector.
    is static;

    NumberOfBisectors(me) returns Integer from Standard
	--- Purpose : Returns the total number of bisectors.
    is static;

fields

    thenumberofbisectors  : Integer;
    thenumberofedges      : Integer;
    semiInfinite          : Boolean;
    theedgelist           : ListOfEdge               from MAT;
    typeofbisectortoremove: DataMapOfIntegerInteger  from TColStd;
    bisectoronetoremove   : DataMapOfIntegerBisector from MAT;
    bisectortwotoremove   : DataMapOfIntegerBisector from MAT;
    bisectormap           : DataMapOfIntegerBisector from MAT;
    roots                 : ListOfBisector           from MAT;
    thecurrentindex       : Integer;
    isDone                : Boolean;             
    
end Mat;
