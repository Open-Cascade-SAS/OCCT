-- Created on: 1994-08-31
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class FaceInfo from Draft

	---Purpose: 

uses Surface  from Geom,
     Curve    from Geom,
     Face     from TopoDS


raises DomainError from Standard

is

    Create
    
    	returns FaceInfo from Draft;


    Create(S: Surface from Geom; HasNewGeometry: Boolean from Standard)
    
    	returns FaceInfo from Draft;


    RootFace(me: in out; F: Face from TopoDS)
    
    	is static;


    NewGeometry(me)
    
    	returns Boolean from Standard
	is static;
	

    Add(me: in out; F: Face from TopoDS)
    
    	is static;

    FirstFace(me)
    
    	returns Face from TopoDS
	---C++: return const&
	is static;


    SecondFace(me)
    
    	returns Face from TopoDS
	---C++: return const&
	is static;


    Geometry(me)
    
    	returns Surface from Geom
	is static;
	---C++: return const&

    ChangeGeometry(me: in out)
    
    	returns Surface from Geom
	is static;
	---C++: return &

    RootFace(me)
    
	---C++: return const&
    	returns Face from TopoDS
	is static;

    ChangeCurve(me: in out)
    
    	returns Curve from Geom
	---C++: return &
	is static;

    Curve(me)
    
    	returns Curve from Geom
	---C++: return const&
	is static;




fields

    myNewGeom : Boolean from Standard;
    myGeom    : Surface from Geom;
    myRootFace: Face    from TopoDS;
    myF1      : Face    from TopoDS;
    myF2      : Face    from TopoDS;
    myCurv    : Curve   from Geom;

end FaceInfo;
