-- Created on: 1992-03-06
-- Created by: Isabelle GRIGNON
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



generic class Iterator from IntWalk (Point as any)
                       

	---Purpose: Template class to describe the exploration argument of the
	--          generic class IWalking 


raises OutOfRange from Standard

is

    Create
    
    	returns Iterator from IntWalk;


    Length(me)
    
    	---Purpose: returns the dimension of the exploration

    	returns Integer from Standard

    	is static;


    Value(me; Index : Integer)
    
    	---Purpose: returns the current point
    	--          an exception is raised if i>NbPoints

    	returns  Point

    	raises OutOfRange from Standard

    	is static;


    Append(me: in out; P: Point)
    
	---Purpose: Adds a point in the iterator.
    
    	is static;
	
	
end Iterator;
