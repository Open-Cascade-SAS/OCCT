-- Created on: 2004-06-11
-- Created by: Alexander SOLOVYOV
-- Copyright (c) 2004-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DrawableMesh from XSDRAWSTLVRML inherits Drawable3D from Draw

	---Purpose:
uses
  Display from Draw,
  Mesh    from MeshVS

is
    Create ( aMesh : Mesh from MeshVS ) returns DrawableMesh from XSDRAWSTLVRML;
    DrawOn(me; dis : in out Display) is redefined virtual;

    GetMesh( me ) returns Mesh;

fields
    myMesh : Mesh;

end DrawableMesh;
