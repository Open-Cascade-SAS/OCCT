-- File:	TDataStd_HDataMapOfStringHArray1OfReal.cdl
-- Created:	Fri Aug 17 17:24:55 2007
-- Author:	Sergey ZARITCHNY
--		<szy@popox.nnov.matra-dtv.fr>
---Copyright:	Open CasCade SA 2007


class HDataMapOfStringHArray1OfReal from TDataStd inherits TShared from MMgt

	---Purpose: Extension of TDataStd_DataMapOfStringHArray1OfReal class  
    	--          to be manipulated by handle.

uses
    DataMapOfStringHArray1OfReal from TDataStd 
    
is
    Create( NbBuckets: Integer from Standard = 1 )  
    returns mutable HDataMapOfStringHArray1OfReal from TDataStd;    
     
    Create( theOther:  DataMapOfStringHArray1OfReal from TDataStd)  
    returns mutable HDataMapOfStringHArray1OfReal from TDataStd;
     
    Map( me ) returns DataMapOfStringHArray1OfReal from TDataStd
	---C++: return const &
        ---C++: inline      
    is static;	    	
	  
    ChangeMap( me: mutable ) returns DataMapOfStringHArray1OfReal from TDataStd 
    	---C++: return &
        ---C++: inline 
    is static; 	    	
 
fields
    
    myMap : DataMapOfStringHArray1OfReal from TDataStd ;  

end HDataMapOfStringHArray1OfReal;
