
-- File:	Graphic2d_CircleMarker.cdl
-- Created:	Tue Jun 22 16:36:51 1993
-- Author:	Jean Louis FRENKEL
--		<jlf@stylox>
-- Modified: TCL G002A, 28-11-00, new section "inquire methods"

---Copyright:	 Matra Datavision 1993

class CircleMarker from Graphic2d inherits VectorialMarker from Graphic2d

	---Purpose: The primitive CircleMarker
	--	    Every marker takes a reference point as an argument in
	--	    its constructor. CircleMarker and EllipsMarker take
	--	    another point as the center and PolylineMarker takes the
	--	    first point of its list as its origin.
	--	    The coordinates of the centre or origin point are offsets
	--	    with respect to the reference point.

	---Keywords: Primitive, CircleMarker
	---Warning:
	---References:

uses
	Drawer		from Graphic2d,
	GraphicObject	from Graphic2d,
	Length		from Quantity,
	PlaneAngle	from Quantity,
	FStream		from Aspect,
	IFStream	from Aspect


raises
	CircleDefinitionError	from Graphic2d

is
	-------------------------
	-- Category: Constructors
	-------------------------

	Create( aGraphicObject: GraphicObject from Graphic2d;
		    aXPosition, aYPosition: Length from Quantity;
		    X, Y: Length from Quantity;
		    Radius: Length from Quantity)
	returns mutable CircleMarker from Graphic2d
	---Level: Public
	---Purpose: Creates a complete circle.
	--	    The reference point is <aXPosition>, <aYPosition>
	--          The center is <X>, <Y>.
	--          The radius is <Radius>.
	--  Warning: Raises CircleDefinitionError if the
	--          radius is null.
	raises CircleDefinitionError from Graphic2d;

	Create( aGraphicObject: GraphicObject from Graphic2d;
		    aXPosition, aYPosition: Length from Quantity;
		    X, Y: Length from Quantity;
		    Radius: Length from Quantity;
		    Alpha , Beta: PlaneAngle from Quantity)
	returns mutable CircleMarker from Graphic2d
	---Level: Public
	---Purpose: Creates an arc.
	--	    The reference point is <aXPosition>, <aYPosition>
	--	    The center is <X>, <Y>.
	--	    The radius is <Radius>.
	--	    Angles are measured counterclockwise with 0 radian
	--	    at 3 o'clock.
	--  Warning: Raises CircleDefinitionError if the
	--          radius is null.
	raises CircleDefinitionError from Graphic2d;


	--------------------------
	-- Category: Draw and Pick
	--------------------------

	Draw (me : mutable; aDrawer: Drawer from Graphic2d)
	is static protected;
	---Level: Internal
	---Purpose: Draws the circle <me>.

	DrawElement( me : mutable; aDrawer: Drawer from Graphic2d;
                 anIndex: Integer from Standard)
        is redefined protected;
    ---Level: Internal
    ---Purpose: Draws element <anIndex> of the circle marker <me>.

    DrawVertex( me : mutable; aDrawer: Drawer from Graphic2d;
                anIndex: Integer from Standard)
        is redefined protected;
    ---Level: Internal
    ---Purpose: Draws vertex <anIndex> of the circle marker <me>.


	Pick (me : mutable; X, Y: ShortReal from Standard;
		aPrecision: ShortReal from Standard;
		aDrawer: Drawer from Graphic2d)
	returns Boolean from Standard is static protected;
	---Level: Internal
	---Purpose: Returns Standard_True if the circle <me> is picked,
	--	    Standard_False if not.

 	--------------------------------------
	-- Category: Inquire methods
	--------------------------------------

    Center( me; X, Y: out Length from Quantity );  
	---Level: Public
	---Purpose: returns the coordinates of center of the circle marker
	
	Radius( me ) returns Length from Quantity;
	---Level: Public
	---Purpose: returns the radius of this circle marker
	
	FirstAngle( me ) returns PlaneAngle from Quantity;
	---Level: Public
	---Purpose: returns the first angle of the arc marker
	
	SecondAngle( me ) returns PlaneAngle from Quantity;
	---Level: Public
	---Purpose: returns the second angle of the arc marker

	----------------------------------------------------------------------

	Save( me; aFStream: in out FStream from Aspect ) is virtual;
	Retrieve( myclass; anIFStream: in out IFStream from Aspect;
		aGraphicObject: GraphicObject from Graphic2d );

fields

	myX           : ShortReal from Standard;
	myY           :	ShortReal from Standard;
	myRadius      :	ShortReal from Standard;
	myFirstAngle  :	ShortReal from Standard;
	mySecondAngle :	ShortReal from Standard;
	myisArc       : Boolean from Standard;
	
end CircleMarker from Graphic2d;
