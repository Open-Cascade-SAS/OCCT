-- Created on: 1994-12-16
-- Created by: Frederic MAUPAS
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class TranslateShell from StepToTopoDS
    inherits Root from StepToTopoDS
    
    ---Purpose:
    --         

uses
    
    Shape               from TopoDS,
    TranslateShellError from StepToTopoDS,
    Tool                from StepToTopoDS,
    ConnectedFaceSet    from StepShape,
    NMTool              from StepToTopoDS

raises NotDone from StdFail
     
is

    Create returns TranslateShell;
    
    Create (CFS    : ConnectedFaceSet from StepShape;
            T      : in out Tool      from StepToTopoDS;
            NMTool : in out NMTool    from StepToTopoDS)
    	returns TranslateShell;
	    
    Init (me     : in out;
          CFS    : ConnectedFaceSet from StepShape;
          T      : in out Tool      from StepToTopoDS;
          NMTool : in out NMTool    from StepToTopoDS);

    Value (me) returns Shape from TopoDS
    	raises NotDone
	is static;
	---C++: return const &

    Error (me) returns TranslateShellError from StepToTopoDS;
    
fields

    myError  : TranslateShellError from StepToTopoDS;
    
    myResult : Shape               from TopoDS;

end TranslateShell;
