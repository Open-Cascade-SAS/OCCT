-- Created by: Peter KURNEV
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class AlgoTools3D from BOPTools
  ---Purpose:  
  --  The class contains handy static functions 
  --  dealing with the topology  
  --  This is the copy of BOPTools_AlgoTools3D.cdl file

uses  
    Pln   from gp, 
    Dir   from gp, 
    Pnt   from gp,   
    Pnt2d from gp,  
    
    Surface from Geom,
    
    Shape from TopoDS, 
    Wire  from TopoDS, 
    Face  from TopoDS,  
    Edge  from TopoDS,
    Solid from TopoDS,
     
    ShapeEnum   from TopAbs,     
    Orientation from TopAbs, 
    State       from TopAbs, 

    ListOfShape from BOPCol,  
     
    Context     from BOPInt,

    IndexedDataMapOfShapeListOfShape from BOPCol

is  

    DoSplitSEAMOnFace (myclass;  
              aSp:  Edge from TopoDS;              
              aF :  Face from TopoDS);
          ---Purpose:  
          -- Make the edge <aSp> seam edge for the face <aF>                            
          --
        
    GetNormalToFaceOnEdge (myclass;  
              aE:  Edge from TopoDS;              
              aF:  Face from TopoDS;   
              aT:  Real from Standard; 
              aD:out Dir from gp); 
          ---Purpose:  
          --- Computes normal to the face <aF> for the point on the edge <aE>  
          --- at parameter <aT>           
          ---
    GetNormalToFaceOnEdge (myclass;  
              aE:  Edge from TopoDS;              
              aF:  Face from TopoDS;   
              aD:out Dir from gp);          
          ---Purpose:  
          --- Computes normal to the face <aF> for the point on the edge <aE>  
          --- at arbitrary intermediate parameter 
          ---
 
    SenseFlag    (myclass;  
             aNF1   :  Dir from gp;
             aNF2   :  Dir from gp) 
          returns Integer from Standard;   
          ---Purpose: 
          --- Returns 1  if scalar product aNF1* aNF2>0.   
          --- Returns 0  if directions aNF1 aNF2 coinside  
          --- Returns -1 if scalar product aNF1* aNF2<0.      
          ---
    GetNormalToSurface    (myclass;  
              aS:  Surface from Geom; 
              U :  Real from Standard;
              V :  Real from Standard; 
              aD:out Dir from gp)
          returns Boolean from Standard;   
          ---Purpose:  
          --- Compute normal <aD> to surface <aS> in point (U,V)  
          --- Returns TRUE if directions aD1U, aD1V coinside 
          ---
 
    GetApproxNormalToFaceOnEdge (myclass;  
              aE:  Edge from TopoDS;              
              aF:  Face from TopoDS;   
              aT:  Real from Standard;  
              aPx:out Pnt from gp;
              aD:out Dir from gp; 
              theContext:out Context from BOPInt); 
          ---Purpose:  
          --- Computes normal to the face <aF> for the 3D-point that 
          --- belonds to the edge <aE> at parameter <aT>. 
          --  Output: 
          --- aPx  -  the 3D-point where the normal computed 
          --- aD   -  the normal; 
          ---
          --  Warning:
          --- The normal is computed not exactly in the point on the 
          --- edge, but in point that is near to the edge towards to 
          --- the face material (so, we'll have approx. normal) 
          --- 
           
    GetApproxNormalToFaceOnEdge(myclass; 
              theE : Edge from TopoDS; 
              theF : Face from TopoDS; 
              aT   : Real from Standard; 
              aP   : out Pnt  from gp; 
              aDNF : out Dir  from gp; 
              aDt2D: Real from Standard);
          
    PointNearEdge   (myclass;   
              aE   :  Edge from TopoDS;              
              aF   :  Face from TopoDS;   
              aT   :  Real from Standard;  
              aDt2D:  Real from Standard;  
              aP2D :out Pnt2d from  gp; 
              aPx  :out Pnt from gp);
          ---Purpose: 
          --- Compute the point <aPx>,  (<aP2D>)  that is near to  
          --- the edge <aE>   at parameter <aT>  towards to the  
          --- material of the face <aF>. The value of shifting in 
          --- 2D is <aDt2D> 
          ---
    PointNearEdge   (myclass;   
              aE:  Edge from TopoDS;              
              aF:  Face from TopoDS;   
              aT:  Real from Standard;  
              aP2D:out Pnt2d from  gp; 
              aPx:out Pnt from gp; 
              theContext:out Context from BOPInt);
          ---Purpose: 
          --- Computes the point <aPx>,  (<aP2D>)  that is near to  
          --- the edge <aE>   at parameter <aT>  towards to the  
          --- material of the face <aF>. The value of shifting in 
          --  2D is  dt2D=BOPTools_AlgoTools3D::MinStepIn2d()
          ---
    PointNearEdge   (myclass;   
              aE:  Edge from TopoDS;              
              aF:  Face from TopoDS;   
              aP2D:out Pnt2d from  gp; 
              aPx:out Pnt from gp; 
              theContext:out Context from BOPInt);
          ---Purpose: 
          --- Compute the point <aPx>,  (<aP2D>)  that is near to  
          --- the edge <aE>   at arbitrary  parameter  towards to the  
          --- material of the face <aF>. The value of shifting in 
          --  2D is  dt2D=BOPTools_AlgoTools3D::MinStepIn2d()
          ---
 
    MinStepIn2d(myclass) 
          returns  Real from Standard;  
          ---Purpose:  
          --- Returns simple step value that is used in 2D-computations 
          --- = 1.e-5 
          ---
    IsEmptyShape(myclass; 
              aS:  Shape from TopoDS) 
          returns Boolean from Standard; 
          ---Purpose: 
          --- Returns TRUE if the shape <aS> does not contain 
          --- geometry information  (e.g. empty compound) 
          ---
 
    OrientEdgeOnFace  (myclass;  
              aE    :  Edge from TopoDS;
              aF    :  Face from TopoDS;  
              aER   : out  Edge from TopoDS); 
          ---Purpose:  
          --- Get the edge <aER> from the face <aF> that is the same as   
          --- the edge <aE>    
          --- 

    PointInFace(myclass;
              theF:Face from TopoDS;
              theP:out Pnt from gp;
              theP2D:out Pnt2d from gp; 
              theContext:out Context from BOPInt) 
          returns Integer from Standard; 
          ---Purpose: Computes a point <theP> inside the face <theF>. <br>
          --          <theP2D> -  2D  representation of <theP> <br>
          --          on the surface of <theF> <br>
          --          Returns 0 in case of success. <br>

end AlgoTools3D;
