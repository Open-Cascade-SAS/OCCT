-- Created on: 1991-04-03
-- Created by: Remi GILET
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class LinPnt2dBisec

from GccAna

	---Purpose: Describes functions for building bisecting curves between a 2D line and a point.
    	-- A bisecting curve between a line and a point is such a
    	-- curve that each of its points is at the same distance from
    	-- the circle and the point. It can be a parabola or a line,
    	-- depending on the relative position of the line and the
    	-- circle. There is always one unique solution.
    	-- A LinPnt2dBisec object provides a framework for:
    	-- - defining the construction of the bisecting curve,
    	-- - implementing the construction algorithm, and
    	-- - consulting the result.

--inherits Storable from Standard

uses Lin2d from gp,
     Pnt2d from gp,
     Bisec from GccInt

raises ConstructionError from Standard,
       NotDone           from StdFail

is

Create(Line1   : Lin2d from gp;
       Point2  : Pnt2d from gp) returns LinPnt2dBisec
raises ConstructionError;
    	---Purpose: Constructs a bisecting curve between the line Line1 and the point Point2.

IsDone(me) returns Boolean from Standard
is static;
    	---Purpose : Returns True if the algorithm succeeded.

ThisSolution(me) returns Bisec from GccInt
    	---Purpose : Returns the number of solutions.
raises NotDone
is static;
    	---Purpose: It raises NotDone if the construction algorithm didn't succeed.

fields

    WellDone : Boolean from Standard;
    	---Purpose:  True if the algorithm succeeded.

    bissol   : Bisec from GccInt;
    	---Purpose : The solutions.

end LinPnt2dBisec;
