-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class OrganizationAssignment from StepBasic 

inherits TShared from MMgt

uses

	Organization from StepBasic, 
	OrganizationRole from StepBasic
is

	Init (me : mutable;
	      aAssignedOrganization : mutable Organization from StepBasic;
	      aRole : mutable OrganizationRole from StepBasic) is virtual;

	-- Specific Methods for Field Data Access --

	SetAssignedOrganization(me : mutable; aAssignedOrganization : mutable Organization);
	AssignedOrganization (me) returns mutable Organization;
	SetRole(me : mutable; aRole : mutable OrganizationRole);
	Role (me) returns mutable OrganizationRole;

fields

	assignedOrganization : Organization from StepBasic;
	role : OrganizationRole from StepBasic;

end OrganizationAssignment;
