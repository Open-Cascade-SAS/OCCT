-- Created on: 1995-10-24
-- Created by: Mister rmi
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Triangulation from PPoly inherits Persistent from Standard

	---Purpose: This class represents a 3d polyhedral triangulation.
	--          
	--          It is defined by :
	--          
	--          * A Deflection : This  is the distance between the
	--          triangulation and the "ideal" surface.
	--          
	--          *  An  Array1 of 3d   nodes  values : Contains the
	--          Points for the 3d  nodes. Two different  nodes may
	--          have the same  3d point if  they are differents in
	--          UV space.
	--          
	--          * An  Array1 of 2d nodes  values : Contains the UV
	--          coordinates  for   the   nodes   in the    surface
	--          parametric  space. This is optionnal.
	--          
	--          * The  Array of  triangles,   each triangle  is  a
	--          triplet of  node indices.  A  triangle is oriented
	--          and the  whole triangulation  must have a coherent
	--          orientation.

uses
   HArray1OfPnt2d    from PColgp,
   HArray1OfPnt      from PColgp,
   HArray1OfTriangle from PPoly

is

    Create(Defl:       Real              from Standard;
    	   Nodes:      HArray1OfPnt      from PColgp;
    	   Triangles:  HArray1OfTriangle from PPoly)
    returns mutable Triangulation from PPoly;
    	---Purpose: Defaults with allocation of Nodes and Triangles.

    Create(Defl:       Real              from Standard;
    	   Nodes:      HArray1OfPnt      from PColgp;
    	   UVNodes:    HArray1OfPnt2d    from PColgp;
    	   Triangles:  HArray1OfTriangle from PPoly)
    returns mutable Triangulation from PPoly;
    	---Purpose: Defaults with allocation of Nodes and Triangles.

    Deflection(me) returns Real;
    
    Deflection(me : mutable; D : Real);

    NbNodes(me) returns Integer;
	---Purpose: Null if the nodes are not yet defined.

    NbTriangles(me) returns Integer;
	---Purpose: Null if the Triangles are not yet defined.

    HasUVNodes(me) returns Boolean;

    Nodes(me) returns HArray1OfPnt from PColgp;
	---Purpose: Const reference on the 3d nodes values.
    	
    UVNodes(me) returns HArray1OfPnt2d from PColgp;
	---Purpose: Const reference on the 2d nodes values.

    Triangles(me) returns HArray1OfTriangle from PPoly;
	---Purpose: Const reference on the triangles.

fields

    myDeflection  : Real;
    myNodes       : HArray1OfPnt      from PColgp;
    myUVNodes     : HArray1OfPnt2d    from PColgp;
    myTriangles   : HArray1OfTriangle from PPoly;

end Triangulation;
