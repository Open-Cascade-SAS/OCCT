-- Created on: 1993-07-13
-- Created by: Jean Louis FRENKEL
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class ViewMapping from Graphic2d inherits TShared from MMgt

	---Version:

	---Purpose: A ViewMapping defines a square region of the model
	--	    space from an origin point and a size in meters.
	--	    This square region is called the "map from".

	---Keywords:
	---Warning:
	---References:

uses
	Length from Quantity,
	Factor from Quantity

is
	-------------------------
	-- Category: Constructors
	-------------------------

	Create
	returns mutable ViewMapping from Graphic2d;
	---Level: Public
	---Purpose: Creates a view mapping with the following default
	--	    values :
	--		XCenter	= 0.
	--		YCenter	= 0.
	--		Size	= 1.
	---Category: Constructors

	---------------------------------------------------
	-- Category: Methods to modify the class definition
	---------------------------------------------------

	SetViewMapping (me: mutable;
		aXCenter, aYCenter: Length from Quantity;
		aSize: Length from Quantity)
	is static;
	---Level: Public
	---Purpose: Sets new values for the view mapping <me>.
	---Category: Methods to modify the class definition

	SetCenter (me: mutable;
		aXCenter, aYCenter: Length from Quantity)
	is static;
	---Level: Public
	---Purpose: Sets new values for the view mapping center.
	---Category: Methods to modify the class definition

	SetSize (me: mutable;
		aSize: Length from Quantity)
	is static;
	---Level: Public
	---Purpose: Sets new value for the view mapping size.

	SetViewMappingDefault (me: mutable)
	is static;
	---Level: Public
	---Purpose: Saves the current mapping which will be the
	--	    reference value for the reset of the mapping
	--	    done by the ViewmappingReset method.
	---Category: Methods to modify the class definition

	ViewMappingReset (me: mutable)
	is static;
	---Level: Public
	---Purpose: Sets the value of the mapping to be the same as
	--	    the mapping saved by the SetViewMappingDefault method.
	---Category: Methods to modify the class definition

	----------------------------
	-- Category: Inquire methods
	----------------------------

	ViewMapping (me; XCenter, YCenter, Size: out Length from Quantity)
	is static;
	---Level: Public
	---Purpose: Returns the current mapping of the view <me>.
	---Category: Inquire methods

	Center (me; XCenter, YCenter: out Length from Quantity)
	is static;
	---Level: Public
	---Purpose: Returns the current center of the view <me>.
	---Category: Inquire methods

	ViewMappingDefault (me;
		XCenter, YCenter, Size: out Length from Quantity)
	is static;
	---Level: Public
	---Purpose: Returns the current reset mapping of the view <me>.
	---Category: Inquire methods

	Zoom (me)
	returns Factor from Quantity
	is static;
	---Level: Public
	---Purpose: Returns the zoom factor (CurrentSize/InitialSize).
	---Category: Inquire methods

fields
	myXCenter:	Length from Quantity;
	myYCenter:	Length from Quantity;
	mySize:		Length from Quantity;

	myInitialXCenter:	Length from Quantity;
	myInitialYCenter:	Length from Quantity;
	myInitialSize:		Length from Quantity;

end ViewMapping from Graphic2d;
