-- Created on: 1993-09-07
-- Created by: Christian CAILLET
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class SpecificModule  from IGESDimen  inherits  SpecificModule from IGESData

    ---Purpose : Defines Services attached to IGES Entities :
    --           Dump & OwnCorrect, for IGESDimen

uses Messenger from Message, IGESEntity, IGESDumper

is

    Create returns mutable SpecificModule from IGESDimen;
    ---Purpose : Creates a SpecificModule from IGESDimen & puts it into SpecificLib

    OwnDump (me; CN : Integer; ent : IGESEntity;
    	      dumper : IGESDumper;  S : Messenger from Message; own : Integer);
    ---Purpose : Specific Dump (own parameters) for IGESDimen

    OwnCorrect (me; CN : Integer; ent : mutable IGESEntity)
    	returns Boolean  is redefined;
    ---Purpose : Performs non-ambiguous Corrections on Entities which support
    --           them (BasicDimension,CenterLine,DimensionDisplayData,
    --           DimensionTolerance,DimensionUnits,DimensionedGeometry,
    --           NewDimensionedGeometry,Section,WitnessLine)

end SpecificModule;
