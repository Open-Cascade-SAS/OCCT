-- Created on: 1992-09-22
-- Created by: Gilles DEBARBOUILLE
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package MAT

uses
    MMgt,
    TCollection,
    TColStd

is

    generic class Tool;
  	--- Purpose: The template class used in Mat.
   
    generic class Mat;
        --- Purpose: The Algorithm of Computation of the Map of 
        --           bisecting locus.


    --------------------------------------------------
    --  Classes of exploration of the Bisecting Locus.
    --------------------------------------------------
    enumeration Side is Left,Right end Side;
    	--- Purpose: Definition on the Left and the Right on the Fig.

    class Graph;
	--- Purpose: Graph of exploration of the Bisecting Locus.

    class Arc;
    	--- Purpose: Arc of Graph. 
    
    class Node;
    	--- Purpose: Node of Graph.
  
    class BasicElt;
	--- Purpose: BasicElt of Graph.
    
    class Zone;
	--- Purpose: Class Zone contains the frontiere of the Zone of proximity
	--           of a BasicElt.

    class SequenceOfBasicElt instantiates Sequence from TCollection
                                                         (BasicElt from MAT); 
						     
    class SequenceOfArc instantiates Sequence from TCollection
                                                         (Arc from  MAT) ;  

    class DataMapOfIntegerArc instantiates
    	DataMap from TCollection(Integer          from Standard,
	    	    	    	 Arc              from MAT     ,
				 MapIntegerHasher from TColStd);

    class DataMapOfIntegerBasicElt instantiates
    	DataMap from TCollection(Integer          from Standard,
	    	    	    	 BasicElt         from MAT     ,
				 MapIntegerHasher from TColStd);
 
    class DataMapOfIntegerNode instantiates
    	DataMap from TCollection(Integer          from Standard,
	    	    	    	 Node             from MAT     ,
				 MapIntegerHasher from TColStd);
 
 
    --------------------------------------------------- 
    --  Classes used for the computation of the Mat.
    --------------------------------------------------- 

    generic class TList, TListNode;

    class Bisector;
	
    class DataMapOfIntegerBisector instantiates
    	DataMap from TCollection(Integer          from Standard,
	    	    	    	 Bisector         from MAT     ,
				 MapIntegerHasher from TColStd);
				 
    class ListOfBisector instantiates TList from MAT (Bisector from MAT);
    
    class Edge;
    
    class ListOfEdge instantiates TList from MAT (Edge from MAT);
    
end MAT;




