-- File:        Edge.cdl
-- Created:     Fri Dec  1 11:11:19 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class Edge from StepShape 

inherits TopologicalRepresentationItem from StepShape 

uses

	Vertex from StepShape, 
	HAsciiString from TCollection
is

	Create returns mutable Edge;
	---Purpose: Returns a Edge


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aEdgeStart : mutable Vertex from StepShape;
	      aEdgeEnd : mutable Vertex from StepShape) is virtual;

	-- Specific Methods for Field Data Access --

	SetEdgeStart(me : mutable; aEdgeStart : mutable Vertex)
    	is virtual;
	EdgeStart (me) returns mutable Vertex
    	is virtual;
	SetEdgeEnd(me : mutable; aEdgeEnd : mutable Vertex)
    	is virtual;
	EdgeEnd (me) returns mutable Vertex
    	is virtual;

fields

	edgeStart : Vertex from StepShape;
	edgeEnd : Vertex from StepShape;

end Edge;
