-- Created on: 1993-02-22
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class Surface from BRepAdaptor inherits Surface from Adaptor3d

	---Purpose: The Surface from BRepAdaptor allows to  use a Face
	--          of the BRep topology look like a 3D surface.
	--          
	--          It  has  the methods  of  the class   Surface from
	--          Adaptor3d.
	--          
	--          It is created or initialized with a Face. It takes
	--          into account the local coordinates system.
	--          
	--          The  u,v parameter range is   the minmax value for
	--          the  restriction,  unless  the flag restriction is
	--          set to false.

uses
    Face            from TopoDS,
    SurfaceType     from GeomAbs,
    HSurface        from Adaptor3d,
    HCurve          from Adaptor3d,
    Surface         from GeomAdaptor,
    Shape           from GeomAbs,
    BezierSurface   from Geom,
    BSplineSurface  from Geom,
    Trsf            from gp,
    Pnt             from gp,
    Vec             from gp,
    Dir             from gp,
    Pln             from gp,
    Cylinder        from gp,
    Sphere          from gp,
    Torus           from gp,
    Cone            from gp,
    Ax1             from gp,
    Array1OfReal    from TColStd


raises 

    OutOfRange   from Standard,
    DomainError  from Standard,
    NoSuchObject from Standard

is

    Create returns Surface from BRepAdaptor;
	---Purpose: Creates an undefined surface with no face loaded.
	
    Create(F : Face from TopoDS;
           R : Boolean = Standard_True) 
    returns Surface from BRepAdaptor;
	---Purpose: Creates a surface to  access the geometry  of <F>.
	--          If  <Restriction> is  true  the parameter range is
	--          the  parameter  range  in   the  UV space  of  the
	--          restriction. 
	
    Initialize(me : in out; F : Face from TopoDS; 
    	    	    	    Restriction : Boolean = Standard_True)
	---Purpose: Sets the surface to the geometry of <F>.
    is static;
    
    Surface(me) returns Surface from GeomAdaptor
	---Purpose: Returns the surface.
	--          
	---C++: return const &
    is static;
    
    ChangeSurface(me : in out) returns Surface from GeomAdaptor
	---Purpose: Returns the surface.
	--          
	---C++: return &
    is static;
    
    Trsf(me) returns Trsf from gp
	---Purpose: Returns the surface coordinate system.
	--          
	---C++: return const &
    is static;
    
    Face(me) returns Face from TopoDS
	---Purpose: Returns the face.
	--          
	---C++: return const &
    is static;
    
    Tolerance(me) returns Real
	---Purpose: Returns the face tolerance.
	--          
    is static;

    --
    --  Methods of Surface from GeomAdaptor
    --              
    
    FirstUParameter(me) returns Real
         ---C++:inline
    is redefined static;

    LastUParameter(me) returns Real
         ---C++:inline
    is redefined static;
    
    FirstVParameter(me) returns Real
         ---C++:inline
    is redefined static;

    LastVParameter(me) returns Real
         ---C++:inline
    is redefined static;
    
    UContinuity(me) returns Shape from GeomAbs
         ---C++:inline
    is redefined static;
    
    VContinuity(me) returns Shape from GeomAbs
         ---C++:inline
    is redefined static;
    
    NbUIntervals(me; S : Shape from GeomAbs) returns Integer
	---Purpose: If necessary, breaks the surface in U intervals of
	--          continuity    <S>.  And   returns  the  number  of
	--          intervals.
        ---C++:inline
    is redefined static;
    
    NbVIntervals(me; S : Shape from GeomAbs) returns Integer
	---Purpose: If necessary, breaks the surface in V intervals of
	--          continuity    <S>.  And   returns  the  number  of
	--          intervals.
        ---C++:inline
    is redefined static;
    
    UIntervals(me; T : in out Array1OfReal from TColStd; 
    	    	   S :        Shape        from GeomAbs ) 
	---Purpose: Returns the  intervals with the requested continuity
	--          in the U direction.
    raises
    	OutOfRange from Standard -- if the Length of the array does
	    	    	         -- have enought slots to accomodate
	    	    	         -- the result.
    is redefined static;

    VIntervals(me; T : in out Array1OfReal from TColStd; 
    	    	   S :        Shape        from GeomAbs ) 
	---Purpose: Returns the  intervals with the requested continuity
	--          in the V direction.
    raises
    	OutOfRange from Standard -- if the Length of the array does
	    	    	         -- have enought slots to accomodate
	    	    	         -- the result.
    is redefined static;
    
    UTrim(me; First, Last, Tol : Real) returns HSurface from Adaptor3d
	---Purpose: Returns    a  surface trimmed in the U direction
	--           equivalent   of  <me>  between
	--          parameters <First>  and <Last>. <Tol>  is used  to
	--          test for 3d points confusion.
    raises
    	OutOfRange from Standard
	---Purpose: If <First> >= <Last> 
    is redefined static ;
    
    VTrim(me; First, Last, Tol : Real) returns HSurface from Adaptor3d
	---Purpose: Returns    a  surface trimmed in the V direction  between
	--          parameters <First>  and <Last>. <Tol>  is used  to
	--          test for 3d points confusion.
    raises
    	OutOfRange from Standard
	---Purpose: If <First> >= <Last> 
    is redefined static ;

    IsUClosed(me) returns Boolean
         ---C++:inline
    is redefined static;
     
    IsVClosed(me) returns Boolean
         ---C++:inline
    is redefined static;
     
    IsUPeriodic(me) returns Boolean
         ---C++:inline
    is redefined static;
    
    UPeriod(me) returns Real
    raises
    	DomainError from Standard -- if the curve is not periodic
         ---C++:inline
    is redefined static;
     
    IsVPeriodic(me) returns Boolean
         ---C++:inline
    is redefined static;
    
    VPeriod(me) returns Real
         ---C++:inline
    raises
    	DomainError from Standard -- if the curve is not periodic
    is redefined static;
     
    Value (me; U, V : Real)  returns Pnt from gp
        --- Purpose : Computes the point of parameters U,V on the surface.
    is redefined static;

    D0 (me; U, V : Real; P : out Pnt from gp)
        --- Purpose : Computes the point of parameters U,V on the surface.
    is redefined static;

    D1 (me; U, V     : Real; 
    	    P        : out Pnt from gp; 
    	    D1U, D1V : out Vec from gp)
        --- Purpose : Computes the point  and the first derivatives on
        --  the surface.
    raises 
    	DomainError from Standard
            --- Purpose   : Raised   if  the continuity  of   the  current
            --  intervals is not C1.
    is redefined static;

    D2 (me; U, V : Real; 
    	    P : out Pnt from gp; 
    	    D1U, D1V, D2U, D2V, D2UV : out Vec from gp)
        --- Purpose  :  Computes   the point,  the  first  and  second
        --  derivatives on the surface.
    raises 
    	DomainError from Standard
            --- Purpose   : Raised  if   the   continuity   of the current
            --  intervals is not C2.
    is redefined static;

    D3 (me; U, V : Real; P : out Pnt from gp; 
    	    D1U, D1V, D2U, D2V, D2UV, D3U, D3V, D3UUV, D3UVV : out Vec from gp)
        --- Purpose : Computes the point,  the first, second and third
        --  derivatives on the surface.
    raises 
    	DomainError from Standard
            --- Purpose   : Raised  if   the   continuity   of the current
            --  intervals is not C3.
    is redefined static;

    DN (me; U, V : Real; Nu, Nv : Integer)   returns Vec from gp
        --- Purpose :  Computes the derivative of order Nu in the direction 
        --  U and Nv in the direction V at the point P(U, V).
    raises 
    	DomainError from Standard,
            --- Purpose : Raised if the current U  interval is not not CNu
            --  and the current V interval is not CNv.
        OutOfRange from Standard
            --- Purpose : Raised if Nu + Nv < 1 or Nu < 0 or Nv < 0.
    is redefined static;
  
    UResolution(me; R3d : Real ) returns Real
         ---Purpose :  Returns the parametric U  resolution corresponding
         --         to the real space resolution <R3d>.
         --         
	---C++:inline
    is redefined static;
  
    VResolution(me; R3d : Real ) returns Real
         ---Purpose :  Returns the parametric V  resolution corresponding
         --         to the real space resolution <R3d>.
         --         
	---C++:inline
    is redefined static;
  
    GetType(me) returns SurfaceType from GeomAbs
	---Purpose: Returns the type of the surface : Plane, Cylinder,
	--          Cone,      Sphere,        Torus,    BezierSurface,
	--          BSplineSurface,               SurfaceOfRevolution,
	--          SurfaceOfExtrusion, OtherSurface
	---C++:inline
    is redefined static;
    
    Plane(me) returns Pln from gp
      raises NoSuchObject from Standard
      
    is redefined static;
    
    Cylinder(me) returns Cylinder from gp
      raises NoSuchObject from Standard
    is redefined static;
    
    Cone(me) returns Cone from gp
      raises NoSuchObject from Standard
    is redefined static;
    
    Sphere(me) returns Sphere from gp
      raises NoSuchObject from Standard
    is redefined static;
    
    Torus(me) returns Torus from gp
      raises NoSuchObject from Standard
    is redefined static;


    UDegree(me) returns Integer 
     raises NoSuchObject from Standard
     ---C++:inline
    is redefined static;

    NbUPoles(me) returns Integer
     raises NoSuchObject from Standard
    ---C++:inline
    is redefined static;

    VDegree(me) returns Integer
     raises NoSuchObject from Standard
	---C++:inline    
    is redefined static;

    NbVPoles(me) returns Integer
     raises NoSuchObject from Standard
	---C++:inline     
    is redefined static;
    
    
    NbUKnots(me) returns Integer
    raises 
       NoSuchObject from Standard
	---C++:inline       
    is redefined static;
    
    
    NbVKnots(me) returns Integer
    raises 
       NoSuchObject from Standard
	---C++:inline       
    is redefined static;
    
    
    IsURational(me) returns Boolean
    raises
    	NoSuchObject from Standard
	---C++:inline	
    is redefined static;
    
    IsVRational(me) returns Boolean
    raises
    	NoSuchObject from Standard
	---C++:inline	
    is redefined static;
    

    Bezier(me) returns BezierSurface from Geom
    	---Purpose: 
--Warning : this will make a copy of the 
    	--           Bezier Surface since it applies
    	--           to it the myTsrf transformation
    	--           Be Carefull when using this method

    raises 
    	NoSuchObject from Standard
    is redefined static;

    BSpline(me) returns BSplineSurface from Geom
    	---Purpose: 
--  Warning : this will make a copy of the 
    	--           BSpline Surface since it applies
    	--           to it the myTsrf transformation
    	--           Be Carefull when using this method

    raises 
    	NoSuchObject from Standard
    is redefined static;
    
    AxeOfRevolution(me) returns Ax1 from gp
    raises 
       NoSuchObject from Standard -- only for SurfaceOfRevolution
    is redefined static;

    Direction(me) returns Dir from gp
    raises 
       NoSuchObject from Standard -- only for SurfaceOfExtrusion
    is redefined static;

    BasisCurve(me) returns HCurve from Adaptor3d
    raises 
       NoSuchObject from Standard
       ---Purpose: only for SurfaceOfExtrusion and SurfaceOfRevolution
       --  Warning: this will make a copy of the underlying curve
       --          since it applies to it the transformation
       --          myTrsf. Be carefull when using this method.
    is redefined static;

    BasisSurface(me) returns HSurface from Adaptor3d
    raises 
       NoSuchObject from Standard -- only for Offset Surface
    is redefined static;

    OffsetValue(me) returns Real from Standard
    raises 
       NoSuchObject from Standard -- only for Offset Surface
    is redefined static;

fields

    mySurf : Surface from GeomAdaptor;
    myTrsf : Trsf from gp;
    myFace : Face from TopoDS;

end Surface;
