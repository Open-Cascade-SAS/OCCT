-- Created on: 1997-02-12
-- Created by: Alexander BRIVIN
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MatrixTransform from Vrml 

	---Purpose: defines a MatrixTransform node of VRML specifying matrix and transform
	--          properties. 
    	--  This  node  defines  3D  transformation  with  a  4  by  4  matrix.
    	--  By  default  :   
    	--  a11=1  a12=0  a13=0  a14=0
    	--  a21=0  a22=1  a23=0  a24=0
    	--  a31=0  a32=0  a33=1  a34=0
    	--  a41=0  a42=0  a43=0  a44=1	
	--  It  is  written  to  the  file  in  row-major  order  as  16  Real numbers 
	--  separated  by  whitespace.  For  example ,  matrix  expressing  a  translation 
	--  of  7.3  units  along  the  X  axis  is  written  as: 
	--  1  0  0  0   0  1  0  0   0  0  1  0   7.3 0  0  1
uses
 
   Trsf   from   gp

is
 
    Create returns  MatrixTransform from Vrml;
 
    Create  ( aMatrix  :  Trsf    from  gp )
        returns  MatrixTransform from Vrml;
   
    SetMatrix ( me : in out;  aMatrix  :  Trsf    from  gp );
    Matrix ( me )  returns  Trsf    from  gp;

    Print  ( me;  anOStream: in out OStream from Standard) returns OStream from Standard;
    ---C++:  return  & 

fields
 
    myMatrix  :  Trsf    from  gp; -- Transformation matrix

end MatrixTransform;

