-- File:        BSplineSurfaceWithKnotsAndRationalBSplineSurface.cdl
-- Created:     Fri Dec  1 11:11:32 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class BSplineSurfaceWithKnotsAndRationalBSplineSurface from StepGeom 

inherits BSplineSurface from StepGeom 


	--- This classe is an implementation of EXPRESS
	--  ANDOR Subtype Declaration.
uses

	BSplineSurfaceWithKnots from StepGeom, 
	RationalBSplineSurface from StepGeom, 
	HAsciiString from TCollection, 
	Integer from Standard, 
	HArray2OfCartesianPoint from StepGeom, 
	BSplineSurfaceForm from StepGeom, 
	Logical from StepData, 
	HArray1OfInteger from TColStd, 
	HArray1OfReal from TColStd, 
	HArray2OfReal from TColStd, 
	KnotType from StepGeom
is

	Create returns mutable BSplineSurfaceWithKnotsAndRationalBSplineSurface;
	---Purpose: Returns a BSplineSurfaceWithKnotsAndRationalBSplineSurface


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aUDegree : Integer from Standard;
	      aVDegree : Integer from Standard;
	      aControlPointsList : mutable HArray2OfCartesianPoint from StepGeom;
	      aSurfaceForm : BSplineSurfaceForm from StepGeom;
	      aUClosed : Logical from StepData;
	      aVClosed : Logical from StepData;
	      aSelfIntersect : Logical from StepData) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aUDegree : Integer from Standard;
	      aVDegree : Integer from Standard;
	      aControlPointsList : mutable HArray2OfCartesianPoint from StepGeom;
	      aSurfaceForm : BSplineSurfaceForm from StepGeom;
	      aUClosed : Logical from StepData;
	      aVClosed : Logical from StepData;
	      aSelfIntersect : Logical from StepData;
	      aBSplineSurfaceWithKnots : mutable BSplineSurfaceWithKnots from StepGeom;
	      aRationalBSplineSurface : mutable RationalBSplineSurface from StepGeom) is virtual;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aUDegree : Integer from Standard;
	      aVDegree : Integer from Standard;
	      aControlPointsList : mutable HArray2OfCartesianPoint from StepGeom;
	      aSurfaceForm : BSplineSurfaceForm from StepGeom;
	      aUClosed : Logical from StepData;
	      aVClosed : Logical from StepData;
	      aSelfIntersect : Logical from StepData;
	      aUMultiplicities : mutable HArray1OfInteger from TColStd;
	      aVMultiplicities : mutable HArray1OfInteger from TColStd;
	      aUKnots : mutable HArray1OfReal from TColStd;
	      aVKnots : mutable HArray1OfReal from TColStd;
	      aKnotSpec : KnotType from StepGeom;
	      aWeightsData : mutable HArray2OfReal from TColStd) is virtual;

	-- Specific Methods for Field Data Access --

	SetBSplineSurfaceWithKnots(me : mutable; aBSplineSurfaceWithKnots : mutable BSplineSurfaceWithKnots);
	BSplineSurfaceWithKnots (me) returns mutable BSplineSurfaceWithKnots;
	SetRationalBSplineSurface(me : mutable; aRationalBSplineSurface : mutable RationalBSplineSurface);
	RationalBSplineSurface (me) returns mutable RationalBSplineSurface;

	-- Specific Methods for ANDOR Field Data Access --

	SetUMultiplicities(me : mutable; aUMultiplicities : mutable HArray1OfInteger);
	UMultiplicities (me) returns mutable HArray1OfInteger;
	UMultiplicitiesValue (me; num : Integer) returns Integer;
	NbUMultiplicities (me) returns Integer;
	SetVMultiplicities(me : mutable; aVMultiplicities : mutable HArray1OfInteger);
	VMultiplicities (me) returns mutable HArray1OfInteger;
	VMultiplicitiesValue (me; num : Integer) returns Integer;
	NbVMultiplicities (me) returns Integer;
	SetUKnots(me : mutable; aUKnots : mutable HArray1OfReal);
	UKnots (me) returns mutable HArray1OfReal;
	UKnotsValue (me; num : Integer) returns Real;
	NbUKnots (me) returns Integer;
	SetVKnots(me : mutable; aVKnots : mutable HArray1OfReal);
	VKnots (me) returns mutable HArray1OfReal;
	VKnotsValue (me; num : Integer) returns Real;
	NbVKnots (me) returns Integer;
	SetKnotSpec(me : mutable; aKnotSpec : KnotType);
	KnotSpec (me) returns KnotType;

	-- Specific Methods for ANDOR Field Data Access --

	SetWeightsData(me : mutable; aWeightsData : mutable HArray2OfReal);
	WeightsData (me) returns mutable HArray2OfReal;
	WeightsDataValue (me; num1 : Integer;  num2 : Integer) returns Real;
	NbWeightsDataI (me) returns Integer;
	NbWeightsDataJ (me) returns Integer;

fields

	bSplineSurfaceWithKnots : BSplineSurfaceWithKnots from StepGeom;
	rationalBSplineSurface : RationalBSplineSurface from StepGeom;

end BSplineSurfaceWithKnotsAndRationalBSplineSurface;
