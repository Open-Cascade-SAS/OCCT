-- Created on: 1992-02-21
-- Created by: Arnaud BOUZY
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



private class Analysis from ExprIntrp 

	---Purpose: 

uses Generator from ExprIntrp,
    GeneralExpression from Expr,
    GeneralRelation from Expr,
    GeneralFunction from Expr,
    StackOfGeneralExpression from ExprIntrp,
    StackOfGeneralRelation from ExprIntrp,
    StackOfGeneralFunction from ExprIntrp,
    StackOfInteger from TColStd,
    SequenceOfGeneralExpression from Expr,
    SequenceOfNamedFunction from ExprIntrp,
    SequenceOfNamedExpression from ExprIntrp,
    NamedFunction from Expr,
    NamedExpression from Expr,
    AsciiString from TCollection,
    StackOfNames from ExprIntrp
    
is

    Create
    returns Analysis;
    
    SetMaster(me : in out; agen : Generator)
    is static;
    
    Push(me : in out; exp : GeneralExpression)
    is static;
    
    PushRelation(me : in out; rel : GeneralRelation)
    is static;
    
    PushName(me : in out; name : AsciiString)
    is static;
    
    PushValue(me : in out; degree : Integer)
    is static;
    
    PushFunction(me : in out; func : GeneralFunction)
    is static;
    
    Pop(me : in out)
    returns GeneralExpression
    is static;
    
    PopRelation(me : in out)
    returns GeneralRelation
    is static;
    
    PopName(me : in out)
    returns AsciiString
    is static;
    
    PopValue(me: in out)
    returns Integer
    is static;
    
    PopFunction(me: in out)
    returns GeneralFunction
    is static;
    
    IsExpStackEmpty(me)
    returns Boolean
    is static;
    
    IsRelStackEmpty(me)
    returns Boolean
    is static;
    
    ResetAll(me : in out)
    is static;
    
    Use(me : in out; func : NamedFunction)
    is static;

    Use(me : in out; named : NamedExpression)
    is static;
        
    GetNamed(me : in out; name : AsciiString)
    returns NamedExpression
    is static;
    
    GetFunction(me : in out; name : AsciiString)
    returns NamedFunction
    is static;
    
fields

    myGEStack : StackOfGeneralExpression;
    myGRStack : StackOfGeneralRelation;
    myGFStack : StackOfGeneralFunction;
    myNameStack : StackOfNames;
    myValueStack : StackOfInteger;
    myFunctions : SequenceOfNamedFunction;
    myNamed : SequenceOfNamedExpression;
    myMaster : Generator;
    
end Analysis;
