-- File:        FaceSurface.cdl
-- Created:     Mon Dec  4 12:02:26 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWFaceSurface from RWStepShape

	---Purpose : Read & Write Module for FaceSurface

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     FaceSurface from StepShape,
     EntityIterator from Interface

is

	Create returns RWFaceSurface;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable FaceSurface from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : FaceSurface from StepShape);

	Share(me; ent : FaceSurface from StepShape; iter : in out EntityIterator);

end RWFaceSurface;
