-- Created on: 1994-11-04
-- Created by: Christian CAILLET
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



generic class Mapper from Transfer
    (TheKey    as  any;
     TheHasher as  any;
     TheInfo   as  any)
        inherits Finder

    ---Purpose : a Mapper defines a Finder for a specific input class
    --           its definition includes the value of the Key to be mapped,
    --           and the HashCoder associated to the class of the Key
    --           
    --           TheKey defines the class to be keyed
    --           TheHasher is the associated Hasher
    --           TheInfo   is an additionnal class which helps to provide
    --             informations on the value (template : see DataInfo)

uses CString

is

    Create (akey : any TheKey) returns mutable Mapper;
    ---Purpose : Creates a Mapper with a Value. This Value can then not be
    --           changed. It is used by the Hasher to compute the HashCode,
    --           which will then be stored for an immediate reading.

    Value (me) returns any TheKey  is static;
    ---Purpose : Returns the contained value
    ---C++ : return const &

    Equates (me; other : Finder) returns Boolean;
    ---Purpose : Specific testof equallity : defined as False if <other> has
    --           not the same true Type, else contents are compared (by
    --           C++ operator ==)

    ValueType    (me) returns Type  is redefined;
    ---Purpose : Returns the Type of the Value. By default, returns the
    --           DynamicType of <me>, but can be redefined

    ValueTypeName (me) returns CString  is redefined;
    ---Purpose : Returns the name of the Type of the Value. Default is name
    --           of ValueType, unless it is for a non-handled object

fields

    theval  : TheKey;

end Mapper;
