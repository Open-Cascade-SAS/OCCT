-- Created on: 1993-04-07
-- Created by: Laurent BUCHARD
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class IntersectionPoint from IntCurveSurface

    ---Purpose: Definition of an interserction point between a 
    --          curve and a surface. 

    ---Level: Public

   
uses
    Pnt                   from gp,
    TransitionOnCurve     from IntCurveSurface

is 

    Create
    	---Purpose: Empty Constructor.
    	returns IntersectionPoint from IntCurveSurface;
	
    Create(P     : Pnt        from gp; 
    	   USurf : Real       from Standard;
	   VSurf : Real       from Standard;
	   UCurv : Real       from Standard;
	   TrCurv: TransitionOnCurve   from IntCurveSurface)
	---Purpose: Create an IntersectionPoint.
	returns IntersectionPoint from IntCurveSurface;
	
    SetValues(me: in out;
             P     : Pnt        from gp; 
      	     USurf : Real       from Standard;
	     VSurf : Real       from Standard;
	     UCurv : Real       from Standard;
	     TrCurv: TransitionOnCurve   from IntCurveSurface)
	 ---Purpose: Set the fields of the current IntersectionPoint.
	 is static;
	 
    Values(me;
    	  P     : out Pnt        from gp; 
    	  USurf : out Real       from Standard;
	  VSurf : out Real       from Standard;
	  UCurv : out Real       from Standard;
	  TrCurv: out TransitionOnCurve   from IntCurveSurface)
	 ---Purpose: Get the fields of the current IntersectionPoint.
	 is static;
	 
    Pnt(me)
    	 ---Purpose: returns the geometric point.
         ---C++: return const & 
         ---C++: inline
         returns Pnt from gp
         is static;

    U(me)
    	 ---Purpose: returns the U parameter on the surface.
         ---C++: inline
         returns Real from Standard
         is static;

    V(me)
    	 ---Purpose: returns the V parameter on the surface.
         ---C++: inline
         returns Real from Standard
         is static;

    W(me)
    	 ---Purpose: returns the parameter on the curve.
         ---C++: inline
         returns Real from Standard
         is static;

    Transition(me)
    	 ---Purpose: returns the Transition of the point.
         ---C++: inline
         returns TransitionOnCurve from IntCurveSurface
         is static;


    Dump(me) 
    	 ---Purpose: Dump all the fields.
    	 is static;

fields

    myP       : Pnt      from gp;
    myUSurf   : Real     from Standard;
    myVSurf   : Real     from Standard;
    myUCurv   : Real     from Standard;
    myTrOnCurv: TransitionOnCurve   from IntCurveSurface;
 
end IntersectionPoint;

