-- Created on: 1996-01-22
-- Created by: Philippe MANGIN
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class DistributionOfEnergy from  FairCurve 
     inherits  FunctionSet from math

	---Purpose: Abstract class to use the Energy of an FairCurve

uses  Vector        from math, 
      FunctionSet   from math,
      HArray1OfReal  from TColStd,
      HArray1OfPnt2d from TColgp   



is

---    redefined methods

    NbVariables(me)
    	---Purpose: returns the number of variables of the function.

    returns Integer is redefined;

    
    NbEquations(me)
    	---Purpose: returns the number of equations of the function.

    returns Integer is redefined;

    
---    new methods
    Initialize( BSplOrder : Integer;
                FlatKnots :  HArray1OfReal;
		Poles     :  HArray1OfPnt2d;
    	    	DerivativeOrder : Integer;
    	    	NbValAux  : Integer = 0);
		
    SetDerivativeOrder(me :in out; DerivativeOrder : Integer); 
		    

fields

MyBSplOrder   : Integer is protected;
MyFlatKnots   : HArray1OfReal is  protected;
MyPoles       : HArray1OfPnt2d  is protected;
MyDerivativeOrder : Integer is protected;
MyNbVar       : Integer is protected;
MyNbEqua      : Integer is protected;
MyNbValAux    : Integer is protected;


end DistributionOfEnergy ;
