-- Created on: 1995-01-27
-- Created by: Marie Jose MARTZ
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class BRSolid from BRepToIGES inherits BREntity from BRepToIGES

    ---Purpose: This class implements the transfer of Shape Entities from Geom
    --          To IGES. These can be :
    --            . Vertex
    --            . Edge
    --            . Wire
  

uses

    Shape                from TopoDS,
    Solid                from TopoDS,
    CompSolid            from TopoDS,
    Compound             from TopoDS,
    IGESEntity           from IGESData,
    BREntity             from BRepToIGES    
    
is 
    
    Create returns BRSolid from BRepToIGES;


    Create (BR : BREntity from BRepToIGES)
    	returns BRSolid from BRepToIGES;    


    TransferSolid (me    : in out;
                   start : Shape from TopoDS)
    	 returns IGESEntity from IGESData;
    ---Purpose :  Transfert a Shape entity from TopoDS to IGES 
    --            this entity must be a Solid or a CompSolid or a Compound. 
    --            If this Entity could not be converted, this member returns a NullEntity.


    TransferSolid (me    : in out;
                   start : Solid from TopoDS)
    	 returns IGESEntity from IGESData;
    ---Purpose :  Transfert a Solid entity from TopoDS to IGES
    --            If this Entity could not be converted, this member returns a NullEntity.


    TransferCompSolid (me    : in out;
                       start : CompSolid from TopoDS)
    	 returns IGESEntity from IGESData;
    ---Purpose :  Transfert an CompSolid entity from TopoDS to IGES
    --            If this Entity could not be converted, this member returns a NullEntity.


    TransferCompound (me    : in out;
                      start : Compound from TopoDS)
    	 returns IGESEntity from IGESData;
    ---Purpose :  Transfert a Compound entity from TopoDS to IGES
    --            If this Entity could not be converted, this member returns a NullEntity.


end BRSolid;


