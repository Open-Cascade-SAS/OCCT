-- Created on: 1993-09-22
-- Created by: Didier PIFFAULT
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package BRepMesh

        ---Purpose: Instantiated   package for the   class of packages

        ---Level : Advanced.  
        --  All methods of all  classes will be advanced.


uses    Standard,
        gp,
        Bnd,
        TColStd,
        TColgp,
        GCPnts,
        BRepAdaptor,
        BRepTopAdaptor,
        TCollection,
        MMgt,
        TopoDS,
        TopAbs,
        TopExp,
        TopTools,
        Poly,
        Geom2d,
        GeomAbs,
        GeomAdaptor,
        TopLoc,
        SortTools,
        Plugin


is    enumeration DegreeOfFreedom is 
        Free,
        InVolume,
        OnSurface,
        OnCurve,
        Fixed,
        Frontier,
        Deleted;

      imported Status from BRepMesh;
       
      enumeration FactoryError is 
        FE_NOERROR,  
        FE_LIBRARYNOTFOUND,
        FE_FUNCTIONNOTFOUND,
        FE_CANNOTCREATEALGO
      end FactoryError;   
      
      class Vertex;

      class Edge;

	  imported Triangle from BRepMesh;
	  
      class ShapeTool;

      class Circ;

      deferred class DiscretRoot; 
      class DiscretFactory;
      --
      pointer PDiscretRoot to DiscretRoot from BRepMesh;
      --
      imported Delaun from BRepMesh;
      imported MapOfIntegerInteger from BRepMesh;
      imported MapOfInteger from BRepMesh;
      imported ListOfInteger from BRepMesh;
      imported BaseAllocator from BRepMesh;
      imported PairOfIndex from BRepMesh;
      imported CircleInspector from BRepMesh;
      imported CellFilter from BRepMesh;
      imported VertexInspector from BRepMesh;
      imported VertexCellFilter from BRepMesh;
      imported VectorOfVertex from BRepMesh;

      primitive PluginEntryType;

      class ComparatorOfVertexOfDelaun;
      class ComparatorOfIndexedVertexOfDelaun;
      class SelectorOfDataStructureOfDelaun;
      class DataStructureOfDelaun;
      class CircleTool;
      class VertexTool;
    
      class Array1OfVertexOfDelaun instantiates Array1 from TCollection
        (Vertex from BRepMesh);

      class HArray1OfVertexOfDelaun instantiates HArray1 from TCollection
        (Vertex from BRepMesh, Array1OfVertexOfDelaun);

      class HeapSortVertexOfDelaun instantiates  HeapSort from SortTools
        (Vertex from BRepMesh, Array1OfVertexOfDelaun,
        ComparatorOfVertexOfDelaun from BRepMesh);

      class HeapSortIndexedVertexOfDelaun instantiates  HeapSort from SortTools
        (Integer, Array1OfInteger from TColStd,
        ComparatorOfIndexedVertexOfDelaun from BRepMesh);

      class LinkHasherOfDataStructureOfDelaun instantiates MapHasher from TCollection
        (Edge from BRepMesh);
      class ElemHasherOfDataStructureOfDelaun instantiates MapHasher from TCollection
        (Triangle from BRepMesh);

      class DataMapOfIntegerListOfInteger     instantiates DataMap from TCollection
        (Integer from Standard, ListOfInteger from BRepMesh, MapIntegerHasher from TColStd);

      class IDMapOfLinkOfDataStructureOfDelaun  instantiates IndexedDataMap from TCollection
        (Edge from BRepMesh,
        PairOfIndex from BRepMesh,
        LinkHasherOfDataStructureOfDelaun);

      class IMapOfElementOfDataStructureOfDelaun instantiates IndexedMap from TCollection
        (Triangle from BRepMesh,
        ElemHasherOfDataStructureOfDelaun);

      class DataMapOfVertexInteger instantiates DataMap from TCollection
          (Vertex from TopoDS, Integer from Standard, ShapeMapHasher from TopTools);

      class ListOfVertex instantiates List from TCollection 
          (Vertex from  BRepMesh);
          
      class ListOfXY instantiates List from TCollection (XY from gp);

      class DataMapOfIntegerListOfXY  instantiates DataMap from TCollection
          (Integer from Standard, ListOfXY from BRepMesh, MapIntegerHasher from TColStd);


      class  VertexHasher  instantiates   MapHasher  from  TCollection(Vertex  from  BRepMesh);

      class IndexedMapOfVertex instantiates IndexedMap from TCollection 
          (Vertex from  BRepMesh,  VertexHasher from  BRepMesh);


      class BiPoint;
  
      class Array1OfBiPoint    instantiates Array1  from TCollection(BiPoint from BRepMesh);

      private class FastDiscretFace;
      
      class FastDiscret;
      
      class FaceAttribute;
  
      class DataMapOfFaceAttribute instantiates DataMap from TCollection
                                            (Face           from TopoDS,
                                             FaceAttribute  from BRepMesh,
                                             ShapeMapHasher from TopTools);
              
      private class Classifier;
      imported ClassifierPtr; -- smart pointer on Classifier

      class IncrementalMesh from BRepMesh;

         ---- classes moved from MeshShape
      class GeomTool;

      class DataMapOfIntegerPnt instantiates
          DataMap from TCollection   (Integer          from Standard,
                                      Pnt              from gp,
                                      MapIntegerHasher from TColStd);

      class PairOfPolygon;

      class DataMapOfShapePairOfPolygon instantiates 
      DataMap from TCollection(Shape          from TopoDS,
                               PairOfPolygon  from BRepMesh,
                               ShapeMapHasher from TopTools);

      Mesh(S: Shape from TopoDS; d: Real from Standard);
      ---Purpose: call to incremental mesh.

  
end BRepMesh;
