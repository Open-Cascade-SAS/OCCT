-- Created on: 1996-01-29
-- Created by: Kernel
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class BaseArray from DBC
inherits Storable from Standard

uses DBVArray from DBC

raises NullObject,
    NegativeValue,
    DimensionMismatch

is
    Create returns BaseArray;
    ---Purpose: Creates an BaseArray of NULL size
    
    Create (Size : Integer) returns BaseArray;
    ---Purpose: Creates  an BaseArray of lower bound 0 and
    --          upper bound <Size>-1.

    Create (BaseArray: BaseArray) returns BaseArray;
    ---Purpose: Creates an array which  is the copy of the given
    --          argument.

    ---C++: alias "  Standard_EXPORT virtual ~DBC_BaseArray();"

    Length (me) returns Integer is static ;
    ---C++: inline

    Upper (me) returns Integer is static;
    ---Purpose: Returns the upper bound
    ---C++: inline
              
    Lock (me) returns Address is static ;
    ---Purpose: Locks the array <me> in memory and 
    --          returns its virtual address
		

    Unlock (me) is static;
    ---Purpose: unlocks the array <me> from memory

fields
    mySize : Integer is protected;
    myData : DBVArray from DBC is protected;
end BaseArray;
