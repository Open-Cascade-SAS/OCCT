-- Created on: 1995-06-13
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class MakeCylindricalHole from BRepFeat inherits Builder from BRepFeat

        ---Purpose: Provides a tool to make cylindrical holes on a shape.

uses Shape                from TopoDS,
     Face                 from TopoDS,
     Ax1                  from gp,
     Status               from BRepFeat


raises NotDone from StdFail,
       ConstructionError from Standard

is

    Create
        ---Purpose: Empty constructor.
            returns MakeCylindricalHole from BRepFeat;
        ---C++: inline


    Init(me: in out; Axis: Ax1 from gp)
        ---Purpose: Sets the axis of the hole(s).
        ---C++: inline
            is static;


    Init(me: in out; S: Shape from TopoDS; Axis: Ax1 from gp)
        ---Purpose: Sets the shape and  axis on which hole(s)  will be
        --          performed.  
        ---C++: inline
            is static;


    Perform(me: in out; Radius: Real from Standard)
        ---Purpose: Performs every  holes of   radius  <Radius>.  This
        --          command  has the  same effect as   a cut operation
        --          with an  infinite cylinder   defined by the  given
        --          axis and <Radius>.

            raises ConstructionError from Standard
        -- The exception is raised when no shape or no axis is defined.
            is static;


    Perform(me: in out; Radius: Real from Standard; 
                        PFrom,PTo: Real from Standard;
                        WithControl: Boolean from Standard = Standard_True)
        ---Purpose: Performs evry   hole  of  radius  <Radius> located
        --          between PFrom  and  PTo  on the  given  axis.   If
        --          <WithControl> is set  to Standard_False no control
        --          are  done  on   the  resulting  shape   after  the
        --          operation is performed.

            raises ConstructionError from Standard
        -- The exception is raised when no shape or no axis is defined.
            is static;


    PerformThruNext(me: in out; 
                     Radius: Real from Standard;
                     WithControl: Boolean from Standard = Standard_True)
        ---Purpose: Performs the first hole of radius <Radius>, in the
        --          direction of  the defined axis. First hole signify
        --          first encountered after the origin of the axis. If
        --          <WithControl> is set  to Standard_False no control
        --          are  done  on   the  resulting  shape   after  the
        --          operation is performed. 

            raises ConstructionError from Standard
        -- The exception is raised when no shape or no axis is defined.
            is static;


    PerformUntilEnd(me: in out; 
                     Radius: Real from Standard;
                     WithControl: Boolean from  Standard = Standard_True)
        ---Purpose: Performs  evry  holes of  radius  <Radius> located
        --          after  the   origin  of   the given    axis.    If
        --          <WithControl> is  set to Standard_False no control
        --          are done   on   the  resulting  shape   after  the
        --          operation is performed.

            raises ConstructionError from Standard
        -- The exception is raised when no shape or no axis is defined.
            is static;


    PerformBlind(me: in out; 
                  Radius: Real from Standard; 
                  Length: Real from Standard;
                  WithControl: Boolean from  Standard = Standard_True)
        ---Purpose: Performs a  blind   hole of radius    <Radius> and
        --          length <Length>.  The length is  measured from the
        --          origin of the given  axis. If <WithControl> is set
        --          to  Standard_False no  control  are done after the
        --          operation is performed.

            raises ConstructionError from Standard
        -- The exception is raised when no shape or no axis is defined.
            is static;


    Status(me)
        ---Purpose: Returns the status after a hole is performed.
        ---C++: inline
            returns Status from BRepFeat
        is static;


--- Redefinition of BRepBuilderAPI_MakeShape methods
--  
--  

    Build(me:out);
        ---Purpose: Builds the    resulting shape  (redefined     from
        --          MakeShape). Invalidates the  given parts  of tools
        --          if  any,   and performs the  result   of the local
        --          operation.


--- Private implementation method


    Validate(me: in out)
    
            returns Status from BRepFeat
        is static private;


fields

    myAxis    : Ax1                  from gp;
    myAxDef   : Boolean              from Standard;
    myStatus  : Status               from BRepFeat;
    myIsBlind : Boolean              from Standard;
    myValidate: Boolean              from Standard;
    myTopFace : Face                 from TopoDS;
    myBotFace : Face                 from TopoDS;


end MakeCylindricalHole;
