-- File:	RWStepRepr_RWProductDefinitionShape.cdl
-- Created:	Mon Jul  3 16:29:03 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class RWProductDefinitionShape from RWStepRepr

    ---Purpose: Read & Write tool for ProductDefinitionShape

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    ProductDefinitionShape from StepRepr

is
    Create returns RWProductDefinitionShape from RWStepRepr;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : ProductDefinitionShape from StepRepr);
	---Purpose: Reads ProductDefinitionShape

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: ProductDefinitionShape from StepRepr);
	---Purpose: Writes ProductDefinitionShape

    Share (me; ent : ProductDefinitionShape from StepRepr;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWProductDefinitionShape;
