-- Created on: 1997-03-03
-- Created by: Jean-Pierre COMBE
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class IdenticRelation from AIS inherits Relation from AIS

	---Purpose: Constructs a constraint by a relation of identity
    	-- between two or more datums figuring in shape
    	-- Interactive Objects.

uses
     Shape                 from TopoDS,
     Vertex                from TopoDS,
     Wire                  from TopoDS,
     Presentation          from Prs3d,
     PresentationManager3d from PrsMgr,
     Selection             from SelectMgr,
     Projector             from Prs3d,
     Transformation         from Geom,
     Plane                 from Geom,
     Curve                 from Geom,
     Line                  from Geom,
     Circle                from Geom,
     Ellipse               from Geom,
     Pnt                   from gp,
     Dir                   from gp

is
    Create(FirstShape  : Shape from TopoDS;
    	   SecondShape : Shape from TopoDS;
	   aPlane      : Plane from Geom)
    returns mutable IdenticRelation from AIS;
    	---Purpose:
    	--   Initializes the relation of identity between the two
    	-- entities, FirstShape and SecondShape. The plane
    	-- aPlane is initialized in case a visual reference is
    	-- needed to show identity.
    
    IsMovable(me) returns Boolean from Standard 
        ---C++: inline       
    	---Purpose:
    	-- Returns true if the interactive object is movable.
    is redefined;     
    
-- Methods from PresentableObject

    Compute(me            : mutable;
    	    aPresentationManager: PresentationManager3d from PrsMgr;
    	    aPresentation : mutable Presentation from Prs3d;
    	    aMode         : Integer from Standard= 0) 
    is redefined private;
    
    Compute(me:mutable;
    	        aProjector: Projector from Prs3d;
                aPresentation: mutable Presentation from Prs3d)
    is redefined static private;     

    Compute(me            : mutable;
    	    aProjector    : Projector from Prs3d;
    	    aTrsf         : Transformation from Geom;
	    aPresentation : mutable Presentation from Prs3d)
    is redefined;
    ---Purpose: computes the presentation according to a point of view
    --          given by <aProjector>. 
    --          To be Used when the associated degenerated Presentations 
    --          have been transformed by <aTrsf> which is not a Pure
    --          Translation. The HLR Prs can't be deducted automatically
    --          WARNING :<aTrsf> must be applied
    --           to the object to display before computation  !!!

-- Methods from SelectableObject

    ComputeSelection(me         : mutable;
    	    	     aSelection : mutable Selection from SelectMgr;
    	    	     aMode      : Integer from Standard)
    is redefined private;

--
--     Computation private methods
--

    ComputeOneEdgeOVertexPresentation(me: mutable;
    	    	    	       aPresentation : mutable Presentation from Prs3d)
    is private;

    ComputeTwoEdgesPresentation(me: mutable;
    	    	    	       aPresentation : mutable Presentation from Prs3d)
    is private;
    
    ComputeTwoLinesPresentation(me: mutable;
    	    	    	       aPresentation : mutable Presentation from Prs3d; 
			       aLin    : Line from Geom;
    	    	    	       Pnt1On1 : in out Pnt  from gp;
			       Pnt2On1 : in out Pnt  from gp;
			       Pnt1On2 : in out Pnt  from gp;
			       Pnt2On2 : in out Pnt  from gp;
			       isInf1  : Boolean from Standard;
			       isInf2  : Boolean from Standard)
    is private; 
    
    ComputeTwoCirclesPresentation(me: mutable;
    	    	    	       aPresentation : mutable Presentation from Prs3d; 
			       aCircle : Circle from Geom;
    	    	    	       Pnt1On1 : Pnt    from gp;
			       Pnt2On1 : Pnt    from gp;
			       Pnt1On2 : Pnt    from gp;
			       Pnt2On2 : Pnt    from gp)
    is private;        
    
    -- jfa 17/10/2000
    ComputeAutoArcPresentation(me: mutable;
    	    	    	       aCircle : Circle from Geom;
    	    	    	       firstp  : Pnt from gp;
    	    	    	       lastp   : Pnt from gp;
    	    	    	       isstatic: Boolean from Standard = Standard_False)
    	---Purpose: Computes the presentation of the identic constraint
    	--          between 2 arcs in the case of automatic presentation 
    is private; 

    ComputeNotAutoCircPresentation(me: mutable;
    	    	    	    	   aCircle : Circle from Geom)
    	---Purpose: Computes the presentation of the identic constraint
    	--          between 2 circles in the case of non automatic presentation 
    is private; 
    
    ComputeNotAutoArcPresentation(me: mutable;
    	    	    	    	  aCircle : Circle from Geom;
    	    	    	    	  pntfirst: Pnt from gp;
    	    	    	    	  pntlast : Pnt from gp)
    	---Purpose: Computes the presentation of the identic constraint
    	--          between 2 arcs in the case of non automatic presentation 
    is private; 
    -- jfa 17/10/2000 end
    
    -- jfa 10/10/2000
    ComputeTwoEllipsesPresentation(me: mutable;
    	    	    		   aPrs    : mutable Presentation from Prs3d; 
			           anEll   : Ellipse from Geom;
    	    	    	           Pnt1On1 : Pnt    from gp;
			           Pnt2On1 : Pnt    from gp;
			           Pnt1On2 : Pnt    from gp;
			           Pnt2On2 : Pnt    from gp)
    is private;        
    -- jfa 10/10/2000 end
    
    -- jfa 18/10/2000
    ComputeAutoArcPresentation(me: mutable;
    	    	    	       theEll  : Ellipse from Geom;
    	    	    	       firstp  : Pnt from gp;
    	    	    	       lastp   : Pnt from gp;
    	    	    	       isstatic: Boolean from Standard = Standard_False)
    	---Purpose: Computes the presentation of the identic constraint
    	--          between 2 arcs in the case of automatic presentation 
    is private; 

    ComputeNotAutoElipsPresentation(me: mutable;
    	    	    	    	    theEll : Ellipse from Geom)
    	---Purpose: Computes the presentation of the identic constraint
    	--          between 2 ellipses in the case of non automatic presentation 
    is private; 

    ComputeNotAutoArcPresentation(me: mutable;
    	    	    	    	  theEll  : Ellipse from Geom;
    	    	    	    	  pntfirst: Pnt from gp;
    	    	    	    	  pntlast : Pnt from gp)
    	---Purpose: Computes the presentation of the identic constraint
    	--          between 2 arcs in the case of non automatic presentation 
    is private; 
    -- jfa 18/10/2000 end
    
    ComputeTwoVerticesPresentation(me: mutable; 
    	    	    	           aPresentation : mutable Presentation from Prs3d)
    is private;    

    ComputeSegSize(me)
    returns Real from Standard
    is private;
    
    ComputeDirection(me; aWire    : Wire    from TopoDS;
    	    	    	 aVertex  : Vertex  from TopoDS;
    	    	    	 aDir     : out Dir from gp)
    returns Boolean from Standard
    is private;

    ComputeLineDirection(me; aLin        : Line from Geom;
    	    	    	     anExtremity : Pnt from gp)
    returns Dir from gp
    is private;
    
    ComputeCircleDirection(me; aCirc           : Circle from Geom;
    	                       ConnectedVertex : Vertex from TopoDS)
    returns Dir from gp
    is private;
        
fields 

    isCircle    : Boolean from Standard;
    myFAttach   : Pnt     from gp;
    mySAttach   : Pnt     from gp;
    myCenter    : Pnt     from gp;

end IdenticRelation;
