-- Created on: 1992-09-28
-- Created by: Remi GILET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MakeSegment from GC inherits Root from GC

    --- Purpose: Implements construction algorithms for a line
    -- segment in 3D space.
    -- Makes a segment of Line from the 2 points <P1> and <P2>.
    -- The result is a Geom_TrimmedCurve curve.
    -- A MakeSegment object provides a framework for:
    -- -   defining the construction of the line segment,
    -- -   implementing the construction algorithm, and
    -- -   consulting the results. In particular, the Value
    --   function returns the constructed line segment.

uses Pnt          from gp,
     Real         from Standard,
     Lin          from gp,
     TrimmedCurve from Geom

raises NotDone from StdFail

is

Create(P1, P2 : Pnt from gp ) returns MakeSegment;
    	---Purpose: Make a segment of Line from the 2 points <P1> and <P2>.
    	--          It returns NullObject if <P1> and <P2> are confused.
	
Create(Line   : Lin  from gp       ;
       U1, U2 : Real from Standard ) returns MakeSegment;
    	---Purpose: Make a segment of Line from the line <Line1> 
    	--          between the two parameters U1 and U2.
    	--          It returns NullObject if <U1> is equal <U2>.

Create(Line   : Lin  from gp       ;
       Point  : Pnt  from gp       ;
       Ulast  : Real from Standard ) returns MakeSegment;
    	---Purpose: Make a segment of Line from the line <Line1> 
    	--          between the point <Point> and the parameter Ulast.
    	--          It returns NullObject if <U1> is equal <U2>.

Create(Line : Lin  from gp ;
       P1   : Pnt  from gp ;
       P2   : Pnt  from gp ) returns MakeSegment;
    	---Purpose: Make a segment of Line from the line <Line1> 
    	--          between the two points <P1> and <P2>.
    	--          It returns NullObject if <U1> is equal <U2>.

Value(me) returns TrimmedCurve from Geom
    raises NotDone
    is static;
    	---Purpose: Returns the constructed line segment.
    	---C++: return const&
        ---C++: alias "operator const Handle(Geom_TrimmedCurve)& () const { return Value(); }"

fields

    TheSegment : TrimmedCurve from Geom;
    --The solution from Geom.
    
end MakeSegment;
