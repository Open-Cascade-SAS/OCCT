-- Created on: 1994-12-12
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class Copy from BRepBuilderAPI inherits ModifyShape from BRepBuilderAPI

	---Purpose: Duplication of a shape.
    	-- A Copy object provides a framework for:
    	-- -   defining the construction of a duplicate shape,
    	-- -   implementing the construction algorithm, and
    	-- -   consulting the result.
        
uses
    Shape             from TopoDS,
    Face              from TopoDS,
    ShapeModification from BRepBuilderAPI,
    ListOfShape       from TopTools


is

    Create
	---Purpose: Constructs an empty copy framework. Use the function
    	-- Perform to copy shapes.
       	returns Copy from BRepBuilderAPI;


    Create(S: Shape from TopoDS; copyGeom: Boolean = Standard_True)
	---Purpose: Constructs a copy framework and copies the shape S.
    	-- Use the function Shape to access the result.
    	-- If copyGeom is False, only topological objects will be copied, while 
    	-- geometry will be shared with original shape.
    	-- Note: the constructed framework can be reused to copy
    	-- other shapes: just specify them with the function Perform.
    	returns Copy from BRepBuilderAPI;


    Perform(me: in out; S: Shape from TopoDS; copyGeom: Boolean = Standard_True)
	---Purpose: Copies the shape S.
    	-- Use the function Shape to access the result.
    	-- If copyGeom is False, only topological objects will be copied, while 
    	-- geometry will be shared with original shape.
    	is static;


end Copy;
