-- Created on: 1993-08-19
-- Created by: Laurent BUCHARD
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



generic class QuadricCurveFunc from IntCurveSurface ( 
    	TheQuadric       as any;    -- as Quadric   from IntCurveSurface
	TheCurve         as any;    
        TheCurveTool     as any)    -- as CurveTool from Adaptor3d
 
inherits  FunctionWithDerivative   from math


        
        ---Purpose: Implements     the function  Q(w)   and its  first
        --          derivative used  by FunctionAllRoots  to  find the
        --          areas where  the distance  between the quadric and
        --          the   parametric   curves is    less than a  given
        --          tolerance.
        --          
    	--   where Q(X,Y,Z) =  0   is the  implicit expression  of   a
    	--   quadric and (X(w),Y(w),Z(w))  the point of parameter w on
    	--   a parametric curve.
    	--

is

    Create(Q: TheQuadric; C:TheCurve)
    
    	---Purpose: Create the function.
    	--          
    	returns QuadricCurveFunc from IntCurveSurface;
	
	
	
    Value(me: in out; Param: Real from Standard; F: out Real from Standard)

      	---Purpose: Computes the value of the signed  distance between
      	--          the  implicit surface and  the point  at parameter
      	--          Param on the parametrised curve.
      	--          Value always returns True. 

    	returns Boolean from Standard
        is redefined static;
	
	
    Derivative(me: in out; Param: Real from Standard; 
               D: out Real from Standard)
	       
    	---Purpose: Computes the derivative of the previous function at
    	--          parameter Param.
    	--          Derivative always returns True.

    	returns Boolean from Standard
        is redefined static;
	
	
    Values(me: in out; Param: Real from Standard; F,D: out Real from Standard)
    
    	---Purpose: Computes the value and the derivative of the function.
    	--          returns True. 

    	returns Boolean from Standard
    	is redefined static;


fields 

    myQuadric       : TheQuadric;    
    myCurve         : TheCurve;
		  
end QuadricCurveFunc;

