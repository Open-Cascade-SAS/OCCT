-- Created on: 1993-10-29
-- Created by: Christophe MARION
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PolyShellData from HLRAlgo inherits TShared from MMgt
	---Purpose: All the PolyData of a Shell

uses
    Address            from Standard,
    Boolean            from Standard,
    Integer            from Standard,
    Array1OfTransient  from TColStd,
    HArray1OfTransient from TColStd,
    ListOfBPoint       from HLRAlgo

is
    Create(nbFace : Integer from Standard)
    returns PolyShellData from HLRAlgo;

    UpdateGlobalMinMax(me        : mutable;
                       TotMinMax : Address from Standard)
    is static;
    
    UpdateHiding(me       : mutable;
  	         nbHiding : Integer from Standard)
    is static;

    Hiding(me) returns Boolean from Standard
	---C++: inline
    is static;

    PolyData(me : mutable) 
	---C++: return &
	---C++: inline
    returns Array1OfTransient from TColStd
    is static;

    HidingPolyData(me : mutable) 
	---C++: return &
	---C++: inline
    returns Array1OfTransient from TColStd
    is static;

    Edges(me : mutable) 
	---C++: return &
	---C++: inline
    returns ListOfBPoint from HLRAlgo
    is static;

    Indices(me : mutable) returns Address from Standard
    	---C++: inline
    is static;

fields
    myMinMax    : Integer            from Standard[2];
    myPolyg     : Array1OfTransient  from TColStd;
    myHPolHi    : HArray1OfTransient from TColStd;
    mySegList   : ListOfBPoint       from HLRAlgo;

end PolyShellData;
