-- File:	IntImp_CSFunction.cdl
-- Created:	Mon Feb 14 11:50:41 1994
-- Author:	Jacques GOUSSARD
--		<jag@topsn2>
---Copyright:	 Matra Datavision 1994



deferred generic class CSFunction from IntImp 
    (ThePSurface as any;
     TheCurve as any
    )
    
inherits FunctionSetWithDerivatives from math

      	---Purpose: This class is the template function for the intersection
      	--          between a curve and a surface.
      	--          It is possible to implement such a function with an
      	--          instantiation of :
      	--           - ZerCSParFunc for the intersection between a 3d curve
      	--             and a surface.
      	--           - ZerCOnSSParFunc for the intersection between a curve
      	--             on surface and another surface.
    	

uses Vector from math,
     Matrix from math,
     Pnt from gp

is
	    
    NbVariables(me) returns Integer from Standard
    ---Purpose: Returns 3.
    is static;
    
    NbEquations(me) returns Integer from Standard
    ---Purpose: Returns 3.
    is static;
    
    Value(me : in out; X : in Vector from math;
    	    	       F : out Vector from math)
    returns Boolean from Standard
    is static;
    
    Derivatives(me : in out;X : in  Vector from math;
    	    	    	    D : out Matrix from math)
    returns Boolean from Standard
    is static;
    
    Values(me : in out;
    	   X  : in Vector from math;
	   F  : out Vector from math; D: out Matrix from math)
    returns Boolean from Standard
    is static;

    Point(me)
    	---C++: return const&
    	returns Pnt from gp
    	is static;
    
    Root(me) returns Real from Standard
    is static;
    
    AuxillarSurface(me)
    	---C++: return const&
    	returns ThePSurface
    	is static;

    AuxillarCurve(me)
    	---C++: return const&
    	returns TheCurve
    	is static;
     
end CSFunction;
