-- Created on: 1998-03-12
-- Created by: Pierre BARRAS
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class SplitCurve2d from ShapeUpgrade inherits SplitCurve from ShapeUpgrade

    	---Purpose: Splits a 2d curve with a criterion.
    
uses     
    Curve          from Geom2d,
    HArray1OfCurve from TColGeom2d
   
is 
 
    Create returns mutable SplitCurve2d from ShapeUpgrade;
    	---Purpose: Empty constructor.

    Init (me: mutable; C: Curve from  Geom2d);
       	---Purpose: Initializes with pcurve with its first and last parameters.
	
    Init (me: mutable; C          : Curve from  Geom2d;
    	    	       First, Last: Real);
       	---Purpose: Initializes with pcurve with its parameters.
	
    Build (me: mutable; Segment: Boolean) is redefined;
       ---Purpose: If Segment is True, the result is composed with
       --  segments of the curve bounded by the SplitValues.  If
       --  Segment is False, the result is composed with trimmed
       --  Curves all based on the same complete curve.
       --  
    GetCurves(me) returns HArray1OfCurve from TColGeom2d;
       ---C++: return const &
       
fields 
 
    myCurve          : Curve from Geom2d is protected;
    myResultingCurves: HArray1OfCurve from TColGeom2d is protected;
    
end;
    
