-- Created on: 1997-10-22
-- Created by: Jean-Louis Frenkel
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MetaData from CDM inherits Transient from Standard

uses ExtendedString from TCollection,Document from CDM,MetaDataLookUpTable from CDM, DocumentPointer from CDM,
Application from CDM
raises NoSuchObject from Standard

is
    
    Create(aFolder,aName, aPath: ExtendedString from TCollection;
           aFileName: ExtendedString from TCollection; ReadOnly:Boolean from Standard)
    returns  MetaData from CDM is private;

    Create(aFolder,aName, aPath, aVersion: ExtendedString from TCollection;
           aFileName: ExtendedString from TCollection; ReadOnly:Boolean from Standard)
    returns  MetaData from CDM is private;



    LookUp(myclass; aFolder,aName, aPath: ExtendedString from TCollection; 
           aFileName: ExtendedString from TCollection; ReadOnly:Boolean from Standard)
    returns  MetaData from CDM;

    LookUp(myclass; aFolder,aName, aPath, aVersion: ExtendedString from TCollection; aFileName: ExtendedString from TCollection; ReadOnly:Boolean from Standard)
    returns  MetaData from CDM;




    IsRetrieved(me) returns Boolean from Standard;

    Document(me) returns Document from CDM;
    
    Folder(me) returns ExtendedString from TCollection;
    ---Purpose: returns the folder in which the meta-data has to be created 
    --          or has to be found.
    --          
    Name(me) returns ExtendedString from TCollection;
    ---Purpose: returns the name under which the meta-data has to be created 
    --          or has to be found.
    --          
    
    Version(me) returns ExtendedString from TCollection
    ---Purpose: returns the version under which the meta-data has to be found.  
    -- Warning: raises NoSuchObject from Standard if no Version has been defined

    raises NoSuchObject from Standard;

    HasVersion(me) returns Boolean from Standard;
    ---Purpose: indicates that the version has to be taken into account when
    --          searching the corresponding meta-data.

    FileName(me) returns ExtendedString from TCollection;
    ---Category: programming facility
    --           
    Print(me; anOStream:  in out OStream from Standard)
    returns OStream from Standard;
    ---C++: return &
    ---C++: alias "Standard_OStream& operator << (Standard_OStream& anOStream);"
    --      

    Path(me) returns ExtendedString from TCollection;
    
   
    ---Category: methods to modify the metadata.
    --           
    SetDocument(me: mutable; aDocument: Document from CDM)
    is private;

    UnsetDocument(me: mutable);

    LookUpTable(myclass) returns MetaDataLookUpTable from CDM
    is private;
    ---C++: return const&
    --      
    DocumentVersion(me: mutable; anApplication: Application from CDM) returns Integer from Standard
    is private;
    
    IsReadOnly(me) returns Boolean from Standard;

    SetIsReadOnly(me: mutable);
    
    UnsetIsReadOnly(me: mutable);
    
fields
    myIsRetrieved: Boolean from Standard;
    myDocument: DocumentPointer from CDM;
    myFolder: ExtendedString from TCollection;
    myName: ExtendedString from TCollection;

    myVersion: ExtendedString from TCollection;
    myHasVersion: Boolean from Standard;

    myFileName: ExtendedString from TCollection;
    myPath: ExtendedString from TCollection;


    myDocumentVersion: Integer from Standard;
    
    myIsReadOnly: Boolean from Standard;

 friends SetMetaData from class Document from CDM(me: mutable; aMetaData: MetaData from CDM),
        class Reference from CDM,
        SetDocumentVersion from class Application from CDM(me; aDocument: Document from CDM; aMetaData: MetaData from CDM)
end MetaData from CDM;
