-- Created on: 1992-05-05
-- Created by: Remi GILET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


package GCE2d

uses gp,
     Geom2d,
     gce,
     StdFail


    ---Level : Public. 
    --  All methods of all  classes will be public.



is

private deferred class Root;

---------------------------------------------------------------------------
--          Constructions of 2d geometrical elements from Geom2d.
---------------------------------------------------------------------------

class MakeLine;
    	---Purpose: Makes a Line from Geom2d.

class MakeCircle;
    	---Purpose: Makes a Circle from Geom2d.

class MakeHyperbola;
    	---Purpose: Makes an hyperbola from Geom2d.

class MakeEllipse;
    	---Purpose: Makes an Ellipse from Geom2d.

class MakeParabola;
    	---Purpose: Makes a parabola from Geom2d.

class MakeSegment;
    	---Purpose: Makes a segment of Line (TrimmedCurve from Geom2d).

class MakeArcOfCircle;
    	---Purpose: Makes an arc of circle (TrimmedCurve from Geom2d).

class MakeArcOfEllipse;
    	---Purpose: Makes an arc of ellipse (TrimmedCurve from Geom2d).

class MakeArcOfParabola;
    	---Purpose: Makes an arc of parabola (TrimmedCurve from Geom2d).

class MakeArcOfHyperbola;
    	---Purpose: Makes an arc of hyperbola (TrimmedCurve from Geom2d).

---------------------------------------------------------------------------
--              Constructions of Transformation from Geom2d.
---------------------------------------------------------------------------

class MakeTranslation;
    	---Purpose: Returns a translation transformation.
 
class MakeMirror;
    	---Purpose: Returns a symmetry transformation. 

class MakeRotation;
    	---Purpose: Returns a rotation transformation.

class MakeScale;
    	---Purpose: Returns a scaling transformation.

    
end GCE2d;



