-- Created on: 1992-05-06
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PntOn2S from IntSurf 

	---Purpose: This class defines the geometric informations
	--          for an intersection point between 2 surfaces :
	--          The coordinates ( Pnt from gp ), and two
	--          parametric coordinates.


uses Pnt from gp

is


    Create
    
	---Purpose: Empty constructor.
    
    	returns PntOn2S from IntSurf;


    SetValue(me: in out; Pt: Pnt from gp)
    
	---Purpose: Sets the value of the point in 3d space.

	---C++: inline

    	is static;


    SetValue(me: in out; Pt: Pnt from gp; OnFirst: Boolean from Standard;
             U,V: Real from Standard)
    
	---Purpose: Sets the values of the point in 3d space, and
	--          in the parametric space of one of the surface.

    	is static;


    SetValue(me: in out; Pt: Pnt from gp; U1,V1,U2,V2: Real from Standard)
    
	---Purpose: Sets the values of the point in 3d space, and
	--          in the parametric space of each surface.

	---C++: inline

    	is static;


    SetValue(me: in out; OnFirst: Boolean from Standard;
                         U,V: Real from Standard)
    
	---Purpose: Set the values of the point in the parametric
	--          space of one of the surface.

    	is static;


    SetValue(me: in out; U1,V1, U2, V2: Real from Standard)
    
	---Purpose: Set the values of the point in the parametric
	--          space of one of the surface.

	---C++: inline

    	is static;


    Value(me)
    
	---Purpose: Returns the point in 3d space.

    	returns Pnt from gp
	---C++: return const&
	---C++: inline

	is static;



    ParametersOnS1(me; U1,V1: out Real from Standard)

	---Purpose: Returns the parameters of the point on the first surface.

	---C++: inline

    	is static;


    ParametersOnS2(me; U2,V2: out Real from Standard)

	---Purpose: Returns the parameters of the point on the second surface.

	---C++: inline

    	is static;


    Parameters(me; U1,V1,U2,V2: out Real from Standard)

	---Purpose: Returns the parameters of the point on both surfaces.

	---C++: inline

    	is static;


fields

    pt  : Pnt     from gp;
    u1  : Real    from Standard;
    v1  : Real    from Standard;
    u2  : Real    from Standard;
    v2  : Real    from Standard;

end PntOn2S;
