-- Created on: 1995-12-01
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DrawableC2D from TestTopOpeDraw inherits Curve2d from DrawTrSurf

uses  

    Interpretor from Draw,
    Curve from Geom2d,
    Color from Draw,
    Display from Draw,
    Text2D from Draw,
    CString from Standard,
    Pnt2d from gp

is

    Create (C : Curve from Geom2d; CColor : Color from Draw)
    returns DrawableC2D from TestTopOpeDraw;

    Create (C : Curve from Geom2d; CColor : Color from Draw;
    	    Text : CString; TextColor : Color from Draw)
    returns DrawableC2D from TestTopOpeDraw;

    Create (C : Curve from Geom2d; CColor : Color from Draw;
    	    Text : CString; TextColor : Color from Draw;
    	    Discret : Integer;
    	    DispOrigin : Boolean = Standard_True;
            DispCurvRadius : Boolean = Standard_False;
	    RadiusMax : Real = 1.0e3;
	    RatioOfRadius : Real = 0.1)
    returns DrawableC2D from TestTopOpeDraw;

    Pnt2d(me) returns Pnt2d from gp is virtual;
    
    ChangePnt2d(me : mutable; P : Pnt2d);
    
    ChangeCurve(me : mutable; C : Curve from Geom2d);
    
    ChangeText(me : mutable; T : CString from Standard);
    
    Name(me : mutable; N : CString) is redefined;
    
    Whatis(me; I : in out Interpretor from Draw) is redefined;
    ---Purpose: For variable whatis command.

    DrawOn(me; dis : in out Display from Draw) is redefined;
    
fields

    myText2D : Text2D from Draw is protected;
    myText : CString from Standard is protected;
    myTextColor : Color from Draw;

end DrawableC2D;
