-- File:	PGeom_OffsetCurve.cdl
-- Created:	Mon Mar  1 13:22:09 1993
-- Author:	Philippe DAUTRY
--		<fid@phylox>
-- Copyright:	 Matra Datavision 1993


class OffsetCurve from PGeom inherits Curve from PGeom

        ---Purpose :
        --  This class implements the basis services for an offset curve
        --  in 3D space.
        --  
	---See Also : OffsetCurve from Geom.

uses Dir      from gp,
     Curve    from PGeom


is
    

  Create returns mutable OffsetCurve from PGeom;
    ---Purpose: Creates an OffsetCurve with default values.
    	---Level: Internal 


  Create (
    	    aBasisCurve : Curve from PGeom;
    	    aOffsetValue : Real from Standard;
    	    aOffsetDirection : Dir from gp)
     returns mutable OffsetCurve from PGeom;
        ---Purpose : <aBasisCurve> is  the basis curve, <aOffsetValue>
        --         is the distance between <me> and the basis curve at
        --         any point.    <aOffsetDirection>  defines the fixed
        --         reference direction (offset direction).
    	---Level: Internal 


  BasisCurve (me : mutable; aBasisCurve : Curve from PGeom);
	---Purpose: Set the field basisCurve with <aBasisCurve>.
    	---Level: Internal 
      

  BasisCurve (me) returns Curve from PGeom; 
        ---Purpose : The basis curve can be an offset curve.
    	---Level: Internal 


  OffsetDirection (me : mutable; aOffsetDirection : Dir from gp);
        ---Purpose : Set the value of  the field offsetDirection with
        --  <aOffsetDirection>.
    	---Level: Internal 


  OffsetDirection (me)  returns Dir from gp;
        ---Purpose : Returns the direction of offset.
    	---Level: Internal 


  OffsetValue (me : mutable; aOffsetValue : Real from Standard);
        ---Purpose : Set the field offsetValue with <aOffsetValue>.
    	---Level: Internal 


  OffsetValue (me) returns Real from Standard;
        ---Purpose : Returns the value of the field offsetValue.
    	---Level: Internal 


fields

  basisCurve      : Curve from PGeom;
  offsetDirection : Dir from gp;
  offsetValue     : Real from Standard;

end;
