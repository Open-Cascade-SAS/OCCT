-- Created on: 1993-02-22
-- Created by: Philippe DAUTRY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class CartesianPoint from PGeom inherits Point from PGeom

        ---Purpose : Point defined  in  3D space with its 3  cartesian
        --         coordinates X, Y, Z.
        --         
    	---See Also : CartesianPoint from Geom.

uses Pnt from gp

is


  Create returns mutable CartesianPoint from PGeom;
        ---Purpose : Returns a CartesianPoint with default values..
    	---Level: Internal 


  Create (aPnt : Pnt from gp) returns mutable CartesianPoint from PGeom;
        ---Purpose : Returns a CartesianPoint built with <aPnt>.
    	---Level: Internal 


  Pnt (me : mutable; aPnt : Pnt from gp);
        ---Purpose : Set the field pnt.
    	---Level: Internal 


  Pnt (me)  returns Pnt;
        ---Purpose : Returns the value of the field pnt.
    	---Level: Internal 


fields

    pnt : Pnt from gp;

end;
