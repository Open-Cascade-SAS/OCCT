-- Created on: 1997-04-29
-- Created by: Stagiaire Francois DUMONT
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class CompCurveToBSplineCurve from Geom2dConvert 

	    ---Purpose: Concat sevral curve in an BSplineCurve

uses
 ParameterisationType from Convert,
 BoundedCurve from Geom2d,
 BSplineCurve from Geom2d

--raises

is

    Create (BasisCurve : BoundedCurve from Geom2d; 
     	    Parameterisation : ParameterisationType from Convert 
    	    	       =  Convert_TgtThetaOver2)
	    ---Purpose: Initialize the algorithme with one curve
	    --        - Parameterisation is used to convert 
    returns CompCurveToBSplineCurve;
    
    Add (me : in out; 
         NewCurve :  BoundedCurve from Geom2d;
         Tolerance:  Real from Standard;
         After      : Boolean from Standard = Standard_False)
	    ---Purpose: Append a curve in the BSpline
	    --          Return False if the curve is not G0 with the BSplineCurve.
	    --          Tolerance is used to check continuity and decrease 
	    --          Multiplicty at the common Knot 
	    --          After is usefull if BasisCurve is a closed curve .
    returns Boolean;
       
    
    Add (me : in out; 
         FirstCurve : in out BSplineCurve from Geom2d;
    	 SecondCurve: in out BSplineCurve from Geom2d;
         After      : Boolean from Standard)
	    ---Purpose: Concat two BSplineCurves.
    	is private;    
    
    BSplineCurve(me) returns BSplineCurve from Geom2d;

fields
 myCurve :  BSplineCurve from Geom2d;
 myTol   :  Real;
 myType  :  ParameterisationType from Convert;

end CompCurveToBSplineCurve;
