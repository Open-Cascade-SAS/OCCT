-- Created on: 1996-02-13
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class GIter from TopOpeBRepBuild

uses

    State from TopAbs,
    GTopo from TopOpeBRepBuild
    
is

    Create returns GIter;
    Create(G : GTopo) returns GIter;

    Find(me : in out) is static private;
    Init(me : in out) is static;
    Init(me : in out; G : GTopo) is static;
    More(me) returns Boolean is static;
    Next(me : in out) is static;
    Current(me; s1,s2 : in out State from TopAbs) is static;

    Dump(me; OS : in out OStream) is static;
    
fields

    myII : Integer;
    mypG : Address; -- (GTopo*)
    
end GIter;
