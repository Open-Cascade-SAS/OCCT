-- Created on: 1991-05-14
-- Created by: Laurent PAINNOT
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class FRPR from math
    	---Purpose:
    	-- this class implements the Fletcher-Reeves-Polak_Ribiere minimization 
    	-- algorithm of a function of multiple variables.
    	-- Knowledge of the function's gradient is required.

uses Vector from math, Matrix from math, 
     MultipleVarFunctionWithGradient from math,
     Status from math,
     OStream from Standard
     
raises DimensionError from Standard,
       NotDone from StdFail

is

    Create(theFunction: in MultipleVarFunctionWithGradient;
           theTolerance: Real;
           theNbIterations: Integer = 200;
           theZEPS: Real = 1.0e-12)
    ---Purpose:
    -- Initializes the computation of the minimum of F.
    -- Warning: constructor does not perform computations.
    returns FRPR;

    Delete(me) is static;
    ---Purpose: Destructor alias.
    ---C++: alias "  Standard_EXPORT virtual ~math_FRPR();"


    Perform(me: in out;
            theFunction: in out MultipleVarFunctionWithGradient; 
            theStartingPoint: Vector)
    ---Purpose:
    -- The solution F = Fi is found when
    -- 2.0 * abs(Fi - Fi-1) <= Tolerance * (abs(Fi) + abs(Fi-1) + ZEPS).
    is static;


    IsSolutionReached(me: in out; theFunction: in out MultipleVarFunctionWithGradient)
    ---Purpose:
    -- The solution F = Fi is found when:
    --   2.0 * abs(Fi - Fi-1) <= Tolerance * (abs(Fi) + abs(Fi-1)) + ZEPS.
    -- The maximum number of iterations allowed is given by NbIterations.
    ---C++:inline
    returns Boolean is virtual;


    IsDone(me)
        ---Purpose: Returns true if the computations are successful, otherwise returns false.
        ---C++: inline
    returns Boolean
    is static;
    
    

    Location(me)
    	---Purpose: returns the location vector of the minimum.
        -- Exception NotDone is raised if the minimum was not found.
        ---C++: inline
        ---C++: return const&
    
    returns Vector
    raises NotDone
    is static;


    Location(me; Loc: out Vector)
    	---Purpose: outputs the location vector of the minimum in Loc.
    	-- Exception NotDone is raised if the minimum was not found.
    	-- Exception DimensionError is raised if the range of Loc is not
    	-- equal to the range of the StartingPoint.
        ---C++: inline
    raises DimensionError,
    	   NotDone
    is static;
    

    Minimum(me)
       	---Purpose: returns the value of the minimum.
       	-- Exception NotDone is raised if the minimum was not found.
       	---C++: inline
    returns Real
    raises NotDone
    is static;
    
    
    Gradient(me)
       ---Purpose: returns the gradient vector at the minimum.
       -- Exception NotDone is raised if the minimum was not found.
       ---C++: inline
       ---C++: return const&
    returns Vector
    raises NotDone
    is static;
    
    
    Gradient(me; Grad: out Vector)
    	---Purpose: outputs the gradient vector at the minimum in Grad.
        -- Exception NotDone is raised if the minimum was not found.
        -- Exception DimensionError is raised if the range of Grad is not
        -- equal to the range of the StartingPoint.
        ---C++: inline
    
    raises DimensionError,
    	   NotDone
    is static;
    
    
    
    NbIterations(me)
	---Purpose: returns the number of iterations really done during the
        -- computation of the minimum.
        -- Exception NotDone is raised if the minimum was not found.
        ---C++: inline
    
    returns Integer
    raises NotDone
    is static;
    

    Dump(me; o: in out OStream)
	---Purpose: Prints on the stream o information on the current state 
    	--          of the object.
    	--          Is used to redefine the operator <<.

    is static;



fields

Done:            Boolean;
TheLocation:     Vector is protected;
TheGradient:     Vector is protected;
TheMinimum:      Real is protected;
PreviousMinimum: Real is protected;
Iter:            Integer;
State:           Integer;
XTol:            Real is protected;
EPSZ:            Real is protected;
TheStatus:       Status;
Itermax:         Integer;

end FRPR;
