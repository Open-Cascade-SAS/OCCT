-- Created on: 2002-12-12
-- Created by: data exchange team
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class FeaModel from StepFEA
inherits Representation from StepRepr

    ---Purpose: Representation of STEP entity FeaModel

uses
    HAsciiString from TCollection,
    HArray1OfRepresentationItem from StepRepr,
    RepresentationContext from StepRepr,
    HArray1OfAsciiString from TColStd

is
    Create returns FeaModel from StepFEA;
	---Purpose: Empty constructor

    Init (me: mutable; aRepresentation_Name: HAsciiString from TCollection;
                       aRepresentation_Items: HArray1OfRepresentationItem from StepRepr;
                       aRepresentation_ContextOfItems: RepresentationContext from StepRepr;
                       aCreatingSoftware: HAsciiString from TCollection;
                       aIntendedAnalysisCode: HArray1OfAsciiString from TColStd;
                       aDescription: HAsciiString from TCollection;
                       aAnalysisType: HAsciiString from TCollection);
	---Purpose: Initialize all fields (own and inherited)

    CreatingSoftware (me) returns HAsciiString from TCollection;
	---Purpose: Returns field CreatingSoftware
    SetCreatingSoftware (me: mutable; CreatingSoftware: HAsciiString from TCollection);
	---Purpose: Set field CreatingSoftware

    IntendedAnalysisCode (me) returns HArray1OfAsciiString from TColStd;
	---Purpose: Returns field IntendedAnalysisCode
    SetIntendedAnalysisCode (me: mutable; IntendedAnalysisCode: HArray1OfAsciiString from TColStd);
	---Purpose: Set field IntendedAnalysisCode

    Description (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Description
    SetDescription (me: mutable; Description: HAsciiString from TCollection);
	---Purpose: Set field Description

    AnalysisType (me) returns HAsciiString from TCollection;
	---Purpose: Returns field AnalysisType
    SetAnalysisType (me: mutable; AnalysisType: HAsciiString from TCollection);
	---Purpose: Set field AnalysisType

fields
    theCreatingSoftware: HAsciiString from TCollection;
    theIntendedAnalysisCode: HArray1OfAsciiString from TColStd;
    theDescription: HAsciiString from TCollection;
    theAnalysisType: HAsciiString from TCollection;

end FeaModel;
