-- Created on: 1995-07-24
-- Created by: Modelistation
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class PoleCurve from StdPrs 

inherits Root from Prs3d
     
  	     
    	---Purpose: A framework to provide display of Bezier or BSpline curves.

uses
    Curve        from Adaptor3d,
    Presentation from Prs3d,
    Drawer       from Prs3d,
    Length       from Quantity 

is

    --- Purpose:
    
    Add(myclass; aPresentation: Presentation from Prs3d; 
    	    	 aCurve       : Curve        from Adaptor3d;
    	    	 aDrawer      : Drawer       from Prs3d);
    	---Purpose: Defines display of BSpline and Bezier curves.
    	-- Adds the 3D curve aCurve to the
    	-- StdPrs_PoleCurve algorithm. This shape is found in
    	-- the presentation object aPresentation, and its display
    	-- attributes are set in the attribute manager aDrawer.
    	-- The curve object from Adaptor3d provides data from
    	-- a Geom curve. This makes it possible to use the
    	-- surface in a geometric algorithm.

		 
    Match(myclass; X,Y,Z    : Length from Quantity;
                   aDistance: Length from Quantity;
    	    	   aCurve   : Curve  from Adaptor3d;
    	    	   aDrawer  : Drawer from Prs3d) 
    returns Boolean from Standard;
    	---Purpose: returns true if the distance between the point (X,Y,Z) and the
    	--          broken line made of the poles is less then aDistance.


    Pick(myclass; X,Y,Z    : Length from Quantity;
    	          aDistance: Length from Quantity;
                  aCurve   : Curve  from Adaptor3d;
    	          aDrawer  : Drawer from Prs3d)
    returns Integer from Standard;
    	---Purpose: returns the pole  the most near of the point (X,Y,Z) and
    	--          returns its range. The distance between the pole and
    	--          (X,Y,Z) must be less then aDistance. If no pole corresponds, 0 is returned.

end PoleCurve from StdPrs;



