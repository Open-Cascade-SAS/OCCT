-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class BSplineSurfaceWithKnots from StepGeom 

inherits BSplineSurface from StepGeom 

uses

	HArray1OfInteger from TColStd, 
	HArray1OfReal from TColStd, 
	KnotType from StepGeom, 
	Integer from Standard, 
	Real from Standard, 
	HAsciiString from TCollection, 
	HArray2OfCartesianPoint from StepGeom, 
	BSplineSurfaceForm from StepGeom, 
	Logical from StepData
is

	Create returns BSplineSurfaceWithKnots;
	---Purpose: Returns a BSplineSurfaceWithKnots


	Init (me : mutable;
	      aName : HAsciiString from TCollection;
	      aUDegree : Integer from Standard;
	      aVDegree : Integer from Standard;
	      aControlPointsList : HArray2OfCartesianPoint from StepGeom;
	      aSurfaceForm : BSplineSurfaceForm from StepGeom;
	      aUClosed : Logical from StepData;
	      aVClosed : Logical from StepData;
	      aSelfIntersect : Logical from StepData) is redefined;

	Init (me : mutable;
	      aName : HAsciiString from TCollection;
	      aUDegree : Integer from Standard;
	      aVDegree : Integer from Standard;
	      aControlPointsList : HArray2OfCartesianPoint from StepGeom;
	      aSurfaceForm : BSplineSurfaceForm from StepGeom;
	      aUClosed : Logical from StepData;
	      aVClosed : Logical from StepData;
	      aSelfIntersect : Logical from StepData;
	      aUMultiplicities : HArray1OfInteger from TColStd;
	      aVMultiplicities : HArray1OfInteger from TColStd;
	      aUKnots : HArray1OfReal from TColStd;
	      aVKnots : HArray1OfReal from TColStd;
	      aKnotSpec : KnotType from StepGeom) is virtual;

	-- Specific Methods for Field Data Access --

	SetUMultiplicities(me : mutable; aUMultiplicities : HArray1OfInteger);
	UMultiplicities (me) returns HArray1OfInteger;
	UMultiplicitiesValue (me; num : Integer) returns Integer;
	NbUMultiplicities (me) returns Integer;
	SetVMultiplicities(me : mutable; aVMultiplicities : HArray1OfInteger);
	VMultiplicities (me) returns HArray1OfInteger;
	VMultiplicitiesValue (me; num : Integer) returns Integer;
	NbVMultiplicities (me) returns Integer;
	SetUKnots(me : mutable; aUKnots : HArray1OfReal);
	UKnots (me) returns HArray1OfReal;
	UKnotsValue (me; num : Integer) returns Real;
	NbUKnots (me) returns Integer;
	SetVKnots(me : mutable; aVKnots : HArray1OfReal);
	VKnots (me) returns HArray1OfReal;
	VKnotsValue (me; num : Integer) returns Real;
	NbVKnots (me) returns Integer;
	SetKnotSpec(me : mutable; aKnotSpec : KnotType);
	KnotSpec (me) returns KnotType;

fields

	uMultiplicities : HArray1OfInteger from TColStd;
	vMultiplicities : HArray1OfInteger from TColStd;
	uKnots : HArray1OfReal from TColStd;
	vKnots : HArray1OfReal from TColStd;
	knotSpec : KnotType from StepGeom; -- an Enumeration

end BSplineSurfaceWithKnots;
