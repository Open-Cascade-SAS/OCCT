-- Created on: 1996-03-15
-- Created by: Christian CAILLET
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ModifReorder  from IFSelect  inherits Modifier

    ---Purpose : This modifier reorders a whole model from its roots, i.e.
    --           according to <rootlast> status, it considers each of its
    --           roots, then it orders all its shared entities at any level,
    --           the result begins by the lower level entities ... ends by
    --           the roots.

uses CString, AsciiString from TCollection,
     InterfaceModel, CopyTool, Protocol from Interface, ContextModif

is

    Create (rootlast : Boolean = Standard_True) returns mutable ModifReorder;
    ---Purpose : Creates a ModifReorder. It may change the graph (it does !)
    --           If <rootlast> is True (D), roots are set at the end of packets
    --           Else, they are set at beginning (as done by AddWithRefs)

    Perform (me; ctx  : in out ContextModif;
    	     target   : mutable InterfaceModel;
    	     protocol : Protocol from Interface;
    	     TC       : in out CopyTool);
    ---Purpose : Acts by computing orders (by method All from ShareTool) then
    --           forcing them in the model. Remark that selection is ignored :
    --           ALL the model is processed in once

    Label (me) returns AsciiString from TCollection;
    ---Purpose : Returns Label as "Reorder, Roots (last or first)"

fields

    thertl : Boolean;

end ModifReorder;
