-- Created on: 1992-04-13
-- Created by: Isabelle GRIGNON
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



package IntImp

	---Purpose: 

uses Standard, TColStd, StdFail, math, gp, IntSurf

is

    enumeration ConstIsoparametric is
                UIsoparametricOnCaro1, VIsoparametricOnCaro1,
                UIsoparametricOnCaro2, VIsoparametricOnCaro2;
		
    deferred generic class PSurfaceTool;

    deferred generic class ISurfaceTool;

    deferred generic class CurveTool;

    deferred generic class CSCurveTool;

    deferred generic class COnSCurveTool;

    generic class ZerImpFunc; -- inherits FunctionSetWithDerivatives
    
    generic class ZerParFunc; -- inherits FunctionSetWithDerivatives

    deferred generic class CSFunction; -- inherits FunctionSetWithDerivatives

    generic class ZerCSParFunc; -- inherits FunctionSetWithDerivatives
    
    generic class ZerCOnSSParFunc; -- inherits FunctionSetWithDerivatives
    
    generic class Int2S,TheFunction;
    
    generic class IntCS;

end IntImp;
