-- File:	StepBasic_NameAssignment.cdl
-- Created:	Wed May 10 15:09:08 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class NameAssignment from StepBasic
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity NameAssignment

uses
    HAsciiString from TCollection

is
    Create returns NameAssignment from StepBasic;
	---Purpose: Empty constructor

    Init (me: mutable; aAssignedName: HAsciiString from TCollection);
	---Purpose: Initialize all fields (own and inherited)

    AssignedName (me) returns HAsciiString from TCollection;
	---Purpose: Returns field AssignedName
    SetAssignedName (me: mutable; AssignedName: HAsciiString from TCollection);
	---Purpose: Set field AssignedName

fields
    theAssignedName: HAsciiString from TCollection;

end NameAssignment;
