-- File:	Dynamic_StringParameter.cdl
-- Created:	Wed Feb  3 15:49:43 1993
-- Author:	Gilles DEBARBOUILLE
--		<gde@bravox>
---Copyright:	 Matra Datavision 1993



class StringParameter from Dynamic

inherits

    Parameter from Dynamic


	---Purpose: This inherited class  from Parameter describes all
	--          the  parameters,  which   are  characterized by  a
	--          string value.

uses

    OStream from Standard,
    CString from Standard,
    HAsciiString from TCollection,
    AsciiString  from TCollection

is

    Create(aparameter : CString from Standard )
    
    ---Level: Public 
    
    ---Purpose: Creates a StringParameter with <aparameter> as name.
    
    returns mutable StringParameter from Dynamic;

    Create(aparameter : CString from Standard ; astring : CString from Standard) 
    
    ---Level: Public 
    
    ---Purpose: With  the name of  the  Parameter <aparameter> and the
    --          string    <astring>,   creates    an    instance    of
    --          StringParameter.
    
    returns mutable StringParameter from Dynamic;
    
    Value(me) returns AsciiString from TCollection
    
    ---Level: Public 
    
    ---Purpose: Returns the value    of  the parameter which     is an
    --          AsciiString.
    
    is static;

    Value (me : mutable ; avalue : CString from Standard)
    
    ---Level: Public 
    
    --- Purpose: Sets the string <avalue> in <me>.

    is static;
    
    Dump(me ; astream : in out OStream from Standard)
    
    ---Level: Internal 
    
    ---Purpose: Useful for debugging.

    is redefined;

fields

    thestring : HAsciiString from TCollection;

end StringParameter;
