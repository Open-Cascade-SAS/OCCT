-- Created on: 1996-02-15
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class FindEdges from LocOpe

	---Purpose: 

uses Shape                      from TopoDS,
     Edge                      from TopoDS,
     ListOfShape               from TopTools,
     ListIteratorOfListOfShape from TopTools
     

raises ConstructionError from Standard,
       NoSuchObject      from Standard,
       NoMoreObject      from Standard

is

    Create
    	returns FindEdges from LocOpe;
	---C++: inline



    Create(FFrom,FTo: Shape from TopoDS)
    
	---C++: inline
    	returns FindEdges from LocOpe
	raises ConstructionError from Standard;
	
	
    Set(me: in out; FFrom, FTo: Shape from TopoDS)
    
	raises ConstructionError from Standard
    	is static;


    InitIterator(me: in out)
    
	---C++: inline
    	is static;


    More(me)
    
    	returns Boolean from Standard
	---C++: inline
	is static;


    EdgeFrom(me)
    
    	returns Edge from TopoDS
	---C++: return const&
	---C++: inline
	raises NoSuchObject from Standard
	is static;


    EdgeTo(me)
    
    	returns Edge from TopoDS
	---C++: return const&
	---C++: inline
	raises NoSuchObject from Standard
	is static;


    Next(me: in out)
    
	---C++: inline
    	raises NoMoreObject from Standard
	is static;


fields

    myFFrom  : Shape                     from TopoDS;
    myFTo    : Shape                     from TopoDS;
    myLFrom  : ListOfShape               from TopTools;
    myLTo    : ListOfShape               from TopTools;
    myItFrom : ListIteratorOfListOfShape from TopTools;
    myItTo   : ListIteratorOfListOfShape from TopTools;

end FindEdges;
