-- File:	QABRGM.cdl
-- Created:	Wed Mar 20 17:10:09 2002
-- Author:	QA Admin
--		<qa@umnox.nnov.matra-dtv.fr>
---Copyright:	 Matra Datavision 2002

package QABRGM
     uses Draw
is
    Commands(DI : in out Interpretor from Draw);
end;
    
