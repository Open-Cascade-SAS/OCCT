-- Created on: 1992-11-17
-- Created by: Christian CAILLET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SelectModelEntities  from IFSelect  inherits SelectBase

    ---Purpose : A SelectModelEntities gets all the Entities of an
    --           InterfaceModel.

uses AsciiString from TCollection, EntityIterator, Graph

is

    Create  returns SelectModelEntities;
    ---Purpose : Creates a SelectModelRoot

    RootResult (me; G : Graph) returns EntityIterator;
    ---Purpose : Returns the list of selected entities : the Entities of the
    --           Model (note that this result assures naturally uniqueness)

    CompleteResult (me; G : Graph) returns EntityIterator  is redefined;
    ---Purpose : The complete list of Entities (including shared ones) ...
    --           is exactly identical to RootResults in this case

    Label (me) returns AsciiString from TCollection;
    ---Purpose : Returns a text defining the criterium : "Model Entities"

end SelectModelEntities;
