-- File:	RWStepRepr_RWCompositeShapeAspect.cdl
-- Created:	Wed Jun  4 14:17:23 2003 
-- Author:	Galina KULIKOVA
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWCompositeShapeAspect from RWStepRepr

    ---Purpose: Read & Write tool for CompositeShapeAspect

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    CompositeShapeAspect from StepRepr

is
    Create returns RWCompositeShapeAspect from RWStepRepr;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : CompositeShapeAspect from StepRepr);
	---Purpose: Reads CompositeShapeAspect

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: CompositeShapeAspect from StepRepr);
	---Purpose: Writes CompositeShapeAspect

    Share (me; ent : CompositeShapeAspect from StepRepr;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWCompositeShapeAspect;
