-- Created on: 1992-06-22
-- Created by: Gilles DEBARBOUILLE
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class MethodDefinitionsDictionary from Dynamic

inherits

    Transient
    
	---Purpose: This  class groups  in   a dictionary  of  all the
	--          various definitions of methods. It also allows the
	--          share of  the  same  definition by  more  than one
	--          MethodInstance to  preserve a global coherence and
	--          also to  manage the memory.   To use this class an
	--          inheritance is necessary with perhaps the overload
	--          of the Switch   method if the parameter  types are
	--          not      of     the      type    BooleanParameter,
	--          IntegerParameter,       RealParameter          and
	--          StringParameter.

uses

    CString from Standard,
    OStream from Standard,
    Boolean from Standard,
    Integer from Standard,
    HAsciiString                from TCollection,
    Parameter                   from Dynamic,
    SequenceOfMethodDefinitions from Dynamic,
    Method                      from Dynamic

is

    Initialize;
    
    ---Level: Internal 
    
    ---Purpose: Deferred constructor of the class.
    
    Creates(me : mutable ; afilename : CString from Standard)
    
    ---Level: Internal 
    
    ---Purpose: Starting with   a file named  <afilename>,  fills  the
    --          dictionary with all the wishes definitions.
    
    is static;
    
    Definition(me : mutable ; adefinition : Method from Dynamic) returns Boolean from Standard
    
    ---Level: Advanced 
    
    ---Purpose: This method sets  the new definition  <adefinition> in
    --          the dictionary. It   returns true if the operation  is
    --          successful, false otherwise.
    
    is static;
    
    Switch(me ; aname , atype , avalue : CString from Standard)
    
    ---Level: Internal 
    
    ---Purpose: This virtual method allows the user to add recognition
    --          of its  own  parameters when reading  the file to fill
    --          the dictionary.
    
    returns Parameter from Dynamic;
    
    Definition(me ; atype       : CString from Standard
                  ; adefinition : out Method from Dynamic) returns Boolean from Standard
        
    ---Level: Public 
    
    ---Purpose: Returns from     the dictionary in  the   out variable
    --          <adefinition> a reference to the right instance of the
    --          definition identified  by its type <atype>. The method
    --          returns true if the definition exist, false otherwise.
    
    is static;
    
    UpToDate(me) returns Boolean from Standard
    
    ---Level: Advanced 
    
    ---Purpose: Returns true if there has  been no modification of the
    --          file  method-definitions.dat since the creation of the
    --          dictionary object, false otherwise.
    
    is static;
    
    NumberOfDefinitions(me) returns Integer from Standard
    
    ---Level: Public 
    
    ---Purpose: Returns    the number  of  definitions  stored  in the
    --          dictionary.
    
    is static;
    
    Definition(me ; anindex : Integer from Standard) returns any Method from Dynamic
    
    ---Level: Public 
    
    ---Purpose: Returns a  reference on the  definition identified  by
    --          the index <anidex>.
    
    is static;
    
    Dump(me ; astream : in out OStream from Standard)
    
    ---Level: Internal 
    
    ---Purpose: Useful for debugging.
    
    is static;

fields

    thefilename                    : HAsciiString                from TCollection;
    thetime                        : Time                        from Standard;
    thesequenceofmethoddefinitions : SequenceOfMethodDefinitions from Dynamic;

end MethodDefinitionsDictionary;
