-- Created on: 1992-02-17
-- Created by: Christian CAILLET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class BinderOfShape from TransferBRep inherits Binder from Transfer

    ---Purpose : Allows direct binding between a starting Object and the Result
    --           of its transfer when it is Unique.
    --           The Result itself is defined as a formal parameter <Shape from TopoDS>           
    --  Warning : While it is possible to instantiate BinderOfShape with any Type
    --           for the Result, it is not advisable to instantiate it with
    --           Transient Classes, because such Results are directly known and
    --           managed by TransferProcess & Co, through
    --           SimpleBinderOfTransient : this class looks like instantiation
    --           of BinderOfShape, but its method ResultType
    --           is adapted (reads DynamicType of the Result)

uses CString,
     Type,
     Shape     from TopoDS,
     ShapeInfo from TransferBRep

raises TransferFailure

is

    Create returns mutable BinderOfShape;
    ---Purpose : normal standard constructor, creates an empty BinderOfShape

    Create (res : any Shape from TopoDS) returns mutable BinderOfShape;
    ---Purpose : constructor which in the same time defines the result

--    IsMultiple (me) returns Boolean;
    ---Purpose : Returns True if a starting object is bound with SEVERAL
    --           results : Here, returns allways False
    --           But it can have next results

    ResultType (me) returns Type;
    ---Purpose : Returns the Type permitted for the Result, i.e. the Type
    --           of the Parameter Class <Shape from TopoDS> (statically defined)

    ResultTypeName (me) returns CString;
    ---Purpose : Returns the Type Name computed for the Result (dynamic)

    SetResult (me : mutable; res : any Shape from TopoDS)
    ---Purpose : Defines the Result
    	raises TransferFailure;
    --           Error if the Result is already used (see class Binder)

    Result (me) returns any Shape from TopoDS
    ---Purpose : Returns the defined Result, if there is one
    	raises TransferFailure;
    --           Error if the Result is not defined (see class Binder)
    ---C++ : return const &

    CResult (me : mutable) returns any Shape from TopoDS;
    ---Purpose : Returns the defined Result, if there is one, and allows to
    --           change it (avoids Result + SetResult).
    --           Admits that Result can be not yet defined
    --  Warning : a call to CResult causes Result to be known as defined
    ---C++ : return &

fields

    theres : Shape from TopoDS;

end BinderOfShape;
