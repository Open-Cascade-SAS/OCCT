-- Created on: 1992-09-01
-- Created by: Remi GILET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MakeMirror2d

from gce

    ---Purpose: This class implements elementary construction algorithms for a
    -- symmetrical transformation in 2D space about a point
    -- or axis. The result is a gp_Trsf2d transformation.
    -- A MakeMirror2d object provides a framework for:
    -- -   defining the construction of the transformation,
    -- -   implementing the construction algorithm, and consulting the result.

uses Pnt2d  from gp,
     Ax2d   from gp,
     Dir2d  from gp,
     Lin2d  from gp,
     Trsf2d from gp,
     Real   from Standard
     
is

Create(Point : Pnt2d from gp) returns MakeMirror2d;
    ---Puprose: Makes a symmetry transformation of center <Point>.

Create(Axis : Ax2d from gp) returns MakeMirror2d;
    ---Puprose: Makes a symmetry transformation of axis <Axis>.

Create(Line : Lin2d from gp) returns MakeMirror2d;
    ---Puprose: Makes a symmetry transformation of axis <Line>.

Create(Point : Pnt2d from gp;
       Direc : Dir2d from gp) returns MakeMirror2d;
    ---Purpose: Makes a symmetry transformation af axis defined by 
    --          <Point> and <Direc>.

Value(me) returns Trsf2d from gp
    is static;
    ---C++: return const&
    ---Purpose: Returns the constructed transformation.

Operator(me) returns Trsf2d from gp
    is static;
    ---C++: return const&
    ---C++: alias "Standard_EXPORT operator gp_Trsf2d() const;"

fields

    TheMirror2d : Trsf2d from gp;

end MakeMirror2d;

