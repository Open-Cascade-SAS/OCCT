-- Created on: 1992-11-17
-- Created by: Remi LEQUETTE
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred generic class Intersection2d from TopClass 
    (TheEdge as any) inherits Intersection from IntRes2d 

	---Purpose: Template  class for  the  intersection   algorithm
	--          required by the 2D classifications.
	--          
	--          The results should be  expressed as the  result of
	--          Intersection   from IntRes2d.   The class used  to
	--          instantiate the Classifier2d can be inherited from
	--          the    Intersection  algorithms   inherited   from
	--          Intersection from IntRes2d.
	--          
	--          It is not necesary to return  all the Intersection
	--          points, the  point with   the   smallest parameter
	--          value on the segment is enough.

uses
    Lin2d from gp,
    Dir2d from gp

is
    Initialize;
	---Purpose: An empty constructor is required.
	
    Perform(me : in out; L : Lin2d from gp; P : Real; Tol : Real; E : TheEdge)
	---Purpose: Performs the intersection   between the  2d   line
	--          segment (<L>, <P>) and  the  Edge <E>.   The  line
	--          segment  is the  part  of  the  2d   line   <L> of
	--          parameter range [0, <P>] (P is positive and can be
	--          RealLast()). Tol is the  Tolerance on the segment.
	--          The order  is relevant, the  first argument is the
	--          segment, the second the Edge.
    is deferred;
	
    LocalGeometry(me; E : TheEdge;  U : Real; 
    	    	      T : out Dir2d from gp; 
    	    	      N : out Dir2d from gp;
                      C : out Real)
	---Purpose: Returns in <T>,  <N> and <C>  the tangent,  normal
	--          and  curvature of the edge  <E> at parameter value
	--          <U>.
    is deferred;

end Intersection2d;
