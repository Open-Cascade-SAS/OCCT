-- Created on: 1992-02-20
-- Created by: Remy GILET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



generic class FunctionTanCuCu from GccIter (
    TheCurve     as any;
    TheCurveTool as any) -- as CurvePGTool from GccInt (TheCurve)

inherits FunctionSetWithDerivatives from math 

    ---Purpose: This abstract class describes a Function of 1 Variable 
    --          used to find a line tangent to two curves.

uses Vector from math,
     Matrix from math,
     Circ2d from gp,
     Pnt2d  from gp,
     Vec2d  from gp,
     Type3  from GccIter

     
raises ConstructionError

is

Create (Curv1 : TheCurve ;
        Curv2 : TheCurve ) returns FunctionTanCuCu from GccIter;

Create (Circ1 : Circ2d   from gp ;
        Curv2 : TheCurve         ) returns FunctionTanCuCu from GccIter;

InitDerivative(me                   : in out                      ;
    	       X                    :        Vector from math     ;
	       Point1,Point2        :    out Pnt2d  from gp       ;
	       Tan1,Tan2,D21,D22    :    out Vec2d  from gp       )
raises ConstructionError
is static;

NbVariables(me) returns Integer;
    ---Purpose: returns the number of variables of the function.

NbEquations(me) returns Integer;
    ---Purpose: returns the number of equations of the function.

Value (me : in out                 ;
       X  :        Vector from math;
       F  :    out Vector from math) returns Boolean;
    ---Purpose: Computes the value of the function F for the variable X.
    --          It returns True if the computation is successfully done,
    --          False otherwise.

Derivatives (me    : in out                 ;
             X     :        Vector from math;
             Deriv :    out Matrix from math) returns Boolean;
    ---Purpose: Computes the derivative of the function F for the variable X.
    --          It returns True if the computation is successfully done,
    --          False otherwise.

Values (me    : in out                 ;
        X     :        Vector from math;
        F     : out    Vector from math;
        Deriv : out    Matrix from math) returns Boolean;
    ---Purpose: Computes the value and the derivative of the function F 
    --          for the variable X.
    --          It returns True if the computation is successfully done,
    --          False otherwise.

fields

TheCurve1     : TheCurve               ;
TheCurve2     : TheCurve               ;
TheCirc1      : Circ2d   from gp       ;
TheType       : Type3    from GccIter  ;

end FunctionTanCuCu;



