-- File:	IGESBasic_ToolSubfigureDef.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolSubfigureDef  from IGESBasic

    ---Purpose : Tool to work on a SubfigureDef. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses SubfigureDef from IGESBasic,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolSubfigureDef;
    ---Purpose : Returns a ToolSubfigureDef, ready to work


    ReadOwnParams (me; ent : mutable SubfigureDef;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : SubfigureDef;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : SubfigureDef;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a SubfigureDef <ent>, from
    --           its specific (own) parameters

    DirChecker (me; ent : SubfigureDef) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : SubfigureDef;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : SubfigureDef; entto : mutable SubfigureDef;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : SubfigureDef;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolSubfigureDef;
