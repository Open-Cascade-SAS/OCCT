-- File:	StepToGeom_MakeSurfaceOfRevolution.cdl
-- Created:	Mon Jun 14 16:20:58 1993
-- Author:	Martine LANGLOIS
---Copyright:	 Matra Datavision 1993

class MakeSurfaceOfRevolution from StepToGeom

    ---Purpose: This class implements the mapping between class
    --          SurfaceOfRevolution from StepGeom which describes a
    --          surface_of_revolution from Prostep and SurfaceOfRevolution
    --          from Geom 

uses SurfaceOfRevolution from Geom,
     SurfaceOfRevolution from StepGeom

is 

    Convert ( myclass; SS : SurfaceOfRevolution from StepGeom;
                       CS : out SurfaceOfRevolution from Geom )
    returns Boolean from Standard;

end MakeSurfaceOfRevolution;
