-- Created on: 2008-07-02
-- Created by: Alexander GRIGORIEV
-- Copyright (c) 2008-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Dummy package header

package NIS
uses
     V3d,
     Bnd
is
    imported Drawer;
    imported DrawList;
    imported InteractiveContext;
    imported InteractiveObject;
    imported ObjectsIterator;
    imported SelectFilter;
    imported Surface;
    imported SurfaceDrawer;
    imported Triangulated;
    imported TriangulatedDrawer;
    imported View;
    
end NIS;
