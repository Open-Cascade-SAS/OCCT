-- Created on: 1993-07-08
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class BoxSort from TopOpeBRepTool

uses

    Box from Bnd,
    BoundSortBox from Bnd,
    HArray1OfBox from Bnd,
    HArray1OfInteger from TColStd,
    ListOfInteger from TColStd,
    ListIteratorOfListOfInteger from TColStd,
    ShapeEnum from TopAbs,
    Shape from TopoDS,
    IndexedMapOfShape from TopTools,
    Box from Bnd,
    HBoxTool from TopOpeBRepTool
    
is

    Create returns BoxSort;
    Create(T:HBoxTool) returns BoxSort;
    SetHBoxTool(me:in out;T:HBoxTool);
    HBoxTool(me) returns HBoxTool;---C++: return const &
    Clear(me:in out);
    AddBoxes(me:in out;S:Shape;TS:ShapeEnum;TA:ShapeEnum=TopAbs_SHAPE);
    MakeHAB(me:in out;S:Shape;TS:ShapeEnum;TA:ShapeEnum=TopAbs_SHAPE);
    HAB(me) returns HArray1OfBox from Bnd;---C++:return const &
    MakeHABCOB(myclass;HAB:HArray1OfBox from Bnd;COB:out Box from Bnd);
    HABShape(me; I:Integer) returns Shape;---C++: return const &
    MakeCOB(me:in out;S:Shape;TS:ShapeEnum;TA:ShapeEnum=TopAbs_SHAPE);
    AddBoxesMakeCOB(me:in out;S:Shape;TS:ShapeEnum;TA:ShapeEnum=TopAbs_SHAPE);
    Compare(me:out;S:Shape) returns ListIteratorOfListOfInteger;---C++:return const&
    TouchedShape(me;I:ListIteratorOfListOfInteger) returns Shape;---C++:return const&
    Box(me;S:Shape) returns Box from Bnd;---C++:return const & 
    
--modified by NIZNHY-PKV Mon Dec 16 10:24:42 2002  f
    Destroy(me: out); 
    ---C++:  alias  "Standard_EXPORT ~TopOpeBRepTool_BoxSort() {Destroy();}"
--modified by NIZNHY-PKV Mon Dec 16 10:25:22 2002  t

fields

    myCOB:Box from Bnd;
    myBSB:BoundSortBox from Bnd;
    myIterator:ListIteratorOfListOfInteger from TColStd;
    myLastCompareShape:Shape from TopoDS;
    myLastCompareShapeBox:Box from Bnd;
    myHBT:HBoxTool from TopOpeBRepTool;
    myHAB:HArray1OfBox from Bnd;
    myHAI:HArray1OfInteger from TColStd;    

end BoxSort;
