-- Created on: 1993-07-21
-- Created by: Martine LANGLOIS
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


private deferred class Root from TopoDSToStep

    ---Purpose : This class implements the common services for
    --           all classes of TopoDSToStep which report error.

uses Real

is

    Initialize;

    Tolerance (me : in out) returns Real;
    ---Purpose : Returns (modifiable) the tolerance to be used for writing
    --           If not set, starts at 0.0001
    ---C++ : return &

    IsDone(me) returns Boolean
    	is static;

fields

    toler    : Real    is protected;
    done     : Boolean is protected;
    --Equal True if everything is ok, False otherwise.

end Root;
