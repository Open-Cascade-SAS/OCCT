-- Created on: 1993-01-28
-- Created by: Gilles DEBARBOUILLE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class InterpretedMethod from Dynamic

inherits

    MethodDefinition from Dynamic

	---Purpose: This class derived from Method, describes an  
	--          interpreted method. The additional field is the 
	--          name of the file to be interpreted.

uses

    CString from Standard,
    HAsciiString from TCollection,
    AsciiString  from TCollection

is

    Create(aname , afile : CString from Standard) returns mutable InterpretedMethod from Dynamic;
    
    ---Level: Public 
    
    ---Purpose: Creates a new  InterpretedMethod with <aname> as  name
    --          and <afile> as file name to be interpreted.
    
    Function(me : mutable ; afile : CString from Standard)
    
    ---Level: Public 
    
    ---Purpose: Sets the the   name of the  file to  be interpreted to
    --          <afile>.
    
    is static;
    
    Function(me) returns AsciiString from TCollection
    
    ---Level: Public 
    
    ---Purpose: Returns the name of the file to be interpreted.
    
    is static;
    
fields

    thefunction : HAsciiString from TCollection;

end InterpretedMethod;
