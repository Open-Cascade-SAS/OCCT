-- Created on: 1996-12-05
-- Created by: Odile Olivier
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DimensionOwner from AIS inherits EntityOwner from SelectMgr

  ---Purpose: The owner is the entity which makes it possible to link
    -- the sensitive primitives and the reference shapes that
    -- you want to detect. It stocks the various pieces of
    -- information which make it possible to find objects. An
    -- owner has a priority which you can modulate, so as to
    -- make one entity more selectable than another. You
    -- might want to make edges more selectable than
    -- faces, for example. In that case, you could attribute sa
    -- higher priority to the one compared to the other. An
    -- edge, could have priority 5, for example, and a face,
    -- priority 4. The default priority is 5.

uses

    SelectableObject       from SelectMgr,
    PresentationManager    from PrsMgr,
    PresentationManager3d  from PrsMgr,
    NameOfColor            from Quantity,
    DimensionSelectionMode from AIS

is

    Create (theSelObject  : SelectableObject;
            theSelMode    : DimensionSelectionMode from AIS;
            thePriority   : Integer from Standard = 0)
    returns DimensionOwner from AIS;
      ---Purpose:
      -- Initializes the dimension owner, theSO, and attributes it
      -- the priority, thePriority.

    SelectionMode (me)
    returns DimensionSelectionMode from AIS;

    HilightWithColor (me       : mutable;
                      thePM    : PresentationManager3d from PrsMgr;
                      theColor : NameOfColor from Quantity;
                      theMode  : Integer  from  Standard = 0)
    is redefined virtual;

    IsHilighted (me;
                 thePM   : PresentationManager from PrsMgr;
                 theMode : Integer  from  Standard  =0)
    returns Boolean from Standard is redefined virtual;
    ---Purpose: Returns true if an object with the selection mode
    -- aMode is highlighted in the presentation manager aPM.

    Hilight(me    : mutable;
            thePM   : PresentationManager from PrsMgr;
            theMode : Integer  from  Standard  =0) is redefined virtual;

    Unhilight(me    : mutable;
              thePM   : PresentationManager from PrsMgr;
              theMode : Integer  from  Standard  =0) is redefined virtual;
    ---Purpose: Removes highlighting from the selected part of dimension.

fields

    mySelectionMode : DimensionSelectionMode from AIS;

end DimensionOwner;
