-- File:	Segment3D.cdl
-- Created:	Thu Apr 25 10:27:04 1991
-- Author:	Arnaud BOUZY
--		<adn@topsn2>
---Copyright:	 Matra Datavision 1991


class Segment3D from Draw inherits Drawable3D from Draw

	---Purpose: 

uses Pnt from gp,
    Color from Draw,
    Display from Draw

is

    Create(p1,p2 : Pnt; col : Color)
    returns mutable Segment3D;
    
    DrawOn(me; dis : in out Display);
    
    First(me) returns Pnt from gp
	---C++: return const&
    is static;

    First(me : mutable; P : Pnt from gp)
    is static;

    Last(me) returns Pnt from gp
	---C++: return const&
    is static;

    Last(me : mutable; P : Pnt from gp)
    is static;

fields

    myFirst : Pnt;
    myLast  : Pnt;
    myColor : Color;
    
end Segment3D;
