-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class TextOrCharacter from StepVisual inherits SelectType from StepData

	-- <TextOrCharacter> is an EXPRESS Select Type construct translation.
	-- it gathers : AnnotationText, CompositeText, TextLiteral

uses

	AnnotationText,
	CompositeText,
	TextLiteral
is

	Create returns TextOrCharacter;
	---Purpose : Returns a TextOrCharacter SelectType

	CaseNum (me; ent : Transient) returns Integer;
	---Purpose: Recognizes a TextOrCharacter Kind Entity that is :
	--        1 -> AnnotationText
	--        2 -> CompositeText
	--        3 -> TextLiteral
	--        0 else

	AnnotationText (me) returns any AnnotationText;
	---Purpose : returns Value as a AnnotationText (Null if another type)

	CompositeText (me) returns any CompositeText;
	---Purpose : returns Value as a CompositeText (Null if another type)

	TextLiteral (me) returns any TextLiteral;
	---Purpose : returns Value as a TextLiteral (Null if another type)


end TextOrCharacter;

