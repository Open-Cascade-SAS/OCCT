-- Created on: 1995-04-24
-- Created by: Modelistation
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class FilSpine from ChFiDS inherits Spine from ChFiDS 

	---Purpose: Provides  data specific to  the fillets -
	--          vector or rule  of evolution (C2).
	--          


uses
    HArray1OfReal from TColStd,  
    HElSpine      from ChFiDS,
    Function      from Law,
    Laws          from Law,
    Composite     from Law,
    Edge          from TopoDS,
    Vertex        from TopoDS,
    SequenceOfXY  from TColgp, 
    XY	          from gp

is

    Create  returns FilSpine from ChFiDS;

    Create(Tol : Real from Standard) returns FilSpine from ChFiDS;

    Reset(me : mutable; AllData : Boolean from Standard = Standard_False)
    is redefined;

    ------------------------------------------------
    -- Update selectif du rayon par edges ou vertex.
    ------------------------------------------------

    SetRadius(me     : mutable;
    	      Radius : Real from Standard;
              E      : Edge from TopoDS) 
    ---Purpose: initializes the constant vector on edge E.
    is static;

    UnSetRadius(me     : mutable;
                E      : Edge from TopoDS) 
    ---Purpose: resets the constant vector  on   edge E.
    is static;

    SetRadius(me     : mutable;
    	      Radius : Real from Standard;
              V      : Vertex from TopoDS) 
    ---Purpose: initializes the  vector on Vertex V.
    is static;

    UnSetRadius(me     : mutable;
                V      : Vertex from TopoDS) 
    ---Purpose: resets the vector on Vertex V.
    is static;

    SetRadius(me     : mutable;
    	      UandR  : XY from gp;
              IinC   : Integer from Standard) 
    ---Purpose: initializes the vector on the point of parameter W.
    is static;

    SetRadius(me : mutable;Radius : Real from Standard) 
    ---Purpose: initializes the constant vector on all spine.
    is static;
    
    SetRadius(me : mutable; 
    	      C      : Function from Law;
              IinC   : Integer from Standard) 
    ---Purpose: initializes the rule of evolution on all spine.
    is static;
    
    IsConstant(me) 
    returns Boolean from Standard
    ---Purpose: returns true if the radius is constant 
    --          all along the spine.
    is static;
    
    IsConstant(me; IE : Integer from Standard) 
    returns Boolean from Standard
    ---Purpose: returns true if the radius is constant 
    --          all along the edge E.
    is static;
    
    Radius(me) returns Real from Standard;
    ---Purpose: returns the radius if the fillet is constant
    --          all along the spine.

    Radius(me; IE : Integer from Standard) 
    returns Real from Standard;
    ---Purpose: returns the radius if the fillet is constant
    --          all along the edge E.

    Radius(me; E : Edge from TopoDS) 
    returns Real from Standard;
    ---Purpose: returns the radius if the fillet is constant
    --          all along the edge E.

    ComputeLaw(me : mutable; Els : HElSpine from ChFiDS) 
    returns Composite from Law
    is private;
    
    AppendElSpine(me : mutable; Els : HElSpine from ChFiDS) 
    is redefined;
    
    AppendLaw(me : mutable; Els : HElSpine from ChFiDS) 
    is private;
    
    Law(me; Els : HElSpine from ChFiDS) 
    returns Composite from Law
    is static;
    
    ChangeLaw(me : mutable; E : Edge from TopoDS) 
    ---C++: return &
    returns Function from Law
    ---Purpose: returns the elementary law 
    is static;

    MaxRadFromSeqAndLaws(me) returns Real from Standard;
    ---Purpose: returns the maximum radius if the fillet is non-constant

fields

--radius    : HArray1OfReal from TColStd;
parandrad : SequenceOfXY  from TColgp;
laws      : Laws          from Law;

end FilSpine;


