-- File:	BOPTools_PaveFiller.cdl
-- Created:	Thu Feb  8 14:07:33 2001
-- Author:	Peter KURNEV
--		<pkv@irinox>
---Copyright:	 Matra Datavision 2001


class PaveFiller from BOPTools 

	---Purpose:  The algorithm that provides  
        ---  1. creation of the data structure (DS)    	 
        ---  2. creation of the interferences' pool   	 
        ---  3. invocation of Perform() to fill the DS 
    	---   
        ---
uses
    
    PShapesDataStructure    from BooleanOperations, 
    
    InterferencePool        from BOPTools,  
    PInterferencePool       from BOPTools,  
    PavePool                from BOPTools, 
    CommonBlockPool         from BOPTools, 
    SplitShapesPool         from BOPTools, 
    
    Pave                    from BOPTools,  
    PaveBlock               from BOPTools,  
    PaveSet                 from BOPTools, 
    Curve                   from BOPTools,
    SSInterference          from BOPTools, 
    ListOfPaveBlock         from BOPTools, 
    IteratorOfCoupleOfShape from BOPTools, 
    SSInterference          from BOPTools, 
    SSIntersectionAttribute from BOPTools, 
    ShrunkRange             from IntTools, 
    Context                 from IntTools, 
    
    ShapeEnum           from  TopAbs, 
    ListOfInteger       from TColStd, 
    IndexedMapOfInteger from TColStd, 
    
    Pnt     from gp,
    Vertex  from TopoDS,
    SetOfInteger  from  TColStd


is 
 
    Create   
    	returns PaveFiller from BOPTools; 
    	---Purpose:  
    	--- Empty Contructor  
    	---
    Create  (aIP: InterferencePool from BOPTools) 
    	returns PaveFiller from BOPTools; 
    	---Purpose:   
    	--- Constructor 
    	---
    Create  (theIP              : InterferencePool from BOPTools;
    	     theSectionAttribute: SSIntersectionAttribute from BOPTools) 
    	returns PaveFiller from BOPTools; 
    	---Purpose:   
    	--- Constructor
    	---
    Destroy (me: in out) 
	is  virtual;     
    	---C++: alias "Standard_EXPORT virtual ~BOPTools_PaveFiller(){Destroy();}"     
    	---Purpose:   
    	--- Destructor
    	---
    Perform    (me:out) 
	is virtual;       
    	---Purpose:
    	--- Fills the DS               
    	---
 
    PartialPerform(me:out; anObjSubSet, aToolSubSet:  SetOfInteger  from  TColStd) 
	is virtual;       
       
    ToCompletePerform(me:out)		   
	is virtual;       
 
    PerformVV  (me:out) 
    	is  virtual protected; 
    	---Purpose:
    	--- Computes Vertex/Vertex interferences                
    	---
    PerformVE  (me:out) 
    	is  virtual protected;  
    	---Purpose:
    	--- Computes Vertex/Edge interferences                
    	---
    PerformVF  (me:out) 
    	is  virtual protected;  
    	---Purpose:
    	--- Computes Vertex/Face interferences                
    	---
    PerformEE  (me:out) 
    	is  virtual protected;  
    	---Purpose:
    	--- Computes Edge/Edge interferences                
    	---
    PerformEF  (me:out) 
    	is  virtual protected; 
    	---Purpose:
    	--- Computes Edge/Face interferences                
    	---
    PerformFF  (me:out) 
    	is  virtual protected;   
    	---Purpose:
    	--- Computes Face/Face interferences                
    	---

    -------------------------------------------------------------- 
    --- 
    ---	  Selectors   
    ---   
    --- 
    SetContext(me:out; 
    	    aContext:  Context from IntTools); 
    	---Purpose:
    	--- Sets the intersecton context                 
    	---   
    Context(me) 
    	 returns Context from IntTools; 
    	---C++:return const &	
    	---Purpose:
    	--- Selector                
    	---
--    ChangeContext(me:out) 
--    	 returns Context from IntTools;  
    	--  C++:return &	
    	---Purpose:
    	--- Selector                
    	---
    SetInterferencePool(me:out; 
    	 aPool:InterferencePool from BOPTools); 
    	---Purpose:
    	--- Selector                
    	---
    IsDone(me) 
    	returns  Boolean  from  Standard;  
    	---Purpose:
    	--- Selector
    	---
    PavePool(me) 
    	returns  PavePool from BOPTools; 
    	---C++:return const &	 
    	---Purpose:
    	--- Selector               
    	---
    ChangePavePool(me:out) 
    	returns  PavePool from BOPTools; 
    	---C++:return &	
   	---Purpose:
    	--- Selector               
    	---
    CommonBlockPool(me) 
    	returns  CommonBlockPool from BOPTools; 
    	---C++:return const &	 
    	---Purpose:
    	--- Selector               
    	---
    ChangeCommonBlockPool(me:out) 
    	returns  CommonBlockPool from BOPTools; 
    	---C++:return &	
    	---Purpose:
    	--- Selector               
    	---
    SplitShapesPool(me)  
    	returns  SplitShapesPool from BOPTools;
    	---C++:return const &	
    	---Purpose:
    	--- Selector               
    	---

    ChangeSplitShapesPool(me:out)  
    	returns  SplitShapesPool from BOPTools;
    	---C++:return  &	
    	---Purpose:
    	--- Selector               
    	---
    DS(me:out) 
    	returns PShapesDataStructure from BooleanOperations;  
    	---Purpose:
    	--- Selector               
    	---
    InterfPool(me:out) 
    	returns PInterferencePool from BOPTools; 
    	---Purpose:
    	--- Selector               
    	---
 
    IteratorOfCoupleOfShape(me)  
    	returns  IteratorOfCoupleOfShape from BOPTools;
    	---C++:return const &	
    	---Purpose:
    	--- Selector               
	---
      
    SectionAttribute(me)
    	returns SSIntersectionAttribute from BOPTools;
    	---C++: return const &
    	---Purpose:
    	--- Selector   
	---

    SetSectionAttribute(me:out; 
    	anAtt  :  SSIntersectionAttribute from BOPTools);
    	---Purpose:
    	--- Selector       
	---
    -------------------------------------------------------------- 
    ---	     
    ---  PaveBlocks for Split Parts of Edges.  
    ---     
    --- 
    SortTypes      (me;   
    	    anInd1:in out Integer from Standard; 
            anInd2:in out Integer from Standard) 
    	is protected;  
    	---Purpose:
    	--- Sorts the types of shapes with DS-indices  
    	--- <anInd1> and  <anInd2> in increasing order of  
    	--- types of the shapes               
    	---
    PerformNewVertices  (me:out) 
    	is protected;     	     
     
    IsSuccesstorsComputed (me;  
    	    iF1:Integer from  Standard; 
    	    iF2:Integer from  Standard) 
    	returns  Boolean from Standard 
    	is protected;    
     
    PrepareEdges  (me:out) 
    	is virtual protected;  
    	---Purpose:   
    	--- Prepare end paves for each edge 
    	---
    PreparePaveBlocks (me:out; 
    	    	    	aType1: ShapeEnum  from  TopAbs; 
    	    	    	aType2: ShapeEnum  from  TopAbs) 
    	is virtual protected; 
    	---Purpose:   
    	--- Prepare PaveBlocks  for  each  edge  (EE-interferences) 
    	---
    PreparePaveBlocks (me:out;   
    	    	       anE:Integer from Standard) 
    	is virtual protected;  
    	---Purpose:  
    	--- Prepare PaveBlocks for given edge (EE-interferences) 
    	---
    RefinePavePool(me:out) 
    	is protected;  
    	---Purpose:  
    	--- Refines myPavePool taking into account new Paves obtained from EE algo 
    	---
    MakeSplitEdges(me:out) 
    	is protected;   
    	---Purpose:  
    	--- Makes split edges from source edges 
    	---
    DoSDEdges(me:out) 
    	is protected;    
    	---Purpose:
    	--- Update Lists of PaveBlocks with info about 
    	--- indices of split edges that are Same Domain 
    	--- with other splits or faces 
    	---
    CorrectShrunkRanges(me:out; 
    	    	    	aSide:  Integer  from  Standard; 
    	    	    	aPave:  Pave from BOPTools; 
    	    	    	aSR  :  out ShrunkRange  from  IntTools)
    	is protected;  
    	---Purpose:
    	--- Update Shrunk  Range <aSR> for Pave <aPave> 
    	---
    SplitIndex  (me:out;  aPB:PaveBlock from BOPTools)  
    	returns Integer from Standard 
    	is protected;  
    	---Purpose:  
    	--- Returns  the Index of Split edge for the PaveBlock <aPB> 
    	--- in  DS. 
    	--- If the PaveBlock is not found, returns 0; 
    	---
    IsBlocksCoinside (me; 
    	aPB1:PaveBlock from BOPTools;
    	aPB2:PaveBlock from BOPTools) 
	returns Boolean from Standard 
    	is protected;   
    	---Purpose: 	 
    	--- Returns  TRUE if the two PaveBlocks have vertices 
    	--- that touch each other in terms of Tolerances of 
    	--- the vertices 	     
    	---
    -------------------------------------------------------------- 
    ---	  
    ---  Some of API FUNCTIONS  
    --- 
    --- 
    SplitsInFace(me:out; 
    	         aBid:Integer from Standard;  
    	         nF1 :Integer from Standard;  
    	         nF2 :Integer from Standard;  
    	         aLs :out ListOfInteger from TColStd) 
    	returns Integer from Standard;  
    	---Purpose:  
    	--- For the face <nF1> get all splits that are IN-2D          
    	--- to  the face <nF2>; The result is in <aLs> 
    	--- Returns 0 if OK; 
    	---
    SplitsInFace(me:out; 
    	         nE1 :Integer from Standard;  
    	         nF2 :Integer from Standard;  
    	         aLs :out ListOfInteger from TColStd) 
    	returns Integer from Standard;  
    	---Purpose:  
    	--- For the edge <nE1> get all splits that are IN-2D          
    	--- to  the face <nF1>; The result is in <aLs> 
    	--- Returns 0 if OK; 
    	---
    SplitsOnEdge(me:out; 
    	         nE1 :Integer from Standard;  
    	         nE2 :Integer from Standard;  
    	         aLs :out ListOfInteger from TColStd) 
    	returns Integer from Standard;  
    	---Purpose:  
    	--- For the edge <nE1> get all splits that are ON-3D          
    	--- to  the edge <nE2>; The result is in <aLs> 
    	--- Returns 0 if OK; 
    	---
    SplitsOnFace(me:out; 
    	         nE1 :Integer from Standard;  
    	         nF2 :Integer from Standard;  
    	         aLs :out ListOfInteger from TColStd) 
    	returns Integer from Standard;  
    	---Purpose:  
    	--- For the edge <nE1> get all splits that are ON-3D          
    	--- to  the face <nF2>; The result is in <aLs> 
    	--- Returns 0 if OK; 
    	---
    SplitsOnFace(me:out;  
    	         aBid:Integer from Standard;  
    	         nF1 :Integer from Standard;  
    	         nF2 :Integer from Standard;  
    	         aLs :out ListOfInteger from TColStd) 
    	returns Integer from Standard;  
    	---Purpose:  
    	--- For the face <nF1> get all splits that are ON-3D          
    	--- to  the face <nF2>; The result is in <aLs> 
    	--- Returns 0 if OK; 
    	---
     
    SplitsInFace(me:out; 
    	         aBid:Integer from Standard;  
    	         nF1 :Integer from Standard;  
    	         nF2 :Integer from Standard;  
    	         aLs :out ListOfPaveBlock from BOPTools) 
    	returns Integer from Standard;  
    	---Purpose:  
    	--- For the face <nF1> get all PaveBlocks that are IN-2D          
    	--- to  the face <nF2>; The result is in <aLs> 
    	--- Returns 0 if OK; 
    	---
     
    SplitsInFace(me:out; 
    	         nE1 :Integer from Standard;  
    	         nF2 :Integer from Standard;  
    	         aLs :out ListOfPaveBlock from BOPTools) 
    	returns Integer from Standard;  
    	---Purpose:   
    	--- For the edge <nE1> get all PaveBlocks that are IN-2D          
    	--- to  the face <nF1>; The result is in <aLs> 
    	--- Returns 0 if OK; 
    	---
     
    SplitsOnEdge(me:out; 
    	         nE1 :Integer from Standard;  
    	         nE2 :Integer from Standard;  
    	         aLs :out ListOfPaveBlock from BOPTools) 
    	returns Integer from Standard;  
    	---Purpose:   
    	--- For the edge <nE1> get all PaveBlocks that are ON-3D          
    	--- to  the edge <nE2>; The result is in <aLs> 
    	--- Returns 0 if OK; 
    	---
     
    SplitsOnFace(me:out; 
    	         nE1 :Integer from Standard;  
    	         nF2 :Integer from Standard;  
    	         aLs :out ListOfPaveBlock from BOPTools) 
    	returns Integer from Standard;  
    	---Purpose:  
    	--- For the edge <nE1> get all PaveBlocks that are ON-3D          
    	--- to  the face <nF2>; The result is in <aLs> 
    	--- Returns 0 if OK; 
    	---

    SplitsOnFace(me:out;  
    	         aBid:Integer from Standard;  
    	         nF1 :Integer from Standard;  
    	         nF2 :Integer from Standard;  
    	         aLs :out ListOfPaveBlock from BOPTools) 
    	returns Integer from Standard;  
    	---Purpose: 
    	--- For the face <nF1> get all PaveBlocks that are ON-3D          
    	--- to  the face <nF2>; The result is in <aLs> 
    	--- Returns 0 if OK; 
    	---
    FindSDVertex (me; 
    	    	    nV:  Integer  from  Standard) 
    	returns Integer from Standard; 
    	---Purpose:
    	--- Find  for the vertex <nV> SD-vertex (if possible) and return  
    	--- its DS-index.  Otherwise it returns 0.
	---
     
    --------------------------------------------------------------- 
    ---	  
    ---   Section  Edges.  Protected Block.
    --- 
    ---	     
    MakeBlocks(me:out) 
    	is protected; 
    	---Purpose: 
    	--- Make Pave Blocks for intersection curves    
    	---
    MakeAloneVertices(me:out) 
    	is protected; 
    	---Purpose: 
    	--- Make vertices that are place of intersection  
    	--- between faces       
    	---
    PutPaveOnCurve(me:out; 
    	    	   aPaveSet: PaveSet from BOPTools; 
		   aTolR3D : Real from Standard; 				   		     
    	    	   aBCurve :out Curve from BOPTools) 
       	is protected;   
    	---Purpose: 
    	--- Among Paves from <aPaveSet> find ones that belong 
    	--- to intersection curve <aBCurve> with 3D-tolerance  
    	--- value <aTolR3D>
    	---
    PutPaveOnCurve(me:out; 
    	    	   aPave   : Pave from BOPTools; 
    	    	   aTolR3D : Real from Standard;  
    	    	   aBCurve :out Curve from BOPTools) 
       	is protected;     
    	---Purpose: 
    	--- Try to put Pave <aPave> on intersection curve <aBCurve>  
    	--- with 3D-tolerance value <aTolR3D>
    	---

    PutPavesOnCurves(me:out)
    	is protected;

    PrepareSetForFace(me:out;  
    	    	    nF1 :Integer from Standard;  
    	    	    nF2 :Integer from Standard;  
	    	    aPaveSet:out PaveSet from BOPTools); 
    	---Purpose:  
    	--- For couple of faces <nF1>, <nF2> prepare set of all paves 
    	--- of all edges <aPaveSet>
    	---
    MakeSectionEdges(me:out) 
    	is protected;  
    	---Purpose:  
    	--- For all inrefered faces make section edges from  
    	--- intersection curves and corresp.  Paves on them      
    	---
    PutBoundPaveOnCurve (me:out; 
    	    	    aBC :out Curve from BOPTools;	 
     	    	    aFF :out SSInterference from BOPTools) 
    	is protected; 
    	---Purpose: 	     
    	--- Try to  put own  bounds of the curve on the curve <aBC> 
    	---
    PutBoundPaveOnCurve (me:out;  
    	    	    aP  : Pnt from  gp; 
		    aT  : Real from Standard; 			 
    	    	    aBC :out Curve from BOPTools;	 
     	    	    aFF :out SSInterference from BOPTools) 
    	is protected;  
    	---Purpose: 	     
    	--- Try to put 3D-point <aP> (parameter aT)  on the curve <aBC> 
    	---
    PutBoundPaveOnCurveSpec (me:out; 
    	    	    aBC :out Curve from BOPTools;	 
     	    	    aFF :out SSInterference from BOPTools) 
    	is protected; 
    	---Purpose: 	     
    	--- Try to  put own  bounds of the curve on the curve <aBC> 
    	--- 
    PutBoundPaveOnCurveSpec (me:out;  
    	    	    aP  : Pnt from  gp; 
		    aT  : Real from Standard; 			 
    	    	    aBC :out Curve from BOPTools;	 
     	    	    aFF :out SSInterference from BOPTools) 
    	is protected;  
    	---Purpose: 	     
    	--- Try to put 3D-point <aP> (parameter aT)  on the curve <aBC> 
    	--- 
 
--modified by NIZNHY-PKV Thu Oct 20 07:17:11 2011f 
    PutClosingPaveOnCurve (me:out; 
    	    	    aBC :out Curve from BOPTools;	 
     	    	    aFF :out SSInterference from BOPTools)  
	is protected; 
	---Purpose: 	     
    	--- Put paves on the curve <aBC> in case when <aBC>   
        --  is closed 3D-curve  
    	---      
--modified by NIZNHY-PKV Thu Oct 20 07:17:11 2011t	 

    FindPave            (me:out; 
		    aP  :Pnt from  gp;  
    	    	    aTpV: Real from Standard;  
    	    	    aPS: PaveSet from BOPTools; 
		    aPV:out Pave from BOPTools) 
    	returns Boolean from Standard
       	is protected; 
    	---Purpose: 	     
    	--- Returns TRUE if 3D-point <aP> coinsides with some Pave 
    	--- from <aPS> (with 3D-tolerance value <aTpV>); 
    	--- In  TRUE case <aPV> will contain the Pave  .      	     
    	---
    CheckCoincidence(me:out;  
    	    	    aPB: PaveBlock      from BOPTools;  
     	    	    aFF: SSInterference from BOPTools) 
    	returns Boolean from Standard 
    	is protected;  
    	---Purpose: 	     
    	--- Returns TRUE if PaveBlock <aPB> lays on the faces 
    	--- from FF-interference <aFF> 
    	---
    CheckIntermediatePoint(me:out;  
    	    	    aPB : PaveBlock      from BOPTools;  
    	    	    aPBR: PaveBlock      from BOPTools;  
     	    	    aTol: Real  from  Standard) 
    	returns Integer from Standard 
    	is protected;  
    	---Purpose: 	     
    	--- Returns 0 if some arbitrary intermediate point from   
    	--- PaveBlock <aPB> lays on the PaveBlock  <aPBR> 
    	--- (with 3D-tolerance value <aTol>)
    	---
 
    CheckFacePaves(me:out;  
    	    	    aV : Vertex  from TopoDS;  
     	    	    nF:  Integer from Standard) 
    	returns Integer from Standard 
    	is protected; 
    	---Purpose: 	 
    	--- Internal  usage 
    	---
    StickVertices (me:out;   
    	    	    nF1:  Integer from Standard;
    	    	    nF2:  Integer from Standard; 
		    aMV:out IndexedMapOfInteger from TColStd) 
	is protected; 	    
    	---Purpose: 	 
    	--- Internal  usage 
    	---
    ExpectedPoolLength(me) 
    	returns  Integer from Standard 
	is protected;
    	---Purpose: 	 
    	--- Returns the value of expected length of array of interferences 
    	---

    RestrictCurveIn2d(me: in out; nE, nF1, nF2    : Integer from Standard;
    	    			theTolerance: Real from Standard;
			     	theBC       : in out Curve from BOPTools)
    	is private;

    RecomputeCommonBlocks(me: in out; nE: Integer from Standard)
    	is private;

    ExtendedTolerance(me:out; 
    	    nV      : Integer from Standard; 
            aTolExt : out Real from Standard) 
	returns Boolean from Standard 		     
	is  protected;		     

fields 
 
    myIntrPool         :  PInterferencePool from BOPTools
    	is protected;
    myDS               :  PShapesDataStructure from BooleanOperations 
    	is protected;   
    myPavePool         :  PavePool from BOPTools 
    	is protected; 
    myPavePoolNew      :  PavePool from BOPTools 
    	is protected; 
    myCommonBlockPool  :  CommonBlockPool from BOPTools 
    	is protected;  
    mySplitShapesPool  :  SplitShapesPool from BOPTools 
    	is protected; 
    mySectionAttribute :  SSIntersectionAttribute from BOPTools 
    	is protected;
    myNbSources        :  Integer from Standard 
    	is protected; 
    myNbEdges          :  Integer from Standard 
    	is protected;      
    myIsDone           :  Boolean from Standard 
    	is protected; 
    myDSIt             :  IteratorOfCoupleOfShape from BOPTools 
    	is protected; 
    myContext           :  Context from IntTools 
    	is protected;  	     

end PaveFiller;
