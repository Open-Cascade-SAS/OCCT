-- Created on: 1993-01-22
-- Created by: Gilles DEBARBOUILLE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class MethodDefinition from Dynamic

inherits

    Method from Dynamic
    
	---Purpose: This  inherited class   is   for  describing   the
	--          definition  of    a  method.   This  definition is
	--          composed by its name which is readable by the type
	--          function   and a  collection   of  variables which
	--          defines the signature  of the method definition in
	--          term of arguments passed  to the function and also
	--          the useful  internal or constant  variables if the
	--          function is a composite method. This class is also
	--          a  deferred  class and can   not be  used directly
	--          because it is  necessary to specify if the  method
	--          is compiled, interpreted or composite.

uses

    CString from Standard,
    OStream from Standard,
    HAsciiString from TCollection,
    AsciiString  from TCollection,
    Parameter    from Dynamic,
    ModeEnum     from Dynamic


is

    Initialize(aname : CString from Standard);
    
    ---Level: Internal 
    
    ---Purpose: Creates a MethodDefinition with <aname> as type.
    
    Type(me) returns AsciiString from TCollection
    
    ---Level: Advanced 
    
    ---Purpose: Returns the name of the method definition.
    
    is redefined;
    
    AddVariable(me : mutable ; aparameter : Parameter from Dynamic ;
                               amode      : ModeEnum  from Dynamic ;
                               agroup     : Boolean = Standard_False)
    
    ---Level: Advanced 
    
    ---Purpose: Adds  a  new  variable   created from    the parameter
    --          <aparameter>, which  defines the  name of the variable
    --          its type and if necessary its  default value, the mode
    --          <amode> which  precise  if it is  an  in,  out, inout,
    --          internal or   constant variable and the  flag <agroup>
    --          for accepting  a  set of homogeneous variables.   with
    --          the parameter value <aparameter>.
    
    is static;
    
    Dump(me ; astream : in out OStream from Standard)
    
    ---Level: Internal 
    
    ---Purpose: Useful for debugging.

    is redefined;
    
fields

    thename : HAsciiString from TCollection;

end MethodDefinition;
