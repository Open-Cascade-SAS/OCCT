-- Created on: 1993-06-14
-- Created by: Martine LANGLOIS
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MakeBSplineCurveWithKnotsAndRationalBSplineCurve from GeomToStep inherits
    Root from GeomToStep

    ---Purpose: This class implements the mapping between classes
    --          BSplineCurve from Geom, Geom2d and the class
    --          BSplineCurveWithKnotsAndRationalBSplineCurve from StepGeom
    --          which describes a rational_bspline_curve_with_knots from
    --          Prostep
  
uses

     BSplineCurve from Geom,
     BSplineCurve from Geom2d,
     BSplineCurveWithKnotsAndRationalBSplineCurve from StepGeom
     
raises

     NotDone from StdFail
     
is 

Create ( Bsplin : BSplineCurve from Geom ) returns
    MakeBSplineCurveWithKnotsAndRationalBSplineCurve;

Create ( Bsplin : BSplineCurve from Geom2d ) returns
    MakeBSplineCurveWithKnotsAndRationalBSplineCurve;
Value (me) returns
    BSplineCurveWithKnotsAndRationalBSplineCurve from StepGeom
    raises NotDone
    is static;
    ---C++: return const&
    
fields

    theBSplineCurveWithKnotsAndRationalBSplineCurve :
    	BSplineCurveWithKnotsAndRationalBSplineCurve from StepGeom;
    	-- The solution from StepGeom
    	
end MakeBSplineCurveWithKnotsAndRationalBSplineCurve;
