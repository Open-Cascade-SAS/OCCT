-- Created on: 1995-03-22
-- Created by: Laurent BUCHARD
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class FClass2d from BRepTopAdaptor

uses  
    Pnt2d             from gp,
    Face              from TopoDS,
    State             from TopAbs,
    SequenceOfInteger from TColStd,
    SeqOfPtr          from BRepTopAdaptor    

is 

    Create(F: Face from TopoDS; Tol: Real from Standard)
    returns FClass2d from BRepTopAdaptor;

    
    PerformInfinitePoint(me) 
    returns State from TopAbs;
    
    Perform(me; Puv: Pnt2d from gp; RecadreOnPeriodic: Boolean from Standard  =  Standard_True) 
    returns State from TopAbs;
    
    Destroy(me: in out);
    	---C++: alias ~
    

    Copy(me; Other: FClass2d from BRepTopAdaptor)
    returns FClass2d from BRepTopAdaptor;
    	---C++: return const &
      	---C++: alias operator=
     --Purpose *** Raise if called ***


    TestOnRestriction(me; Puv: Pnt2d from gp; 
                          Tol: Real from Standard;
                          RecadreOnPeriodic: Boolean from Standard  =  Standard_True) 
    returns State from TopAbs;
    ---Purpose: Test a point with +- an offset (Tol) and returns
    --          On if some points are OUT an some are IN
    --          (Caution: Internal use . see the code for more details)




fields 

    TabClass    : SeqOfPtr          from BRepTopAdaptor;
    TabOrien    : SequenceOfInteger from TColStd;
    Toluv       : Real              from Standard;
    Face        : Face              from TopoDS;
    U1          : Real              from Standard;
    V1          : Real              from Standard;    
    U2          : Real              from Standard;
    V2          : Real              from Standard;
    
    Umin        : Real              from Standard;  
    Umax        : Real              from Standard;
    Vmin        : Real              from Standard;  
    Vmax        : Real              from Standard;


end FClass2d from BRepTopAdaptor;
