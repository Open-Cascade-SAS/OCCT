-- Created on: 1999-04-01
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Marker from TopOpeBRepDS inherits TShared from MMgt    	
uses
    HArray1OfBoolean from TColStd,
    AsciiString from TCollection
is
    Create returns mutable Marker;
    Reset(me:mutable);
    Set(me:mutable;i:Integer;b:Boolean);
    Set(me:mutable;b:Boolean;n:Integer;a:Address);
    GetI(me;i:Integer) returns Boolean;
    Allocate(me:mutable;n:Integer);    
fields
    myhe : HArray1OfBoolean from TColStd;
    myne : Integer;   
end Marker from TopOpeBRepDS;
