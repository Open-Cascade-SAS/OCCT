-- Created on: 1993-07-06
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class Curve3D from BRep inherits GCurve from BRep

	---Purpose: Representation of a curve by a 3D curve.

uses
    Pnt                 from gp,
    Location            from TopLoc,
    Curve               from Geom,
    CurveRepresentation from BRep

is

    Create(C : Curve    from Geom;
    	   L : Location from TopLoc) 
    returns mutable Curve3D from BRep;

    D0(me; U : Real; P : out Pnt from gp);
	---Purpose: Computes the point at parameter U.

    IsCurve3D(me) returns Boolean
	 ---Purpose: Returns True.
    is redefined;
	
    Curve3D(me) returns any Curve from Geom
	---C++: return const &
    is redefined;

    Curve3D(me : mutable; C : Curve from Geom)
    is redefined;
	
    Copy(me) returns mutable CurveRepresentation from BRep;
	---Purpose: Return a copy of this representation.

fields
    
    myCurve : Curve from Geom;

end Curve3D;
