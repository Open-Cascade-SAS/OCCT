-- Created on: 1993-02-22
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class LineOn2S from IntSurf 

	---Purpose: 

inherits TShared from MMgt


uses Allocator         from IntSurf,
     PntOn2S           from IntSurf,
     SequenceOfPntOn2S from IntSurf

raises OutOfRange from Standard

is

    Create (theAllocator: Allocator from IntSurf = 0)
    
    	returns LineOn2S from IntSurf;
	

    Add(me: mutable; P: PntOn2S from IntSurf)
    
	---Purpose: Adds a point in the line.

	---C++: inline

    	is static;


    NbPoints(me)
    
	---Purpose: Returns the number of points in the line.

    	returns Integer from Standard
	---C++: inline
	
	is static;


    Value(me; Index: Integer from Standard)
    
	---Purpose: Returns the point of range Index in the line.
    
    	returns PntOn2S from IntSurf
	---C++: inline
	---C++: return const&
	
	raises OutOfRange from Standard
	--- The exception OutOfRange is raised when Index <= 0 or
	--  Index > NbPoints.
	
	is static;


    Reverse(me: mutable)
    
	---Purpose: Reverses the order of points of the line.

	---C++: inline

    	is static;



    Split(me: mutable;Index: Integer from Standard)

	---Purpose: Keeps in <me> the points 1 to Index-1, and returns
	--          the items Index to the end.

    	returns LineOn2S from IntSurf

    	raises OutOfRange from Standard
	--- The exception OutOfRange is raised when Index <= 0 or
	--  Index > NbPoints.

	is static;


    Value(me: mutable; Index: Integer from Standard; P: PntOn2S from IntSurf)
    
	---Purpose: Replaces the point of range Index in the line.
    
	raises OutOfRange from Standard
	--- The exception OutOfRange is raised when Index <= 0 or
	--  Index > NbPoints.
	
	---C++: inline
        
	is static;
	
	
    SetUV(me: mutable; Index: Integer from Standard;
    	               OnFirst: Boolean from Standard;
		       U,V: Real from Standard)
    
	---Purpose: Sets the parametric coordinates on one of the surfaces
	--          of the point of range Index in the line.
    
	---C++: inline
        
	raises OutOfRange from Standard
	--- The exception OutOfRange is raised when Index <= 0 or
	--  Index > NbPoints.
	
	is static;
	
	
    Clear(me: mutable)
    
	---C++: inline
        
    	is static;


    InsertBefore(me:mutable; I: Integer from Standard; P: PntOn2S from IntSurf) 
    
    	is static;

    RemovePoint(me:mutable; I: Integer from Standard)
    
    	is static;


fields

    mySeq: SequenceOfPntOn2S from IntSurf;

end LineOn2S;
