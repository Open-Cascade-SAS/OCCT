-- File:        FunctionSet.cdl
-- Created:     Mon May 13 15:21:04 1991
-- Author:      Laurent PAINNOT
--              <lpa@topsn3>
--Copyright:     Matra Datavision 1991


deferred class FunctionSet from math
    	---Purpose:
    	-- This abstract class describes the virtual functions associated to
    	-- a set on N Functions of M independant variables.

uses Vector from math

is

    Delete(me:out) is virtual;
    	---C++: alias "Standard_EXPORT virtual ~math_FunctionSet(){Delete();}"
    
    NbVariables(me)
    	---Purpose: Returns the number of variables of the function.

    returns Integer
    is deferred;
    
    
    NbEquations(me)
    	---Purpose: Returns the number of equations of the function.

    returns Integer
    is deferred;
    
    
    Value(me: in out; X: Vector; F: out Vector)
    	---Purpose: Computes the values <F> of the functions for the 
    	--          variable <X>.
    	--          returns True if the computation was done successfully, 
    	--          False otherwise.

    returns Boolean
    is deferred;
    

    GetStateNumber(me: in out)
    	---Purpose: Returns the state of the function corresponding to the
    	--          latestcall of any methods associated with the function.
    	--          This function is called by each of the algorithms 
    	--          described later which define the function Integer 
    	--          Algorithm::StateNumber(). The algorithm has the 
    	--          responsibility to call this function when it has found
    	--          a solution (i.e. a root or a minimum) and has to maintain
    	--          the association between the solution found and this
    	--          StateNumber.
    	--          Byu default, this method returns 0 (which means for the 
    	--          algorithm: no state has been saved). It is the 
    	--          responsibility of the programmer to decide if he needs
    	--          to save the current state of the function and to return
    	--          an Integer that allows retrieval of the state.

    returns Integer
    is virtual;
    
end FunctionSet;


