-- Created on: 1992-11-05
-- Created by: Remi LEQUETTE
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Torus from BRepPrim inherits Revolution from BRepPrim

	---Purpose: Implements the torus primitive

uses
    Face from TopoDS,
    
    Pnt from gp,
    Ax2 from gp    

raises
    DomainError

is
    Create(Position : Ax2 from gp; Major : Real; Minor : Real)
    returns Torus from BRepPrim
	   ---Purpose: the STEP definition
	   --          Position : center and axes
	   --          Major, Minor : Radii
	   --          
	   --          Errors : Major < Resolution
	   --                   Minor < Resolution
    raises DomainError;

    Create(Major,Minor : Real)
    returns Torus from BRepPrim
	---Purpose: Torus centered at origin
    raises DomainError;
    
    Create(Center : Pnt from gp; Major, Minor : Real)
    returns Torus from BRepPrim
	---Purpose: Torus at Center
    raises DomainError;
    
    MakeEmptyLateralFace(me) returns Face from TopoDS
	---Purpose: The surface normal should be directed  towards the
	--          outside.
    is redefined;
    
    SetMeridian(me : in out)
    is static private;
    
fields
    myMajor     : Real;
    myMinor     : Real;

end Torus;
