-- Created on: 1996-09-13
-- Created by: DCB
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Driver from CGM inherits PlotterDriver from PlotMgt
  ---Purpose: This class defines a CGM (Computer Graphic Metafile) plotter Driver.
  ---         All necessary information about methods (purpose, level, category, etc.)
  ---         can be found in CDL files from the inheritance tree (PlotMgt_PlotterDriver,
  ---         Aspect_Driver).

uses
  Plotter                 from PlotMgt,
  ExtendedString          from TCollection,
  ColorMap                from Aspect,
  TypeMap                 from Aspect,
  WidthMap                from Aspect,
  TypeOfText              from Aspect,
  TypeOfColorSpace        from Aspect,
  PlaneAngle              from Quantity,
  Length                  from Quantity,
  Factor                  from Quantity,
  Ratio                   from Quantity,
  Array1OfShortReal       from TShort


is
  Create(aPlotter          : Plotter from PlotMgt;
         aName             : CString from Standard;
         aDX,aDY           : Length from Quantity;
         aTypeOfColorSpace : TypeOfColorSpace from Aspect = Aspect_TOCS_RGB) 
  returns mutable Driver from CGM;


  Create(aName             : CString from Standard;
         aDX,aDY           : Length from Quantity;
         aTypeOfColorSpace : TypeOfColorSpace from Aspect = Aspect_TOCS_RGB) 
  returns mutable Driver from CGM;


  BeginFile(me: mutable;
            aPlotter          : Plotter from PlotMgt;
            aDX,aDY           : Length from Quantity;
            aTypeOfColorSpace : TypeOfColorSpace from Aspect)
  is private;
  
  Close(me: mutable)
  is redefined protected;
  ---C++: alias ~ 


  BeginDraw (me: mutable)
  is redefined;


  EndDraw (me: mutable; dontFlush: Boolean = Standard_False)
  is redefined;


  ---------------------------------------------
  -- Category: Methods to define the attributes
  ---------------------------------------------
  InitializeColorMap(me: mutable; aColorMap: ColorMap from Aspect) 
  is redefined protected;


  InitializeTypeMap(me: mutable; aTypeMap: TypeMap from Aspect)
  is redefined protected;


  InitializeWidthMap(me: mutable; aWidthMap: WidthMap from Aspect)
  is virtual protected;


  -----------------------------------------
  -- Category: Methods to manage the images
  -----------------------------------------
  SizeOfImageFile (me; anImageFile: CString from Standard;
                       aWidth,aHeight: out Integer from Standard)
  returns Boolean from Standard is redefined;


  --------------------------------
  -- Actual set graphic attributes
  --------------------------------
  PlotLineAttrib (me: mutable;
    ColorIndex: Integer from Standard;
    TypeIndex: Integer from Standard;
    WidthIndex: Integer from Standard)
  is redefined protected;


  PlotPolyAttrib (me: mutable;
    ColorIndex: Integer from Standard;
    TileIndex: Integer from Standard;
    DrawEdge: Boolean from Standard)
  is redefined protected;


  -----------------------------------------------
  -- Category: Private methods to draw primitives
  -----------------------------------------------
  PlotPoint (me : mutable; X, Y: ShortReal from Standard)
  returns Boolean from Standard
  is redefined protected;


  PlotSegment (me : mutable;
      X1, Y1: ShortReal from Standard;
      X2, Y2: ShortReal from Standard)
  returns Boolean from Standard
  is redefined protected;


  PlotPolyline (me : mutable;
      xArray : Address from Standard;
      yArray : Address from Standard;
      nPts   : Address from Standard;
      nParts : Integer from Standard)
  returns Boolean from Standard
  is redefined protected;


  PlotPolygon (me : mutable;
      xArray : Address from Standard;
      yArray : Address from Standard;
      nPts   : Address from Standard;
      nParts : Integer from Standard)
  returns Boolean from Standard
  is redefined protected;


  PlotArc (me : mutable; X,Y : ShortReal from Standard;
      anXradius,anYradius : ShortReal from Standard;
      sAngle: ShortReal from Standard;
      oAngle: ShortReal from Standard)
  returns Boolean from Standard
  is redefined protected;


  PlotPolyArc (me : mutable; X,Y : ShortReal from Standard;
      anXradius,anYradius : ShortReal from Standard;
      sAngle: ShortReal from Standard;
      oAngle: ShortReal from Standard)
  returns Boolean from Standard
  is redefined protected;


  PlotImage (me: mutable; 
      aX, aY, aWidth:  ShortReal from Standard;
      aHeight, aScale: ShortReal from Standard;
      anImageFile:     CString   from Standard;
      anArrayOfPixels: Address   from Standard;
      aLineIndex:      Integer   from Standard = -1)
  returns Boolean from Standard
  is redefined protected;


  InitializeDriver  (me:  mutable; aName: CString from Standard)
  is  private;


  WriteData (me: mutable; 
    aCode:      Integer  from  Standard;
    pLongData:  Address  from  Standard;
    pFloatData: Address  from  Standard;
    pCharData:  Address  from  Standard)
  is private;


fields
  myBKIndex:          Integer   from Standard;
  myCurrentPage:      Integer   from Standard;
  myFileIsOpened:     Boolean   from Standard;
  myFillIndex:        Integer   from Standard; 
  myEdgeColor:        Integer   from Standard;
  myEdgeType:         Integer   from Standard;
  myEdgeWidth:        Integer   from Standard; 
  myInteriorStyle:    Integer   from Standard; 
  myEdgeVisibility:   Integer   from Standard;

end Driver from CGM;
