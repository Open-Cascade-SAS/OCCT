-- Created on: 1992-04-06
-- Created by: Christophe MARION
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class WiresBlock from HLRAlgo inherits TShared from MMgt

	---Purpose: A WiresBlock is a set of Blocks. It is used by the
	--          DataStructure to structure the Edges.
	--          
	--          A WiresBlock contains :
	--          
	--          * An Array  of Blocks.

uses
    Address           from Standard,
    Boolean           from Standard,
    Integer           from Standard,
    EdgesBlock        from HLRAlgo,
    Array1OfTransient from TColStd
    
is
    Create(NbWires : Integer from Standard)
	---Purpose: Create a Block of Blocks.
    returns mutable WiresBlock from HLRAlgo;

    NbWires(me) returns Integer from Standard
    is static;
    
    Set(me : mutable; I  : Integer     from Standard;
		      W  : EdgesBlock  from HLRAlgo)
    is static;		   

    Wire(me : mutable; I : Integer from Standard)
    returns any EdgesBlock from HLRAlgo
	---C++: return &
    is static;
    
    UpdateMinMax(me : mutable; TotMinMax : Address from Standard)
    is static;

    MinMax(me) returns Address from Standard
	---C++: inline
    is static;

fields
    myWires  : Array1OfTransient from TColStd;
    myMinMax : Integer           from Standard[16];

end WiresBlock;
