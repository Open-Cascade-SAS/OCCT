-- Created on: 1999-06-11
-- Created by: Sergey RUIN
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class UAttribute from TDataStd inherits Attribute from TDF


uses Attribute       from TDF,
     Label           from TDF,
     GUID            from Standard,
     DataSet         from TDF,
     RelocationTable from TDF

is    


    ---Purpose: api class methods
    --          =============
    
    Set (myclass ; label : Label from TDF; LocalID : GUID from Standard)
    ---Purpose: Find, or create, a UAttribute attribute with <LocalID> as Local GUID.
    -- The UAttribute attribute is returned.
    returns UAttribute from TDataStd ;    


    ---Purpose: UAttribute methods
    --          ============

    Create
    returns mutable UAttribute from TDataStd;
    
    SetID (me: mutable; LocalID : GUID from Standard);
    
    ID (me)
    ---C++: return const & 
    returns GUID from Standard;
    
    ---Category: methodes of TDF_Attribute
    --           =========================
 
    Restore (me: mutable; with : Attribute from TDF);

    NewEmpty (me)
    returns mutable Attribute from TDF;

    Paste (me; into : mutable Attribute from TDF;
	       RT   : mutable RelocationTable from TDF);       

    References (me; DS : DataSet from TDF) is redefined;   

    Dump(me; anOS : in out OStream from Standard)
    returns OStream from Standard
     is redefined;
	---C++: return &
fields
   
   myID:    GUID from Standard;
	
end UAttribute;
