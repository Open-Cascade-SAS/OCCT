-- Created on: 1992-09-28
-- Created by: Remi GILET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MakeRotation

from GCE2d

    	---Purpose: This class implements an elementary construction algorithm for
    	-- a rotation in 2D space. The result is a Geom2d_Transformation transformation.
    	-- A MakeRotation object provides a framework for:
    	-- -   defining the construction of the transformation,
    	-- -   implementing the construction algorithm, and
    	-- -   consulting the result.

uses Pnt2d          from gp,
     Transformation from Geom2d,
     Real           from Standard

is

Create(Point : Pnt2d  from gp      ;
       Angle : Real from Standard) returns MakeRotation;
    	---Purpose: Constructs a rotation through angle Angle about the center Point.
        
Value(me) returns Transformation from Geom2d
    is static;
      	---C++: return const&
      	---Purpose:  Returns the constructed transformation.

Operator(me) returns Transformation from Geom2d
    is static;
    	---C++: return const&
    	---C++: alias "Standard_EXPORT operator Handle_Geom2d_Transformation() const;"

fields

    TheRotation : Transformation from Geom2d;

end MakeRotation;


