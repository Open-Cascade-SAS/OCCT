-- Created on: 1993-01-09
-- Created by: CKY / Contract Toubro-Larsen ( TCD )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class LineFontPredefined from IGESGraph  inherits IGESEntity

        ---Purpose: defines IGESLineFontPredefined, Type <406> Form <19>
        --          in package IGESGraph
        --
        --          Provides the ability to specify a line font pattern
        --          from a predefined list rather than from
        --          Directory Entry Field 4

uses  Integer  -- no one specific type


is

        Create returns mutable LineFontPredefined;

        -- Specific Methods pertaining to the class

        Init (me                   : mutable;
              nbProps              : Integer;
              aLineFontPatternCode : Integer);
        ---Purpose : This method is used to set the fields of the class
        --           LineFontPredefined
        --       - nbProps              : Number of property values (NP = 1)
        --       - aLineFontPatternCode : Line Font Pattern Code

        -- Specific Access Methods : According to each type of Entity

        NbPropertyValues (me) returns Integer;
        ---Purpose : returns the number of property values in <me>

        LineFontPatternCode (me) returns Integer;
        ---Purpose : returns the Line Font Pattern Code of <me>

fields

--
-- Class    : IGESGraph_LineFontPredefined
--
-- Purpose  : Declaration of the variables specific to a
--            LineFontPredefined property.
--
-- Reminder : A LineFontPredefined property is defined by :
--                  - Number of property values
--                  - Line Font Pattern Code
--

        theNbPropertyValues    : Integer;

        theLineFontPatternCode : Integer;

end LineFontPredefined;
