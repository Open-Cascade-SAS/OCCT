-- File:	StepAP214_AppliedOrganizationAssignment.cdl
-- Created:	Wed Mar 10 10:16:54 1999
-- Author:	data exchange team
--		<det@androx.nnov.matra-dtv.fr>
---Copyright:	 Matra Datavision 1999


class AppliedOrganizationAssignment from StepAP214 
inherits OrganizationAssignment from StepBasic
       
uses
    	HArray1OfOrganizationItem from StepAP214, 
	OrganizationItem from StepAP214, 
	Organization from StepBasic,
	OrganizationRole from StepBasic


is
    
    Create returns mutable AppliedOrganizationAssignment;
	---Purpose: Returns a AppliedOrganizationAssignment


	Init (me : mutable;
	      aAssignedOrganization : mutable Organization from StepBasic;
	      aRole : mutable OrganizationRole from StepBasic) is redefined;

	Init (me : mutable;
	      aAssignedOrganization : mutable Organization from StepBasic;
	      aRole : mutable OrganizationRole from StepBasic;
	      aItems : mutable HArray1OfOrganizationItem from StepAP214) is virtual;

	-- Specific Methods for Field Data Access --

	SetItems(me : mutable; aItems : mutable HArray1OfOrganizationItem);
	Items (me) returns mutable HArray1OfOrganizationItem;
	ItemsValue (me; num : Integer) returns OrganizationItem;
	NbItems (me) returns Integer;
    
fields

    	items : HArray1OfOrganizationItem from StepAP214; -- a SelectType

end AppliedOrganizationAssignment;
