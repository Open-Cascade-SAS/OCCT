-- Created on: 2008-12-10
-- Created by: Pavel TELKOV
-- Copyright (c) 2008-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DimTol from PXCAFDoc inherits  Attribute from PDF

	---Purpose: 
uses
    Integer       from Standard,
    HAsciiString  from PCollection,
    HArray1OfReal from PColStd
is
    Create returns DimTol from PXCAFDoc;

    Create (theKind : Integer from Standard;
    	    theVal  : HArray1OfReal from PColStd;
    	    theName : HAsciiString from PCollection;
    	    theDescr: HAsciiString from PCollection)
    returns DimTol from PXCAFDoc;
    
    GetKind (me) returns Integer from Standard;

    GetVal (me) returns HArray1OfReal from PColStd;

    GetName (me) returns HAsciiString from PCollection;

    GetDescription (me) returns HAsciiString from PCollection;

    Set (me : mutable; theKind : Integer from Standard;
    	    	       theVal  : HArray1OfReal from PColStd;
    	    	       theName : HAsciiString from PCollection;
    	    	       theDescr: HAsciiString from PCollection);
    
fields

    myKind : Integer from Standard;
    myVal  : HArray1OfReal from PColStd;
    myName : HAsciiString from PCollection;
    myDescr: HAsciiString from PCollection;

end DimTol from PXCAFDoc;
