-- Created on: 2002-12-10
-- Created by: data exchange team
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V2.0

class SymmetricTensor23d from StepFEA
inherits SelectType from StepData

    ---Purpose: Representation of STEP SELECT type SymmetricTensor23d

uses
    SelectMember from StepData,
    HArray1OfReal from TColStd,
    HArray1OfReal from TColStd

is
    Create returns SymmetricTensor23d from StepFEA;
	---Purpose: Empty constructor

    CaseNum (me; ent: Transient) returns Integer;
	---Purpose: Recognizes a kind of SymmetricTensor23d select type
	--          return 0 

    CaseMem (me; ent: SelectMember from StepData) returns Integer is redefined;
	---Purpose: Recognizes a items of select member SymmetricTensor23dMember
	--          1 -> IsotropicSymmetricTensor23d
	--          2 -> OrthotropicSymmetricTensor23d
	--          3 -> AnisotropicSymmetricTensor23d
	--          0 else


     NewMember(me) returns SelectMember from StepData is redefined;
	---Purpose: Returns a new select member the type SymmetricTensor23dMember

    SetIsotropicSymmetricTensor23d(me: in out; aVal :Real);
	---Purpose: Set Value for IsotropicSymmetricTensor23d

    IsotropicSymmetricTensor23d (me) returns Real;
	---Purpose: Returns Value as IsotropicSymmetricTensor23d (or Null if another type)

    SetOrthotropicSymmetricTensor23d(me: in out; aVal :HArray1OfReal from TColStd);
	---Purpose: Set Value for OrthotropicSymmetricTensor23d

    OrthotropicSymmetricTensor23d (me) returns HArray1OfReal from TColStd;
	---Purpose: Returns Value as OrthotropicSymmetricTensor23d (or Null if another type)

    SetAnisotropicSymmetricTensor23d(me: in out; aVal :HArray1OfReal from TColStd);
	---Purpose: Set Value for AnisotropicSymmetricTensor23d

    AnisotropicSymmetricTensor23d (me) returns HArray1OfReal from TColStd;
	---Purpose: Returns Value as AnisotropicSymmetricTensor23d (or Null if another type)

end SymmetricTensor23d;
