-- Created by: NW,JPB,CAL
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class AspectLine3d from Graphic3d inherits AspectLine from Aspect

	---Version:

	---Purpose: Creates and updates a group of attributes
	--	    for 3d line primitives. This group contains the
	--	    colour, the type of line, and its thickness.
	

uses

	Color          from Quantity,
	TypeOfLine     from Aspect,
	ShaderProgram  from Graphic3d

is

	Create
		returns AspectLine3d from Graphic3d;
	---Level: Public
	---Purpose: Creates a context table for line primitives
	--	    defined with the following default values:
	--
	--	    Colour	: NOC_YELLOW
	--	    Line type	: TOL_SOLID
	--	    Width	: 1.0

	Create ( AColor	: Color from Quantity;
		 AType	: TypeOfLine from Aspect;
		 AWidth	: Real from Standard )
		returns AspectLine3d from Graphic3d;
	---Level: Public
	---Purpose: Creates a context table for line primitives
	--	    defined with the specified values.
	--  Warning: <AWidth> is the "linewidth scale factor".
	--	    The nominal line width is 1 pixel. The width of
	--	    the line is determined by applying the linewidth scale
	--	    factor to this nominal line width.
	--	    The supported linewidths vary by 1-pixel units.

  SetShaderProgram ( me  :  mutable; 
                     theProgram  :  ShaderProgram from Graphic3d );
  ---Level: Public
  ---Purpose: Sets up OpenGL/GLSL shader program.

  ShaderProgram ( me )
  returns ShaderProgram from Graphic3d;
  ---C++: return const &

fields

--
-- Class	:	Graphic3d_AspectLine3d
--
-- Purpose	:	Declaration of context-specific variables
--			for drawing 3d lines
--
-- Reminder	:	A context for drawing 3d lines inherits:
--			- the colour
--			- the type of line
--			- the thickness
--			defined by AspectLine.
--

  MyShaderProgram  :  ShaderProgram  from  Graphic3d; 

end AspectLine3d;
