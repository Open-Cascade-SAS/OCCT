-- Created on: 1993-07-27
-- Created by: Jean Louis FRENKEL
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


package ImageUtility


uses
	TCollection,
	Image,
	AlienImage,
	OSD,
	Aspect

is

	class XPR ;
		--- Purpose : perform a "xpr " with a XAlienImage build
		-- 		 from any Image , any AlienImage .

	class XWUD ;
		--- Purpose : perform a "xwud " with a XAlienImage build
		-- 		 from any Image , any AlienImage .

	class XWD ;
		--- Purpose : perform a "xwd " and create Image and XAlienImage.

	class X11Dump ;
		--- Purpose : Create a X11 Window and perform a XPutImage on it,
		--            from any Image , any AlienImage .

	imported X11Window ;
		--- Xlib.h : Window type

	imported X11Display ;
		--- Xlib.h : Display type

	imported X11XImage ;
		--- Xlib.h : XImage type

	imported X11GC ;
		--- Xlib.h : XImage type

	PixelDiff( aImage       : immutable Image from Image ;
	           anotherImage : immutable Image from Image ) 
		returns mutable PseudoColorImage from Image
		--- Purpose : Create a Black & White Image from two Image.
		--	      Resulting Image Pixel is set to 0 if Pixel from
		--	      both Image are the same else set to 1 .
		raises TypeMismatch from Standard;

	PixelColorDiff( aImage       : immutable Image from Image ;
	                anotherImage : immutable Image from Image ) 
		returns mutable PseudoColorImage from Image
		--- Purpose : Create a Black & White Image from two Image.
		--	      Resulting Image Pixel is set to 0 if PixelColor 
		--	      from both Image are the same else set to 1 .
		raises TypeMismatch from Standard;

	PixelColorDiff( aImage       : immutable Image from Image ;
	                anotherImage : immutable Image from Image ;
			aCRColorMap  : immutable ColorRampColorMap from Aspect )
		returns mutable PseudoColorImage from Image
		--- Purpose : Create a ColorRamp Image from two Image.
		--	      Resulting Image Pixel Index is proportional
		--	      to the (Red+Green_Blue)Image Differences scaling
		--	      to the ColorRamp range.
		raises TypeMismatch from Standard;

	PixelColorDiff( aImage       : immutable Image from Image ;
	                anotherImage : immutable Image from Image ;
			aCRColorMap  : immutable ColorRampColorMap from Aspect ;
			RedDiff      : out mutable PseudoColorImage from Image ;
			GreenDiff    : out mutable PseudoColorImage from Image ;
			BlueDiff     : out mutable PseudoColorImage from Image )
		--- Purpose : Create a ColorRamp Images from two Image.
		--	      Resulting Image Pixel Index is proportional
		--	      to the Image Differences scaling to the 
		--	      ColorRamp range.
		raises TypeMismatch from Standard;


end ;
