-- Created on: 1991-12-06
-- Created by: Remi LEQUETTE
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


package HLRTest 

	---Purpose: This package   is  a test  of  the    Hidden Lines
	--          algorithms instantiated on the BRep Data Structure
	--          and using the Draw package to display the results.

uses
    Standard,
    MMgt,
    TCollection,
    gp,
    TopoDS,
    HLRAlgo,
    HLRBRep,
    HLRTopoBRep,
    Draw

is
    class ShapeData;
    
    class DrawableEdgeTool;
	---Purpose: Used to display the results.

    class DrawablePolyEdgeTool;
	---Purpose: Used to display the results.

    class Projector;
	---Purpose: Draw Variable Projector to test
	
    class OutLiner;
	---Purpose: Draw Variable Outliner to test

    Set(Name : CString;
        P    : Projector from HLRAlgo);
	---Purpose: Set a Projector Variable

    GetProjector(Name : in out CString;
                 P :    in out Projector from HLRAlgo) 
    returns Boolean; 
	---Purpose: Get a projector variable
	--          Returns false if the variable is not a projector

    Set(Name : CString;
        S    : Shape from TopoDS);
	---Purpose: Set a OutLiner Variable

    GetOutLiner(Name : in out CString)  
    	returns OutLiner from HLRTopoBRep;
	---Purpose: Get a outliner variable
	--          Returns a null handle if the variable is not a outliner

    Commands(I : in out Interpretor from Draw);
	---Purpose: Defines commands to test the Hidden Line Removal

end HLRTest;
