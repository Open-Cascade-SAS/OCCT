-- Created on: 1998-08-04
-- Created by: Christian CAILLET
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class AutoDesignOrganizationItem  from StepAP214    
    inherits AutoDesignGeneralOrgItem  from StepAP214

    -- adds : document,  physically_modelled_product_definition

uses
    Document from StepBasic,
    PhysicallyModeledProductDefinition from StepBasic

is

    Create returns AutoDesignOrganizationItem;

    CaseNum (me; ent : Transient) returns Integer  is redefined;
    -- adds : 9  Document
    --       10  PhysicallyModeledProductDefinition

    Document (me) returns Document;

    PhysicallyModeledProductDefinition (me) returns PhysicallyModeledProductDefinition;

end AutoDesignOrganizationItem;
