-- Created on: 2001-05-03
-- Created by: Igor FEOKTISTOV
-- Copyright (c) 2001-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Limitation from QANewModTopOpe inherits MakeShape from BRepBuilderAPI

---Purpose: provides  cutting  shape  by  face  or  shell;

uses

    Shape from TopoDS, 
    ListOfShape from TopTools, 
    ModeOfLimitation  from  QANewModTopOpe, 
    State  from  TopAbs,  
    CutPtr  from  QANewModTopOpe, 
    CommonPtr  from  QANewModTopOpe
is 
  
    Create(theObjectToCut,  theCutTool : Shape from TopoDS;
    	    theMode : ModeOfLimitation  from  QANewModTopOpe = QANewModTopOpe_Forward)
    ---Purpose: initializes and  fills data structure for  cutting and
    --          makes  cutting according to orientation theCutTool and
    --          theMode.
    --          if theCutTool is not face or shell does nothing.
    
    returns Limitation from QANewModTopOpe;    
     
    Cut(me  :  in  out);
    ---Purpose: makes cutting  according to  orientation theCutTool
    --          and  current value   of  myMode.  Does nothing  if
    --          result already  exists.

    SetMode(me  :  in  out;  theMode  :  ModeOfLimitation  from  QANewModTopOpe); 
     
    GetMode(me)  returns  ModeOfLimitation  from  QANewModTopOpe;  
     
    Shape1(me)  returns  Shape  from  TopoDS
    ---Purpose: Returns the first shape.
    ---C++: return const &
    ---Level: Public
    is static;
     
    Shape2(me)  returns  Shape  from  TopoDS
    ---Purpose: Returns the second shape.
    ---C++: return const &
    ---Level: Public
    is static; 
    
    Modified (me: in out; S : Shape from TopoDS)
    	---Purpose: Returns the list  of shapes modified from the shape
    	--          <S>. 
        ---C++: return const & 
        ---Level: Public
    returns ListOfShape from TopTools
    is redefined;

    Generated (me: in out; S : Shape from TopoDS)
    	returns ListOfShape from TopTools
	is redefined;
    	---Purpose: Returns the list  of shapes generated from the shape <S>.
    	---         For use in BRepNaming.
    	---C++:  return const &
    
    HasModified (me)
    	returns Boolean from Standard
	is virtual;
    	---Purpose: Returns true if there is at least one modified shape.
    	---         For use in BRepNaming.

    HasGenerated (me)
    	returns Boolean from Standard
	is virtual;
    	---Purpose: Returns true if there is at least one generated shape.
    	---         For use in BRepNaming.

    HasDeleted (me)
    	returns Boolean from Standard
	is virtual;
    	---Purpose: Returns true if there is at least one deleted shape.
    	---         For use in BRepNaming.

    IsDeleted (me: in out; S : Shape from TopoDS)
    returns Boolean from Standard
    is redefined;
      
    Delete(me  :  in  out)  is  redefined; 
    ---C++:  alias  "Standard_EXPORT  ~QANewModTopOpe_Limitation()  {Delete();}"
  

fields 

    myResultFwd     :  Shape  from  TopoDS;  
    myResultRvs     :  Shape  from  TopoDS;  
    myObjectToCut   :  Shape  from  TopoDS;  
    myCutTool       :  Shape  from  TopoDS;  
    myCut           :  CutPtr  from  QANewModTopOpe;
    myCommon        :  CommonPtr  from  QANewModTopOpe;
    myFwdIsDone     :  Boolean  from  Standard;
    myRevIsDone     :  Boolean  from  Standard;  
    myMode          :  ModeOfLimitation  from  QANewModTopOpe;
    
end  Limitation;
