-- Created on: 1995-07-24
-- Created by: Modelistation
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class WFPoleSurface from StdPrs

inherits Root from Prs3d
    	--- Purpose: The number of lines to be drawn is controlled 
    	-- by the NetworkNumber of the given Drawer.
uses
    Surface      from Adaptor3d,
    Presentation from Prs3d,
    Drawer       from Prs3d
    	

is
   
 
    Add(myclass; aPresentation: Presentation from Prs3d;  
    	    	 aSurface     : Surface      from Adaptor3d;
    	    	 aDrawer      : Drawer       from Prs3d);
    	---Purpose: Adds the surface aSurface to the presentation object aPresentation.
    	-- The shape's display attributes are set in the attribute manager aDrawer.
    	-- The surface aSurface is a surface object from
    	-- Adaptor3d, and provides data from a Geom surface.
    	-- This makes it possible to use the surface in a geometric algorithm.
end WFPoleSurface;



