-- Created on: 1992-02-03
-- Created by: Christian CAILLET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



package Transfer

    ---Purpose : Defines general Transfer engine, which provides tools and
    --           workframe for all kinds of file (non-direct) Interfaces.
    --           Works on the basis of data provided by package Interface
    --           (especially InterfaceModel).

uses TCollection, TColStd, MMgt, Standard, Dico, MoniTool, Interface,  Message

is

    class DataInfo;  -- used in Mapper

    deferred class Finder;
    	generic class Mapper;
	class TransientMapper  instantiates Mapper
    	    (Transient, MapTransientHasher from TColStd, DataInfo);
    class FindHasher;

    deferred class Binder;
    	class VoidBinder;
    	generic class SimpleBinder;
    	class SimpleBinderOfTransient;
	class BinderOfTransientInteger;
        class TransientListBinder;
    	class MultipleBinder;

    class ResultFromTransient;
    class ResultFromModel;

    class TransferIterator;
    generic class TransferProcess;
    generic class TransferMap;
    generic class Iterator;
    generic class Actor;

    class ProcessForTransient   instantiates TransferProcess
    	(Transient,  MapTransientHasher from TColStd,
    	 HSequenceOfTransient  from TColStd);
    ---Purpose : Manages Transfer of Transient Objects. Produces also
    --           ActorOfTransientProcess       (deferred class),
    --           IteratorOfTransientProcess    (for Results),
    --           TransferMapOfTransientProcess (internally used)
    --           Normally uses as TransientProcess, which adds some specifics

    class TransientProcess;    -- inherits TransferForTransient
    class ActorOfTransientProcess;

    class SequenceOfFinder instantiates
    	 Sequence from TCollection (Finder);
    class HSequenceOfFinder instantiates
    	HSequence from TCollection (Finder,SequenceOfFinder);

    class ProcessForFinder      instantiates TransferProcess
    	(Finder,     FindHasher,   HSequenceOfFinder);

    class FinderProcess;
    class ActorOfFinderProcess;

    class TransferOutput;
    class TransferInput;

    class DispatchControl;
    class TransferDispatch;
    class ActorDispatch;
    
    class MapContainer;

    class SequenceOfBinder instantiates
    	 Sequence from TCollection (Binder);
    class HSequenceOfBinder instantiates
    	HSequence from TCollection (Binder,SequenceOfBinder);

    enumeration StatusResult is  StatusVoid, StatusDefined, StatusUsed;
    ---Purpose : result status of transferring an entity (see Transcriptor)

    enumeration StatusExec is
    	StatusInitial, StatusRun, StatusDone, StatusError,StatusLoop;
    ---Purpose : execution status of an individual transfer (see Transcriptor)

    enumeration UndefMode is
    	UndefIgnore, UndefFailure, UndefContent, UndefUser;
    ---Purpose : used on processing Undefined Entities (see TransferOutput)

    	-- --  Exceptions  -- --

    exception TransferFailure   inherits InterfaceError  from Interface;
    exception TransferDeadLoop  inherits TransferFailure from Transfer;

end Transfer;
