-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class TextLiteral from StepVisual 

inherits GeometricRepresentationItem from StepGeom

uses

	HAsciiString from TCollection, 
	Axis2Placement from StepGeom, 
	TextPath from StepVisual, 
	FontSelect from StepVisual
is

	Create returns mutable TextLiteral;
	---Purpose: Returns a TextLiteral


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aLiteral : mutable HAsciiString from TCollection;
	      aPlacement : Axis2Placement from StepGeom;
	      aAlignment : mutable HAsciiString from TCollection;
	      aPath : TextPath from StepVisual;
	      aFont : FontSelect from StepVisual) is virtual;

	-- Specific Methods for Field Data Access --

	SetLiteral(me : mutable; aLiteral : mutable HAsciiString);
	Literal (me) returns mutable HAsciiString;
	SetPlacement(me : mutable; aPlacement : Axis2Placement);
	Placement (me) returns Axis2Placement;
	SetAlignment(me : mutable; aAlignment : mutable HAsciiString);
	Alignment (me) returns mutable HAsciiString;
	SetPath(me : mutable; aPath : TextPath);
	Path (me) returns TextPath;
	SetFont(me : mutable; aFont : FontSelect);
	Font (me) returns FontSelect;

fields

	literal : HAsciiString from TCollection;
	placement : Axis2Placement from StepGeom; -- a SelectType
	alignment : HAsciiString from TCollection;
	path : TextPath from StepVisual; -- an Enumeration
	font : FontSelect from StepVisual; -- a SelectType

end TextLiteral;
