-- Created on: 1997-10-01
-- Created by: Christian CAILLET
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class SelectFaces  from IGESSelect  inherits SelectExplore

    ---Purpose : This selection returns the faces contained in an IGES Entity
    --           or itself if it is a Face
    --           Face means :
    --           - Face (510) of a ManifoldSolidBrep
    --           - TrimmedSurface (144)
    --           - BoundedSurface (143)
    --           - Plane with a Bounding Curve (108, form not 0)
    --           - Also, any Surface which is not in a TrimmedSurface, a
    --             BoundedSurface, or a Face (FREE Surface)
    --           -> i.e. a Face for which Natural Bounds will be considered

uses AsciiString from TCollection, Transient, EntityIterator, Graph

is


    Create returns mutable  SelectFaces;


    Explore (me; level : Integer; ent : Transient; G : Graph;
    	     explored : in out EntityIterator)
    	returns Boolean;
    ---Purpose : Explores an entity, to take its faces
    --           Works recursively


    ExploreLabel (me) returns AsciiString from TCollection;
    ---Purpose : Returns a text defining the criterium : "Faces"

end SelectFaces;
