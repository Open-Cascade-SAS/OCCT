-- Created on: 1992-08-24
-- Created by: Ramin BARRETO
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class Transient from Standard 

    ---Purpose: Abstract class which forms the root of the entire 
    --          Transient class hierarchy.
    ---Warning: This CDL file is actually a stub, even if it attempts to be correct. 
    --          See actual header in Standard_Transient_proto.hxx

uses
    Type from Standard,
    Boolean from Standard,
    Integer from Standard
    
is

        Initialize;
    	    ---Purpose: Empty constructor
	    ---Warning: Copy constructor and assignment operators cannot be 
	    --          declared cleanly in CDL, so we use "C++ alias" for that
    	    ---C++: alias "Standard_Transient(const Standard_Transient&) : count(0) {}"
    	    ---C++: alias "Standard_Transient& operator= (const Standard_Transient&) { return *this; }"

	HashCode (me; Upper : Integer ) returns Integer is virtual;
	    ---Purpose: Returns a hashed value denoting <me>. This value is in
	    --         the range 1..<Upper>.
	    ---C++:  function call
	    ---Level: Advanced

        Delete(me) is  virtual;
            ---Purpose: Memory deallocator for transient classes
            ---Level: Advanced
    	    ---C++: alias "Standard_EXPORT virtual ~Standard_Transient();"
            
	DynamicType (me) returns Type is virtual;
            ---Purpose: Returns a type information object about this object.
            ---Level: Advanced
            
	IsInstance (me; TheType : Type) returns Boolean is static;
            ---Purpose: Returns a true value if this is an instance of Type.
            ---Level: Advanced
            
	IsInstance (me; TheTypeName : CString) returns Boolean is static;
            ---Purpose: Returns a true value if this is an instance of TypeName.
            ---Level: Advanced
            
	IsKind (me; TheType : Type) returns Boolean is static;
	    ---Purpose: Returns true if this is an instance of Type or an
	    --          instance of any class that inherits from Type.
	    --          Note that multiple inheritance is not supported by OCCT RTTI mechanism.
	    ---Level: Advanced
	    
	IsKind (me; TheTypeName : CString) returns Boolean is static;
	    ---Purpose: Returns true if this is an instance of TypeName or an
	    --         instance of any class that inherits from TypeName.
	    --          Note that multiple inheritance is not supported by OCCT RTTI mechanism.
	    ---Level: Advanced
	    
	This (me) returns mutable Transient
	    ---Purpose: Returns a Handle which references this object.
	    ---Warning: Must never be called to objects created in stack.
	    ---Level: Advanced
	is virtual protected;
 
 ---Level: Advanced 

        GetRefCount(me) 
	    ---Purpose: get the reference counter
	    --          of this object.
	    returns  Integer  from  Standard; 

     fields
        count : Integer from Standard;
	
end Transient from Standard;



