-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PlanarExtent from StepVisual 

inherits GeometricRepresentationItem from StepGeom

uses

	Real from Standard, 
	HAsciiString from TCollection
is

	Create returns PlanarExtent;
	---Purpose: Returns a PlanarExtent


	Init (me : mutable;
	      aName : HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      aName : HAsciiString from TCollection;
	      aSizeInX : Real from Standard;
	      aSizeInY : Real from Standard) is virtual;

	-- Specific Methods for Field Data Access --

	SetSizeInX(me : mutable; aSizeInX : Real);
	SizeInX (me) returns Real;
	SetSizeInY(me : mutable; aSizeInY : Real);
	SizeInY (me) returns Real;

fields

	sizeInX : Real from Standard;
	sizeInY : Real from Standard;

end PlanarExtent;
