-- Created on: 1995-09-21
-- Created by: Bruno DUMORTIER
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

private class ApproxSeewing from BRepFill 

	---Purpose: Evaluate the 3dCurve  and the PCurves described in
	--          a MultiLine from BRepFill.  The parametrization of
	--          those curves is  not  imposed by  the Bissectrice.
	--          The  parametrization  is given  approximatively by
	--          the abscissa of the curve3d. 

uses

    MultiLine from BRepFill,
    Curve from Geom,
    Curve from Geom2d
    
raises

    NotDone from StdFail
    
is
    Create returns ApproxSeewing from BRepFill;
    
    Create( ML : MultiLine from BRepFill) 
    returns ApproxSeewing from BRepFill;
    
    Perform(me : in out;
    	    ML : MultiLine from BRepFill)
    is static;
    
    IsDone(me) 
    returns Boolean from Standard
    is static;
    
    Curve(me) 
    	---Purpose: returns the approximation of the 3d Curve
	---C++: return const &
    returns Curve from Geom
    raises
    	NotDone from StdFail
    is static;
    
    CurveOnF1(me) 
    	---Purpose: returns the  approximation  of the  PCurve  on the
    	--          first face of the MultiLine
	---C++: return const &
    returns Curve from Geom2d
    raises
    	NotDone from StdFail
    is static;
    
    CurveOnF2(me) 
    	---Purpose: returns the  approximation  of the  PCurve  on the
    	--          first face of the MultiLine
	---C++: return const &
    returns Curve from Geom2d
    raises
    	NotDone from StdFail
    is static;
    
fields
    myML      : MultiLine from BRepFill;
    myIsDone  : Boolean   from Standard;
    myCurve   : Curve     from Geom;
    myPCurve1 : Curve     from Geom2d;
    myPCurve2 : Curve     from Geom2d;

end ApproxSeewing;
