-- Created on: 1993-02-22
-- Created by: Philippe DAUTRY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Circle from PGeom inherits Conic from PGeom

        ---Purpose : Defines a circle in 3D space.
        --         
	---See Also : Circle from Geom.

uses Ax2 from gp

is


  Create returns mutable Circle from PGeom;
	---Purpose : Creates a circle with default values.
    	---Level: Internal 


  Create (aPosition : Ax2 from gp; aRadius : Real from Standard)
    returns mutable Circle from PGeom;
        ---Purpose : Creates a Circle with <aPosition> and <aRadius> as field
        --         values.
    	---Level: Internal 


  Radius (me : mutable; aRadius : Real from Standard);
	---Purpose: Set the value of the field radius with <aRadius>.
    	---Level: Internal 


  Radius (me) returns Real from Standard;
	---Purpose: Returns the value of the field radius.
    	---Level: Internal 


fields

  radius : Real from Standard;

end;

