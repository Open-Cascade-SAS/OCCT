-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DimensionalExponents from StepBasic 

inherits TShared from MMgt

uses

	Real from Standard
is

	Create returns DimensionalExponents;
	---Purpose: Returns a DimensionalExponents

	Init (me : mutable;
	      aLengthExponent : Real from Standard;
	      aMassExponent : Real from Standard;
	      aTimeExponent : Real from Standard;
	      aElectricCurrentExponent : Real from Standard;
	      aThermodynamicTemperatureExponent : Real from Standard;
	      aAmountOfSubstanceExponent : Real from Standard;
	      aLuminousIntensityExponent : Real from Standard) is virtual;

	-- Specific Methods for Field Data Access --

	SetLengthExponent(me : mutable; aLengthExponent : Real);
	LengthExponent (me) returns Real;
	SetMassExponent(me : mutable; aMassExponent : Real);
	MassExponent (me) returns Real;
	SetTimeExponent(me : mutable; aTimeExponent : Real);
	TimeExponent (me) returns Real;
	SetElectricCurrentExponent(me : mutable; aElectricCurrentExponent : Real);
	ElectricCurrentExponent (me) returns Real;
	SetThermodynamicTemperatureExponent(me : mutable; aThermodynamicTemperatureExponent : Real);
	ThermodynamicTemperatureExponent (me) returns Real;
	SetAmountOfSubstanceExponent(me : mutable; aAmountOfSubstanceExponent : Real);
	AmountOfSubstanceExponent (me) returns Real;
	SetLuminousIntensityExponent(me : mutable; aLuminousIntensityExponent : Real);
	LuminousIntensityExponent (me) returns Real;

fields

	lengthExponent : Real from Standard;
	massExponent : Real from Standard;
	timeExponent : Real from Standard;
	electricCurrentExponent : Real from Standard;
	thermodynamicTemperatureExponent : Real from Standard;
	amountOfSubstanceExponent : Real from Standard;
	luminousIntensityExponent : Real from Standard;

end DimensionalExponents;
