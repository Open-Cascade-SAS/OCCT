-- Created on: 2002-12-12
-- Created by: data exchange team
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class ParametricSurface3dElementCoordinateSystem from StepFEA
inherits FeaRepresentationItem from StepFEA

    ---Purpose: Representation of STEP entity ParametricSurface3dElementCoordinateSystem

uses
    HAsciiString from TCollection

is
    Create returns ParametricSurface3dElementCoordinateSystem from StepFEA;
	---Purpose: Empty constructor

    Init (me: mutable; aRepresentationItem_Name: HAsciiString from TCollection;
                       aAxis: Integer;
                       aAngle: Real);
	---Purpose: Initialize all fields (own and inherited)

    Axis (me) returns Integer;
	---Purpose: Returns field Axis
    SetAxis (me: mutable; Axis: Integer);
	---Purpose: Set field Axis

    Angle (me) returns Real;
	---Purpose: Returns field Angle
    SetAngle (me: mutable; Angle: Real);
	---Purpose: Set field Angle

fields
    theAxis: Integer;
    theAngle: Real;

end ParametricSurface3dElementCoordinateSystem;
