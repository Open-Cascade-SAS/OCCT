-- Created on: 1996-12-03
-- Created by: Arnaud BOUZY/Odile Olivier
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class LengthDimension from AIS inherits Relation from AIS

	---Purpose: A framework to display lengths.
    	-- These can be lengths along a face or edge, or
    	-- between two faces or two edges.
    	-- The value of the length is given in a text figuring in this display.

uses Shape                 from TopoDS,
     Face                  from TopoDS,
     Presentation          from Prs3d,
     PresentationManager3d from PrsMgr,
     Selection             from SelectMgr,
     Dir                   from gp,
     Pnt                   from gp,
     Projector             from Prs3d,
    Transformation        from Geom,
     PresentationManager2d from PrsMgr,
     GraphicObject         from Graphic2d,
     ExtendedString        from TCollection,
     Plane                 from Geom,
     TypeOfDist            from AIS,
     ArrowSide             from DsgPrs,
     KindOfDimension       from AIS,
     Drawer                from Prs3d,
     Edge                  from TopoDS,
     Box                   from Bnd,
     Drawer                from AIS,
     Vertex                from TopoDS
is



    Create (aFirstFace  : Face           from TopoDS;
    	    aSecondFace : Face           from TopoDS;
	    aVal        : Real           from Standard; -- is defined while first compute, may be any Real
	    aText       : ExtendedString from TCollection)    
	    ---Purpose: Constructs a length display object defined by the first
    	    -- face aFShape, the second face aSShape, the dimension aVal, and the text aText.
        
    returns mutable LengthDimension from AIS;

    Create (aFirstFace  : Face           from TopoDS;
    	    aSecondFace : Face           from TopoDS;
	    aVal        : Real           from Standard; -- is defined while first compute, may be any Real
	    aText       : ExtendedString from TCollection;    
	    aPosition   : Pnt            from gp;
	    aSymbolPrs  : ArrowSide      from DsgPrs;    
    	    anArrowSize : Real           from Standard = 0.0)
	    ---Purpose: Constructs a length display object defined by the first
    	    -- face aFShape, the second face aSShape, the
    	    -- dimension aVal, the position aPosition, the arrow
    	    -- aSymbolPrs with the size anArrowSize and the text aText.
    returns mutable LengthDimension from AIS;

    Create (Face      : Face           from TopoDS;
    	    Edge      : Edge           from TopoDS;
	    Val       : Real           from Standard;
	    Text      : ExtendedString from TCollection)
	    ---Purpose: Constructs a length display object defined by the first
    	    -- edge or vertex aFShape, the second edge or vertex
    	    -- aSShape, the dimension aVal,and the plane aPlane.
    returns mutable LengthDimension from AIS;
     
    Create (aFShape     : Shape          from TopoDS;
    	    aSShape     : Shape          from TopoDS;
            aPlane      : Plane          from Geom;
	    aVal        : Real           from Standard;
	    aText       : ExtendedString from TCollection)  
	    ---Purpose: -- Constructs a length display object defined by the first
    	    -- edge or vertex aFShape, the second edge or vertex
    	    -- aSShape, the dimension aVal,and the plane aPlane.
    returns mutable LengthDimension from AIS;

    Create (aFShape     : Shape          from TopoDS;
    	    aSShape     : Shape          from TopoDS;
            aPlane      : Plane          from Geom;
	    aVal        : Real           from Standard;
	    aText       : ExtendedString from TCollection;    
	    aPosition   : Pnt            from gp;
	    aSymbolPrs  : ArrowSide      from DsgPrs;    
	    aTypeDist   : TypeOfDist     from AIS;    
    	    anArrowSize : Real           from Standard = 0.0)
	    ---Purpose: Constructs a length display object defined by the first
    	    -- edge or vertex aFShape, the second edge or vertex
    	    -- aSShape, the dimension aVal, the position aPosition,
    	    -- the type of distance aTypeDist, the type of arrow
    	    -- aSymbolPrs with the size anArrowSize, and the plane aPlane.
    returns mutable LengthDimension from AIS;

    SetFirstShape( me: mutable; aFShape : Shape from TopoDS )
    is redefined static;

    SetSecondShape( me: mutable; aSShape : Shape from TopoDS )
    is redefined static;

    KindOfDimension(me) 
    returns KindOfDimension from AIS 
    is redefined;
    	    ---Purpose: Indicates that we are concerned with a length.
        
    IsMovable(me) returns Boolean from Standard 
    is redefined;    
    	    ---Purpose: Returns true if the length dimension is movable.
   
     TypeOfDist (me) 
            ---C++: inline   
    	    --- Purpose:
    	    -- Returns the type of distance of the length primitive.
    returns TypeOfDist from AIS
    is static;

    SetTypeOfDist(me: mutable;aTypeDist: TypeOfDist from AIS)
	    ---C++: inline       
	    --- Purpose:
    	    -- Returns true if the length dimension is movable.
    is static;

     
    	-- Methods from PresentableObject

    Compute(me : mutable;
    	    aPresentationManager :         PresentationManager3d from PrsMgr;
    	    aPresentation        : mutable Presentation          from Prs3d;
    	    aMode                :         Integer               from Standard= 0) 
    is redefined private;
    
    Compute(me : mutable;
    	    aProjector    :         Projector    from Prs3d;
            aPresentation : mutable Presentation from Prs3d)
    is redefined static private;     

    Compute(me:mutable;
    	    aPresentationManager: PresentationManager2d from PrsMgr;
            aPresentation: mutable GraphicObject from Graphic2d;
            aMode: Integer from Standard = 0)
    is redefined static private;

    Compute(me            : mutable;
    	    aProjector    : Projector from Prs3d;
    	    aTrsf         : Transformation from Geom;
	    aPresentation : mutable Presentation from Prs3d)
    is redefined;
    	---Purpose: computes the presentation according to a point of view
    	--          given by <aProjector>. 
    	--          To be Used when the associated degenerated Presentations 
    	--          have been transformed by <aTrsf> which is not a Pure
    	--          Translation. The HLR Prs can't be deducted automatically
    	--          WARNING :<aTrsf> must be applied
    	--           to the object to display before computation  !!!


    	-- Methods from SelectableObject

    ComputeSelection(me : mutable;
    	    	     aSelection : mutable Selection from SelectMgr;
    	    	     aMode      :         Integer   from Standard)
    is redefined private;



    	--     Computation private methods

    ComputeOneFaceLength(me : mutable; 
    	    	    	 aPresentation : mutable Presentation from Prs3d)
    is private;
    
    ComputeOneEdgeLength(me : mutable;
    	    	    	 aPresentation : mutable Presentation from Prs3d)
    is private;
    
    ComputeTwoFacesLength(me: mutable;
    	    	    	  aPresentation : mutable Presentation from Prs3d)
    is private;
    

    ComputeEdgeFaceLength (me: mutable;
    	    	    	   aPresentation : mutable Presentation from Prs3d)
    is private;


    ComputeTwoEdgesLength (myclass;
    	    	    	   aPresentation : mutable Presentation   from Prs3d; 
			   aDrawer       :         Drawer         from AIS; 
			   aText         :         ExtendedString from TCollection; 
			   ArrowSize     :         Real           from Standard;
			   FirstEdge     :         Edge           from TopoDS;
			   SecondEdge    :         Edge           from TopoDS;
			   Plane         :         Plane          from Geom;
			   AutomaticPos  :         Boolean        from Standard;
			   IsSetBndBox   :         Boolean        from Standard;
			   BndBox        :         Box            from Bnd;
			   ExtShape      : out     Integer        from Standard;
			   Val           : out     Real           from Standard;
			   DirAttach     : out     Dir            from gp;
			   Position      : out     Pnt            from gp;
			   FirstAttach   : out     Pnt            from gp;
			   SecondAttach  : out     Pnt            from gp;
			   SymbolPrs     : out     ArrowSide      from DsgPrs );
    
    ComputeOneEdgeOneVertexLength(myclass; 
    	    	    	          aPresentation : mutable Presentation   from Prs3d;
			          aDrawer       :         Drawer         from AIS; 
			          aText         :         ExtendedString from TCollection; 
			          ArrowSize     :         Real           from Standard;
			          FirstShape    :         Shape          from TopoDS;
			          SecondShape   :         Shape          from TopoDS;
			          Plane         :         Plane          from Geom;
			          AutomaticPos  :         Boolean        from Standard;
			          IsSetBndBox   :         Boolean        from Standard;
			          BndBox        :         Box            from Bnd;
			          ExtShape      : out     Integer        from Standard;
			          Val           : out     Real           from Standard;
			          DirAttach     : out     Dir            from gp;
			          Position      : out     Pnt            from gp;
			          FirstAttach   : out     Pnt            from gp;
			          SecondAttach  : out     Pnt            from gp;
			          SymbolPrs     : out     ArrowSide      from DsgPrs );
    
    ComputeTwoVerticesLength(myclass; 
    	    	    	     aPresentation : mutable Presentation   from Prs3d;
			     aDrawer       :         Drawer         from AIS; 
			     aText         :         ExtendedString from TCollection; 
			     ArrowSize     :         Real           from Standard;
			     FirstVertex   :         Vertex         from TopoDS;
			     SecondVertex  :         Vertex         from TopoDS;
			     Plane         :         Plane          from Geom;
			     AutomaticPos  :         Boolean        from Standard;
			     IsSetBndBox   :         Boolean        from Standard;
			     BndBox        :         Box            from Bnd;
			     TypeDist      :         TypeOfDist     from AIS;
			     ExtShape      : out     Integer        from Standard;
			     Val           : out     Real           from Standard;
			     DirAttach     : out     Dir            from gp;
			     Position      : out     Pnt            from gp;
			     FirstAttach   : out     Pnt            from gp;
			     SecondAttach  : out     Pnt            from gp;
			     SymbolPrs     : out     ArrowSide      from DsgPrs );

    
--
--      Computation Selection private methods
--      

    ComputeFaceSelection(me         : mutable;
    	    	         aSelection : mutable Selection from SelectMgr) 
    is private;
    
    ComputeEdgeVertexSelection( me         : mutable;
    	    	     	        aSelection : mutable Selection from SelectMgr) 
    is private;
			 
    
fields

    myNbShape  : Integer from Standard;
    myFAttach  : Pnt     from gp;
    mySAttach  : Pnt     from gp;
    myDirAttach: Dir     from gp;       
    myTypeDist : TypeOfDist from AIS;
    
end LengthDimension;
