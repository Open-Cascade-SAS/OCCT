-- File:	RWStepBasic_RWActionRequestAssignment.cdl
-- Created:	Fri Nov 26 16:26:30 1999 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0
-- Copyright:	Matra Datavision 1999

class RWActionRequestAssignment from RWStepBasic

    ---Purpose: Read & Write tool for ActionRequestAssignment

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    ActionRequestAssignment from StepBasic

is
    Create returns RWActionRequestAssignment from RWStepBasic;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : ActionRequestAssignment from StepBasic);
	---Purpose: Reads ActionRequestAssignment

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: ActionRequestAssignment from StepBasic);
	---Purpose: Writes ActionRequestAssignment

    Share (me; ent : ActionRequestAssignment from StepBasic;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWActionRequestAssignment;
