-- Created on: 1996-11-14
-- Created by: Philippe MANGIN
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PrefAndRec from AdvApprox inherits Cutting from AdvApprox

    ---Purpose : 
    -- inherits class Cutting; contains a list of preferential points (pi)i
    -- and a list of Recommended points used in cutting management.
    

uses Array1OfReal from TColStd

raises DomainError from Standard
    
is
    Create(RecomendedCut : Array1OfReal;
           PrefferedCut  : Array1OfReal;
           Weight        : Real = 5 ) 
    returns PrefAndRec 
    raises DomainError;  -- if  Weight <= 1
    
    Value(me; a,b : Real;
              cuttingvalue : out Real)
    returns Boolean 
    ---Purpose: 
    --     cuting value is
    --    - the recommended point nerest of (a+b)/2 
    --      if pi is in ]a,b[ or else
    --   -  the preferential point nearest of (a+b) / 2
    --     if pi is in ](r*a+b)/(r+1) , (a+r*b)/(r+1)[ where r = Weight
    --   -  or (a+b)/2 else.
    is redefined;


fields
    myRecCutting : Array1OfReal from TColStd;
    myPrefCutting: Array1OfReal from TColStd;
    myWeight     : Real;
end PrefAndRec;
