-- Created on: 2001-06-25
-- Created by: Michael KLOKOV
-- Copyright (c) 2001-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class SolidBuilder from BOP
     
    ---Purpose: 
    ---   Construct Solids from a Shell Faces  Set (SFS)
    ---
uses

    Shell            from TopoDS,
    Face             from TopoDS,
    ShapeSet         from BOP,
    LoopSet          from BOP,
    ShellFaceSet     from BOP,
    BlockBuilder     from BOP,
    BlockIterator    from BOP,
    SolidAreaBuilder from BOP

is

    Create returns SolidBuilder from BOP;
    	---Purpose:  
    	--- Empty constructor; 
    	---
    Create(theSFS: in out ShellFaceSet from BOP;
    	   theForceClassFlag: Boolean from Standard = Standard_False)
	   returns SolidBuilder from BOP;
    	---Purpose:  
    	--- The constructor that just calls the method  
    	--- InitSolidBuilder() below 
    	---
    InitSolidBuilder(me : in out;
    	    	     theSFS: in out ShellFaceSet from BOP;
		     theForceClassFlag: Boolean from Standard);
    	---Purpose: 
    	--- Launches the algorithm consisting of four steps 
    	--- 1.  Split the SFS on shells ( BOP_SFSCorrector object)      
    	--- 2.  Make Loops from shells  ( this->MakeLoops() )      
    	--- 3.  Make Areas from Loops   ( BOP_SolidAreaBuilder object)            
    	--- 4.  Make Solids from Areas  ( see methods below )   
    	---

    ---
    ---             O  u  t  p  u  t     m  e  t  h  o  d  s  
    ---
    ---  Iterator on  Solids  
    ---
    InitSolid(me: in out) 
	returns Integer from Standard;

    MoreSolid(me) 
    	returns Boolean from Standard;
    
    NextSolid(me : in out);
    ---
    ---  Iterator on  Shells  
    ---
    InitShell(me : in out) 
    	returns Integer from Standard;
    
    MoreShell(me) 
    	returns Boolean from Standard;
    
    NextShell(me : in out);

    IsOldShell(me) 
    	returns Boolean from Standard;

    OldShell(me) returns Shell from TopoDS;
    ---
    ---  Iterator on  Shells  
    ---
    InitFace(me : in out) 
    	returns Integer from Standard;

    MoreFace(me) 
    	returns Boolean from Standard;

    NextFace(me : in out);
    
    Face(me) 
    	returns Face from TopoDS; 
    	---C++: return const &
    	---Purpose:  
    	--- Returns current new face of current new shell.
    	---

    ------------------------------------------------------
    --             P  r  i  v  a  t  e    b  l  o  c  k   
    --
    MakeLoops(me: in out; theSFS: in out ShapeSet from BOP)
    	is private;

fields

    myLoopSet         : LoopSet          from BOP;
    myBlockIterator   : BlockIterator    from BOP;
    myBlockBuilder    : BlockBuilder     from BOP;
    mySolidAreaBuilder: SolidAreaBuilder from BOP;

end SolidBuilder from BOP;
