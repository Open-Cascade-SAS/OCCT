-- Created on: 1991-06-25
-- Created by: Christophe MARION
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




package BRepTest 

	---Purpose: Provides commands to test BRep.
	--          
uses
    Draw,
    TCollection
    
is
   	
    AllCommands(DI : in out Interpretor from Draw);
	---Purpose: Defines all the topology commands.

    BasicCommands(DI : in out Interpretor from Draw);
	---Purpose: Defines the basic commands.

    CurveCommands(DI : in out Interpretor from Draw);
	---Purpose: Defines the commands to build edges and wires.
	
    Fillet2DCommands(DI : in out Interpretor from Draw);
	---Purpose:  Defines the  commands  to perform add  fillets on
	--          wires and  edges.
   
    SurfaceCommands(DI : in out Interpretor from Draw);
	---Purpose: Defines the commands to build faces and shells.

    PrimitiveCommands(DI : in out Interpretor from Draw);
	---Purpose: Defines the commands to build primitives.
	
    FillingCommands(DI : in out Interpretor from Draw);
	---Purpose: Defines the commands to build primitives.
	
    SweepCommands(DI : in out Interpretor from Draw);
	---Purpose: Defines the commands to sweep shapes.
	
    TopologyCommands(DI : in out Interpretor from Draw);
	---Purpose: Defines  the    commands   to perform  topological
	--          operations. 

    FilletCommands(DI : in out Interpretor from Draw);
	---Purpose: Defines  the commands  to perform  add  fillets on
	--          shells.
   
    ChamferCommands(DI : in out Interpretor from Draw);
	---Purpose: Defines  the commands  to perform  add chamfers on
	--          shells.
	
    GPropCommands(DI : in out Interpretor from Draw);
	---Purpose: Defines commands to compute global properties.
	
    MatCommands(DI : in out Interpretor from Draw);
    	---Purpose: Defines commands to compute and to explore the map of the
    	--          Bisecting locus.


    DraftAngleCommands(DI : in out Interpretor from Draw);
	---Purpose: Defines the commands to modify draft angles of the
	--          faces of a shape.


    FeatureCommands(DI : in out Interpretor from Draw);
	---Purpose: Defines the commands to create features on a shape.


    OtherCommands(DI : in out Interpretor from Draw);
	---Purpose: Defines the auxiliary topology commands.
	

    ExtremaCommands(DI : in out Interpretor from Draw);
	---Purpose: Defines the extrema commands.
	

    CheckCommands(DI : in out Interpretor from Draw);
	---Purpose: Defines the checkshape command.

    PlacementCommands(DI : in out Interpretor from Draw);
	---Purpose: Defines the placement  command.
	--          

    ProjectionCommands(DI : in out Interpretor from Draw);
	---Purpose: Defines the commands to project a wire on a shape.
	--          
    ShellCommands(DI : in out Interpretor from Draw);
	---Purpose: Defines the commands to prepare shell commands.

end BRepTest;

