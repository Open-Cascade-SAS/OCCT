-- Created on: 1993-08-11
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




deferred class PointRepresentation from PBRep inherits Persistent

	---Purpose: Root class for points representations.

uses
    Location from PTopLoc

is
    Initialize(P : Real;
    	       L : Location from PTopLoc);
    	---Level: Internal 
	       
    Location(me) returns Location from PTopLoc
    is static;
    	---Level: Internal 
		
    Parameter(me) returns Real
    is static;
    	---Level: Internal 
		
    Parameter(me : mutable; P : Real)
    is static;
    	---Level: Internal 
		
    Next(me) returns PointRepresentation from PBRep
    is static;
    	---Level: Internal 
		
    Next(me : mutable; N :  PointRepresentation from PBRep)
    is static;
    	---Level: Internal 

    ------------------------------------------------------
    -- What kind of representation : used to speed Mapping
    ------------------------------------------------------

    IsPointOnCurve(me)          returns Boolean
	---Purpose: A point on a 3d curve.
    is virtual;
	
    IsPointOnCurveOnSurface(me) returns Boolean
	---Purpose: A point on a 2d curve on a surface.
    is virtual;

    IsPointOnSurface(me)        returns Boolean
	---Purpose: A point on a surface.
    is virtual;
    
fields
    
    myLocation  : Location from PTopLoc;
    myParameter : Real;
    myNext      : PointRepresentation from PBRep;

end PointRepresentation;
