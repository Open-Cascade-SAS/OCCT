-- Created on: 1995-12-11
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Edge from BRepCheck inherits Result from BRepCheck

	---Purpose: 

uses Shape               from TopoDS,
     Edge                from TopoDS,
     CurveRepresentation from BRep,
     HCurve              from Adaptor3d,
     Status              from BRepCheck

is

    Create(E: Edge from TopoDS)
    
    	returns Edge from BRepCheck;


    InContext(me: mutable; ContextShape: Shape from TopoDS);
    


    Minimum(me: mutable);
    

    
    Blind(me: mutable);


    GeometricControls(me)
    
    	returns Boolean from Standard
	is static;


    GeometricControls(me: mutable; B: Boolean from Standard)
    
	is static;

    Tolerance(me: mutable) returns Real from Standard 

    	is static;

    SetStatus(me: mutable;
              theStatus:Status from BRepCheck)

          --- Purpose: Sets status of Edge;
	is static;

    CheckPolygonOnTriangulation(me: mutable; theEdge: Edge from TopoDS)
	  --- Purpose: Checks, if polygon on triangulation of heEdge
     -- is out of 3D-curve of this edge.
        returns Status from BRepCheck
	is static;

fields

    myCref   : CurveRepresentation from BRep;
    myHCurve : HCurve              from Adaptor3d;
    myGctrl  : Boolean from Standard;

end Edge;
