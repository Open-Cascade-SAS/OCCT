-- Created on: 1995-12-07
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.





class ReadWriteModule from RWStepAP214  inherits ReadWriteModule from StepData

	---Purpose : General module to read and write StepAP214 entities

uses Transient,
     SequenceOfAsciiString    from TColStd,
     AsciiString              from TCollection,
     Check                    from Interface,
     StepReaderData           from StepData,
     StepWriter               from StepData

is

	Create returns mutable ReadWriteModule from RWStepAP214;

	CaseStep (me; atype : AsciiString from TCollection) returns Integer;
	---Purpose : associates a positive Case Number to each type of StepAP214 entity,
	-- given as a String defined in the EXPRESS form

	CaseStep(me; types : SequenceOfAsciiString from TColStd) returns Integer is redefined;
	---Purpose : associates a positive Case Number to each type of StepAP214 Complex entity,
	-- given as a String defined in the EXPRESS form

	IsComplex (me; CN : Integer) returns Boolean is redefined;
	---Purpose : returns True if the Case Number corresponds to a Complex Type

	StepType (me; CN : Integer) returns AsciiString from TCollection;
	---Purpose : returns a StepType (defined in EXPRESS form which belongs to a 
	-- Type of Entity, identified by its CaseNumber determined by Protocol
	---C++ : return const &

	ComplexType (me; CN : Integer;
                 types : in out SequenceOfAsciiString from TColStd)
            returns Boolean  is redefined;

	ReadStep (me; CN : Integer; data : StepReaderData; num : Integer;
	            ach : in out Check; ent : mutable Transient);

	WriteStep (me; CN : Integer; SW : in out StepWriter; ent : Transient);

end ReadWriteModule;
