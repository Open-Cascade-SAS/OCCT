-- Created on: 1994-09-14
-- Created by: Christian CAILLET
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class WorkLibrary  from StepSelect  inherits WorkLibrary  from IFSelect

    ---Purpose : Performs Read and Write a STEP File with a STEP Model
    --           Following the protocols, Copy may be implemented or not

uses CString, Transient, 
     CheckIterator, InterfaceModel, Protocol from Interface,
     Messenger from Message,
     EntityIterator, CopyTool,
     ContextWrite

is

    Create (copymode : Boolean = Standard_True)
    	 returns WorkLibrary from StepSelect;
    ---Purpose : Creates a STEP WorkLibrary
    --           <copymode> precises whether Copy is implemented or not

    SetDumpLabel (me : mutable; mode : Integer);
    ---Purpose : Selects a mode to dump entities
    --           0 (D) : prints numbers, then displays table number/label
    --           1 : prints labels, then displays table label/number
    --           2 : prints labels onky

    ReadFile (me; name : CString;
    	      model    : out InterfaceModel;
    	      protocol : Protocol from Interface)
    	  returns Integer;
    ---Purpose : Reads a STEP File and returns a STEP Model (into <mod>),
    --           or lets <mod> "Null" in case of Error
    --           Returns 0 if OK, 1 if Read Error, -1 if File not opened

    WriteFile (me; ctx : in out ContextWrite)  returns Boolean;
    ---Purpose : Writes a File from a STEP Model
    --           Returns False (and writes no file) if <ctx> does not bring a
    --           STEP Model

    CopyModel (me;
    	       original : InterfaceModel;
	       newmodel : InterfaceModel;
	       list     : EntityIterator;
	       TC       : in out CopyTool)
	returns Boolean  is redefined;
    ---Purpose : Performs the copy of entities from an original model to a new
    --           one. Works according <copymode> :
    --           if True, standard copy is run
    --           else nothing is done and returned value is False

    DumpEntity (me;
    	    	model    : InterfaceModel;
		protocol : Protocol from Interface;
		entity   : Transient;
		S        : Messenger from Message;
		level    : Integer);
    ---Purpose : Dumps an entity under STEP form, i.e. as a part of a Step file
    --           Works with a StepDumper.
    --           Level 0 just displays type; level 1 displays the entity itself
    --           and level 2 displays the entity plus its shared ones (one
    --           sub-level : immediately shared entities)

fields

    thecopymode : Boolean;
    thelabmode  : Integer;

end WorkLibrary;
