-- Created on: 2005-01-21
-- Created by: Alexander SOLOVYOV
-- Copyright (c) 2005-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SensitivePolyhedron from MeshVS inherits SensitiveEntity from Select3D

uses
    EntityOwner                from SelectBasics,
    Projector                  from Select3D,
    Location                   from TopLoc,
    Real                       from Standard,
    Boolean                    from Standard,
    Array1OfPnt2d              from TColgp,
    SequenceOfInteger          from TColStd,
    Box2d                      from Bnd,
    Lin                        from gp,
    ListOfBox2d                from SelectBasics,
    PickArgs                   from SelectBasics,
    Array1OfPnt                from TColgp,
    HArray1OfPnt               from TColgp,
    HArray1OfPnt2d             from TColgp,
    HArray1OfSequenceOfInteger from MeshVS,
    XY                         from gp

is
    Create( Owner : EntityOwner from SelectBasics;
            Nodes : Array1OfPnt from TColgp;
            Topo  : HArray1OfSequenceOfInteger from MeshVS ) returns SensitivePolyhedron from MeshVS;

    Project( me:mutable; aProjector: Projector from Select3D ) is redefined;

    GetConnected( me:mutable; aLocation: Location from TopLoc ) returns SensitiveEntity from Select3D 
       is redefined;
   
    Matches (me : mutable;
             thePickArgs : PickArgs from SelectBasics;
             theMatchDMin, theMatchDepth : out Real from Standard)
      returns Boolean is redefined;

    Matches( me                  : mutable; 
             XMin,YMin,XMax,YMax : Real from Standard;
             aTol                : Real from Standard ) returns Boolean from Standard is redefined;

    Matches( me       : mutable; 
             Polyline : Array1OfPnt2d from TColgp;
	     aBox     : Box2d from Bnd;
             aTol     : Real from Standard ) returns Boolean from Standard is redefined;

    GetBox2d( me; aBox : out Box2d from Bnd ) is protected;

    FindIntersection( me; NodesIndices : SequenceOfInteger from TColStd;
                          EyeLine      : Lin from gp ) returns Real is protected;

    ComputeDepth( me; EyeLine: Lin from gp ) returns Real from Standard is virtual;

--  ComputeSize( me ) returns Real from Standard is redefined;

    Areas( me: mutable; aResult : in out ListOfBox2d from SelectBasics ) is redefined;

fields
    myNodes   : HArray1OfPnt from TColgp;
    myNodes2d : HArray1OfPnt2d from TColgp;
    myTopo    : HArray1OfSequenceOfInteger from MeshVS;
    myCenter  : XY from gp;

end SensitiveEntity;

