-- Created on: 1993-07-13
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class Curve2d from BRepAdaptor inherits Curve from Geom2dAdaptor

	---Purpose: The Curve2d from BRepAdaptor allows to use an Edge
	--          on   a Face like   a  2d   curve. (curve  in   the
	--          parametric space).
	--          
	--          It  has  the methods    of the class Curve2d  from
	--          Adpator. 
	--          
	--          It  is created or  initialized with a  Face and an
	--          Edge.  The methods are  inherited from  Curve from
	--          Geom2dAdaptor. 

uses
    Face from TopoDS,
    Edge from TopoDS

raises
    NullObject from Standard

is

    Create returns Curve2d from BRepAdaptor;
	---Purpose: Creates an uninitialized curve2d.

    Create(E : Edge from TopoDS; F : Face from TopoDS)
    returns Curve2d from BRepAdaptor
	---Purpose: Creates with the pcurve of <E> on <F>.
    raises
    	NullObject from Standard; -- if <E> has no pcurve on <F>
	
    Initialize(me : in out; E : Edge from TopoDS; F : Face from TopoDS)
	---Purpose: Initialize with the pcurve of <E> on <F>.
    raises
    	NullObject from Standard -- if <E> has no pcurve on <F>
    is static;
    
    Edge(me) returns Edge from TopoDS
	---Purpose: Returns the Edge.
	--          
	---C++: return const &
    is static;

    Face(me) returns Face from TopoDS
	---Purpose: Returns the Face.
	--          
	---C++: return const &
    is static;

fields

    myEdge : Edge from TopoDS;
    myFace : Face from TopoDS;
	
end Curve2d;
