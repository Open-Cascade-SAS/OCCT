-- Created on: 1993-08-12
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class AncestorsTool from TopOpeBRepTool

	-- as AncestorsTool from TopOpeInter 
	--  (Shape from TopoDS,
	--   IndexedDataMapOfShapeListOfShape from TopTools)
	
	---Purpose: Describes the ancestors tool needed by 
	--          the class DSFiller from TopOpeInter.
	--          
	-- This class has been created because it is not possible
	-- to instantiate the argument TheAncestorsTool (of
	-- DSFiller from TopOpeInter) with a  package (TopExp)
	-- giving services as package methods.

uses

    Shape from TopoDS,
    ShapeEnum from TopAbs,
    IndexedDataMapOfShapeListOfShape from TopTools

is

    MakeAncestors(myclass;
    	    	  S  : Shape from TopoDS;
		  TS : ShapeEnum from TopAbs;
		  TA : ShapeEnum from TopAbs;
		  M  : in out IndexedDataMapOfShapeListOfShape from TopTools); 
		  
	---Purpose: same as package method TopExp::MapShapeListOfShapes()
		  
      		      
end AncestorsTool;
