-- Created on: 1994-04-01
-- Created by: Laurent BUCHARD
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class Intersector3d from BRepClass3d 
    
    
uses 
    Lin               from gp,
    Pnt               from gp,
    Face              from TopoDS,
    Shape             from TopoDS,
    State             from TopAbs,
    TransitionOnCurve from IntCurveSurface
    
is

    Create returns Intersector3d from BRepClass3d;
    	---Purpose: Empty constructor.
    	          
    Perform(me: in out;  L    : Lin     from gp;
    	                 Prm  : Real    from Standard;
			 Tol  : Real    from Standard;
			 F    : Face    from TopoDS) 
	---Purpose: Perform the intersection between the 
	--          segment L(0) ... L(Prm) and the Shape <Sh>.
	--          
	--          Only the point with the smallest parameter on the 
	--          line is returned. 
	--          
	--          The Tolerance <Tol> is used to determine if the 
	--          first point of the segment is near the face. In 
	--          that case, the parameter of the intersection point 
	--          on the line can be a negative value (greater than -Tol).
    is static;
    
    
    IsDone(me)  
    	---Purpose: True is returned when the intersection have been computed.
    	---C++: inline
    returns Boolean from Standard
    is static;
    
    
    HasAPoint(me) 
    	---Purpose: True is returned if a point has been found.
    	---C++: inline
    returns Boolean from Standard
    is static;
    
	 
    UParameter(me) 
    	---Purpose: Returns the U parameter of the intersection point 
    	--          on the surface.
    	---C++: inline
    returns Real from Standard
    is static;

    VParameter(me) 
    	---Purpose: Returns the V parameter of the intersection point 
    	--          on the surface.
    	---C++: inline
    returns Real from Standard
    is static;

    WParameter(me) 
    	---Purpose: Returns the parameter of the intersection point 
    	--          on the line.
    	---C++: inline
    returns Real from Standard
    is static;


    Pnt(me)
	---Purpose: Returns the geometric point of the intersection 
	--          between the line and the surface.
    	---C++: inline
	---C++: return const &
    returns Pnt from gp
    is static;
    
    
    Transition(me) 
    	---Purpose: Returns the transition of the line on the surface.
    	---C++: inline
    returns TransitionOnCurve from IntCurveSurface
    is static;
    

    State(me) 
    	---Purpose: Returns the state of the point on the face.
    	--          The values can be either TopAbs_IN 
    	--             ( the point is in the face)
    	--           or TopAbs_ON
    	--             ( the point is on a boudary of the face).
    	---C++: inline
       
    returns State from TopAbs
    is static;
    
    Face(me) 
    	---Purpose: Returns the significant face used to determine
    	--          the intersection. 
    	--          
    	---C++: inline
    	---C++: return const &
    returns Face from TopoDS
    is static;
    
    
	---------------------- Local Geometry avec courbureS dans une 
	--                     direction et la direction normale     

fields

    pnt                :  Pnt                 from gp;
    U                  :  Real                from Standard;
    V                  :  Real                from Standard;
    W                  :  Real                from Standard;
    transition         :  TransitionOnCurve   from IntCurveSurface;
    done               :  Boolean             from Standard;
    hasapoint          :  Boolean             from Standard;
    state              :  State               from TopAbs;
    face               :  Face                from TopoDS;

end Intersector3d;

   






