-- File:        CartesianPoint.cdl
-- Created:     Mon Dec  4 12:02:24 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWCartesianPoint from RWStepGeom

	---Purpose : Read & Write Module for CartesianPoint

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     CartesianPoint from StepGeom

is

	Create returns RWCartesianPoint;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable CartesianPoint from StepGeom);

	WriteStep (me; SW : in out StepWriter; ent : CartesianPoint from StepGeom);

end RWCartesianPoint;
