-- Created on: 1993-02-05
-- Created by: Gilles DEBARBOUILLE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class DynamicDerivedClass from Dynamic 


inherits

    DynamicClass from Dynamic
    
	---Purpose: The object of  this class is  to allow, as in  the
	--          C++ language,    the  possibility  to   define   a
	--          DynamicDerivedClass  which  inherits from   one or
	--          more DynamicClass.

uses

    CString from Standard,
    Method            from Dynamic,
    DynamicInstance   from Dynamic,
    SequenceOfClasses from Dynamic

is

    Create(aname : CString from Standard) returns mutable DynamicDerivedClass from Dynamic;
    
    ---Level: Public 
    
    ---Purpose: Creates a new instance of this class with <aname> as name.
    
    AddClass(me : mutable ; aclass : any DynamicClass from Dynamic)
    
    ---Level: Public 
    
    ---Purpose: Adds another class <aclass> to the sequence of derived
    --          classes.
    
    is static;
    
    Method(me ; amethod : CString from Standard) returns any Method from Dynamic
    
    ---Level: Public 
    
    ---Purpose: Starting with  the name of  a method,  this  redefined
    --          method searches for   the  right method object  in the
    --          sequence of methods  of  the derived class and  in all
    --          the inherited classes.

    is redefined;
    
    Instance(me) returns mutable DynamicInstance from Dynamic
    
    ---Level: Public 
    
    ---Purpose: Defines an instance of this class definition.

    is redefined;

fields

    thesequenceofclasses : SequenceOfClasses from Dynamic;

end DynamicDerivedClass;
