-- Created on: 2011-06-02
-- Created by: Oleg AGASHIN
-- Copyright (c) 2011-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class VertexTool from BRepMesh 

  ---Purpose: Describes the data structure necessary for the
  --          mesh algorithm and contains the vertices in UV space.

  uses    Boolean from Standard,
          Integer from Standard,
          Real from Standard,
          XY from gp,
          ListOfInteger from BRepMesh,
          VertexCellFilter from BRepMesh,
          VertexInspector from BRepMesh,
          BaseAllocator from BRepMesh,
          Vertex from BRepMesh,
          DataMapOfIntegerListOfInteger from BRepMesh,
          Array1OfReal from TColStd

  is      Create (theAlloc : in BaseAllocator from BRepMesh)
          returns VertexTool from BRepMesh;


          Create     (nbComp   : in Integer from Standard;
                      theAlloc : in BaseAllocator from BRepMesh)
             ---Purpose: Constructs a VertexTool with an  evaluation of the
             --          number of vertices.
             returns VertexTool from BRepMesh;

          SetCellSize(me                 : in out;
                      theSize            : in Real from Standard)
            ---Purpose: Sets new size for cellfilter.
            is static;
            
          SetCellSize(me                 : in out;
                       theXSize            : in Real from Standard;
                       theYSize            : in Real from Standard)
             ---Purpose: Sets new size for cellfilter.
             is static;

          SetTolerance(me                 : in out;
                      theTol            : in Real from Standard)
            ---Purpose: Sets new size for cellfilter.
            is static;
            
          SetTolerance(me                 : in out;
                       theTolX            : in Real from Standard;
                       theTolY            : in Real from Standard)
             ---Purpose: Sets new size for cellfilter.
             is static;

          Add       (me       : in out;
                     theVertex: in Vertex from BRepMesh;
                     theParams: in ListOfInteger from BRepMesh)
            ---Purpose: Adds a vertex to the tool.
            returns Integer from Standard is static;

          Add       (me       : in out;
                     theVertex: in Vertex from BRepMesh)
            ---Purpose: Adds a vertex to the tool.
            returns Integer from Standard is static;

          Delete   (me : in out; theIndex : Integer from Standard) 
            ---Purpose: Deletes a vertex from the tool.
            is static;

          FindFromIndex   (me; theIndex : Integer from Standard)
            ---Purpose: Returns data assigned to theIndex.
            ---C++: alias operator() 
            ---C++: return &
            returns ListOfInteger from BRepMesh is static;
          
          FindKey   (me: out; theIndex: Integer from Standard)
            ---Purpose: Selects the vertex by theIndex.
            ---C++: return const &
            returns Vertex from BRepMesh is static;
            
          FindIndex (me: out;
	  	     theVertex: Vertex from BRepMesh)
            ---Purpose: Returns an index of theVertex.
            returns Integer from Standard is static;
            
          Extent    (me)
            ---Purpose: Returns a number of vertices.
            returns Integer from Standard is static;
            
          IsEmpty   (me)
            ---Purpose: Returns True when the map contains no keys.
            returns Boolean from Standard is static;
          
          Substitute(me: in out; Index: Integer from Standard;
                     theVertex: Vertex from BRepMesh;
                     theData  : ListOfInteger from BRepMesh)
            ---Purpose: Substitutes vertex with Index on
            --          theVertex with attributes theData.
            is static;
            
          RemoveLast(me: out)
            ---Purpose: Remove last node from the structure.
            is static;
            
          GetListOfDelNodes(me)
            ---Purpose: Returns the list with indexes of
            --          vertices that have Movability attribute
            --          equal to BRepMesh_Deleted and can be 
            --          replaced with another node.
            ---C++: return const &
            returns ListOfInteger from BRepMesh
            is static;
            
          ExpandPoint(me: in out;
                      thePnt: in XY from gp;
                      theMinPnt: out XY from gp;
                      theMaxPnt: out XY from gp)
            is static private;
            
          Statistics(me; S: in out OStream from Standard)
            ---Purpose: Prints statistics.
            is static;
            
  fields  myAllocator    : BaseAllocator from BRepMesh;
          myCellFilter   : VertexCellFilter from BRepMesh;
          mySelector     : VertexInspector from BRepMesh;
          myLinksMap     : DataMapOfIntegerListOfInteger from BRepMesh;
          myTol          : Array1OfReal from TColStd;

end CircleTool;
