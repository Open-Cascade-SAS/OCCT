-- Created on: 1993-01-09
-- Created by: CKY / Contract Toubro-Larsen ( TCD )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class TabulatedCylinder from IGESGeom  inherits IGESEntity

        ---Purpose: defines IGESTabulatedCylinder, Type <122> Form <0>
        --          in package IGESGeom
        --          A tabulated cylinder is a surface formed by moving a line
        --          segment called generatrix parallel to itself along a curve
        --          called directrix. The curve may be a line, circular arc,
        --          conic arc, parametric spline curve, rational B-spline
        --          curve or composite curve.

uses

        Pnt         from gp,
        XYZ         from gp

is

        Create returns mutable TabulatedCylinder;

        -- Specific Methods pertaining to the class

        Init (me         : mutable;
              aDirectrix : IGESEntity;
              anEnd      : XYZ);
        ---Purpose : This method is used to set the fields of the class
        --           TabulatedCylinder
        --       - aDirectrix : Directrix Curve of the tabulated cylinder
        --       - anEnd      : Coordinates of the terminate point of the
        --                      generatrix
        -- The start point of the directrix is identical to the start
        -- point of the generatrix

        Directrix (me) returns IGESEntity;
        ---Purpose : returns the directrix curve of the tabulated cylinder

        EndPoint(me) returns Pnt;
        ---Purpose : returns end point of generatrix of the tabulated cylinder

        TransformedEndPoint(me) returns Pnt;
        ---Purpose : returns end point of generatrix of the tabulated cylinder
        -- after applying Transf. Matrix

fields

--
-- Class    : IGESGeom_TabulatedCylinder
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class TabulatedCylinder.
--
-- Reminder : A TabulatedCylinder instance is defined by :
--            A directrix curve and the coordinates of end points of
--            directrix curve

        theDirectrix : IGESEntity;
        theEnd       : XYZ;

end TabulatedCylinder;
