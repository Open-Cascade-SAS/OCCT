-- Created on: 1998-08-17
-- Created by: Philippe MANGIN
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ShapeLaw from BRepFill inherits  SectionLaw  from  BRepFill

	---Purpose: Build Section Law, with an Vertex, or an Wire
        ---Level: Advanced
       
uses 
 SectionLaw          from GeomFill,  
 HArray1OfSectionLaw from  GeomFill, 
 HArray1OfShape      from  TopTools,  
 Shape               from  GeomAbs,
 Vertex              from  TopoDS, 
 Wire                from  TopoDS,  
 Edge                from  TopoDS,  
 Shape               from  TopoDS, 
 Function            from  Law

is  
  Create (V:  Vertex  from  TopoDS;   
          Build  :  Boolean = Standard_True )  
    ---Purpose: Construct an constant Law  
  returns  ShapeLaw  from BRepFill;   

  Create (W:Wire  from  TopoDS;   
          Build :  Boolean = Standard_True)   
     ---Purpose: Construct an constant Law   
  returns ShapeLaw from BRepFill;  
   
  Create  (W:  Wire  from  TopoDS;  
           L:  Function  from  Law; 
           Build :  Boolean = Standard_True)   
    ---Purpose: Construct an evolutive Law         
  returns ShapeLaw from BRepFill;      

  IsVertex(me) 
    ---Purpose: Say if the input shape is a  vertex. 
  returns  Boolean   
  is  redefined; 
   
  IsConstant(me) 
    ---Purpose: Say if the Law is  Constant.        
  returns  Boolean   
  is  redefined;        

  ConcatenedLaw(me)  
   ---Purpose: Give the law build on a concaneted section         
  returns SectionLaw from GeomFill 
  is  redefined;    
  
  Continuity(me; Index  :  Integer; 
    	         TolAngular  :  Real)
  returns  Shape  from  GeomAbs  
  is  redefined;  
   
  VertexTol(me; Index  :  Integer;   
                Param  :  Real) 
  returns  Real   
  is  redefined;  
  
  Vertex(me;  Index  :  Integer; 
              Param  :  Real) 
  returns Vertex  from  TopoDS 
  is  redefined;	    
   
  D0(me:mutable;  Param  :  Real;   
     S  :  out  Shape  from  TopoDS)   
    is  redefined;  
   
  Edge(me; Index  :  Integer)  
   ---C++: return const &
   ---C++: inline
  returns  Edge  from  TopoDS;  
   
  Init(me  :  mutable;  B  :  Boolean)  is  private;
   
fields
  myShape:  Shape          from  TopoDS;
  myEdges:  HArray1OfShape from  TopTools;   
  TheLaw :  Function       from  Law;   
  vertex :  Boolean        from  Standard is  protected; 
end ShapeLaw;
