-- Created on: 1993-09-30
-- Created by: Denis PASCAL
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SC from GraphTools inherits TShared from MMgt

    ---Purpose: This  class is used  to  identify a  Strong Component.
    --          The user has not to used its methods.

uses SCList            from GraphTools,
     SequenceOfInteger from TColStd

raises OutOfRange   from Standard,
       NoSuchObject from Standard
    
is

    Create returns mutable SC;
	
    Reset (me : mutable);
    ---Level: Public

    AddVertex (me : mutable; V : Integer from Standard); 
    ---Level: Public

    NbVertices (me) returns Integer from Standard;
    ---Level: Public

    GetVertex (me; index: Integer from Standard) 
    ---Level: Public
    returns Integer from Standard;
	
    AddFrontSC (me : mutable; SC : SC from GraphTools);
    ---Level: Public
 
    GetFrontSC (me) returns SCList from GraphTools;
    ---Level: Public
    ---C++: return const & 	
	
    AddBackSC (me : mutable; SC : SC from GraphTools);
    ---Level: Public

    GetBackSC (me) returns SCList from GraphTools;
    ---Level: Public
    ---C++: return const & 	

fields
	
    myBackSC   : SCList            from GraphTools;
    myVertices : SequenceOfInteger from TColStd;
    myFrontSC  : SCList            from GraphTools;

end SC;


