-- Created on: 1995-12-07
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




deferred class Result from BRepCheck inherits TShared from MMgt

	---Purpose: 

uses Shape                                       from TopoDS,
     ListOfStatus                                from BRepCheck,
     DataMapOfShapeListOfStatus                  from BRepCheck,
     DataMapIteratorOfDataMapOfShapeListOfStatus from BRepCheck

raises NoSuchObject from Standard

is

    Initialize;

    Init(me: mutable; S: Shape from TopoDS);


    InContext(me: mutable; ContextShape: Shape from TopoDS)
    
    	is deferred;


    Minimum(me: mutable)
    
    	is deferred;

    
    Blind(me: mutable)
    
    	is deferred;

    SetFailStatus(me: mutable; S: Shape from TopoDS);


    Status(me)
    
    	returns ListOfStatus from BRepCheck
	---C++: return const&
	---C++: inline
	is static;

    IsMinimum(me)
    
    	returns Boolean from Standard
	---C++: inline
	is static;


    IsBlind(me)
    
    	returns Boolean from Standard
	---C++: inline
	is static;


    StatusOnShape(me: mutable; S: Shape from TopoDS)
	---Purpose: If  not  already   done,  performs the   InContext
	--          control and returns the list of status.
    	returns ListOfStatus from BRepCheck
	---C++: return const&
	raises
	    NoSuchObject from Standard
	is static;


    InitContextIterator(me: mutable)
    
    	is static;


    MoreShapeInContext(me)
    
    	returns Boolean from Standard
	---C++: inline
	is static;


    ContextualShape(me)
    
    	returns Shape from TopoDS
	---C++: return const&
	---C++: inline
	raises
	    NoSuchObject from Standard
	is static;


    StatusOnShape(me)
    
    	returns ListOfStatus from BRepCheck
	---C++: return const&
	---C++: inline
	raises
	    NoSuchObject from Standard
	is static;


    NextShapeInContext(me: mutable)
    
    	is static;


fields

    myShape : Shape                      from TopoDS    is protected;
    myMin   : Boolean                    from Standard  is protected;
    myBlind : Boolean                    from Standard  is protected;
    myMap   : DataMapOfShapeListOfStatus from BRepCheck is protected;
    myIter  : DataMapIteratorOfDataMapOfShapeListOfStatus from BRepCheck;

end Result;
