-- Created on: 1991-09-18
-- Created by: Arnaud BOUZY
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class UnknownIterator from Expr 

	---Purpose: Describes an iterator on NamedUnknowns contained 
	--          in any GeneralExpression.
        ---Level : Internal

uses GeneralExpression from Expr,
    NamedUnknown from Expr,
    MapOfNamedUnknown from Expr

raises NoMoreObject from Standard,
    NoSuchObject from Standard

is

    Create(exp : GeneralExpression)
    returns UnknownIterator;
    
    Perform(me: in out; exp : GeneralExpression)
    is static private;
    
    More(me)
    returns Boolean
    is static;
    
    Next(me : in out)
    raises NoMoreObject
    is static;
    
    Value(me)
    returns NamedUnknown
    raises NoSuchObject
    is static;

fields

    myMap : MapOfNamedUnknown;
    myCurrent : Integer;

end UnknownIterator;
