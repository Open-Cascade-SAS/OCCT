-- Created on: 1997-02-06
-- Created by: Kernel
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class TypeData from Storage 

inherits TShared from MMgt

uses HSequenceOfAsciiString from TColStd,
     PType from Storage,
     AsciiString from TCollection,
     Error from Storage
     
raises NoSuchObject from Standard
is
    Create returns mutable TypeData from Storage;
    
    NumberOfTypes(me) returns Integer from Standard;
    
    IsType(me; aName : AsciiString from TCollection) returns Boolean from Standard;
    
    Types(me) returns HSequenceOfAsciiString from TColStd;

    ErrorStatus(me) returns Error from Storage;
    ErrorStatusExtension(me) returns AsciiString from TCollection;
   
    ClearErrorStatus(me : mutable);

    Clear(me : mutable); 
	
    -- PRIVATE

    AddType(me : mutable; aName : AsciiString from TCollection; aTypeNum : Integer from Standard) is private;
    ---Purpose: add a type to the list
    
    Type(me; aTypeNum : Integer from Standard) returns AsciiString from TCollection
      raises NoSuchObject is private;
    ---Purpose: returns the name of the type with number <aTypeNum>
    
    Type(me; aTypeName : AsciiString from TCollection) returns Integer from Standard
      raises NoSuchObject is private;
    ---Purpose: returns the name of the type with number <aTypeNum>

    SetErrorStatus(me : mutable; anError : Error from Storage) is private;
    SetErrorStatusExtension(me : mutable; anErrorExt : AsciiString from TCollection) is private;    
    
    fields
    
      myPt                 : PType from Storage;      
      myErrorStatus        : Error from Storage;
      myErrorStatusExt     : AsciiString      from TCollection;
     
    friends class Schema from Storage
    
end;
