-- Created by: Peter KURNEV
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

class IndexRange from BOPDS 

	---Purpose: 
    	-- The class BOPDS_IndexRange is to store  
    	-- the information about range of two indices 
--uses
--raises

is 
    Create 
    	returns IndexRange from BOPDS; 
    ---C++: alias "Standard_EXPORT virtual ~BOPDS_IndexRange();"   
    ---C++: inline 
    	---Purpose:  
    	--- Empty contructor  
    	--- 
	 
    SetFirst(me:out; 
    	    theI1:Integer from Standard); 
    ---C++: inline		 
     	---Purpose: 
    	--- Modifier   
	--- Sets the first index <theI1>  of the range  
	
    SetLast(me:out; 
    	    theI2:Integer from Standard);	 
    ---C++: inline 
    	---Purpose: 
    	--- Modifier   
	--- Sets the second index <theI2>  of the range   
     
    First(me) 
    	returns Integer from Standard; 
    ---C++: inline
	---Purpose: 
    	--- Selector   
	--- Returns the first index of the range  
	
    Last(me) 
    	returns Integer from Standard; 				     
    ---C++: inline
     	---Purpose: 
    	--- Selector   
	--- Returns the second index of the range  
	 
    SetIndices(me:out; 
    	    theI1:Integer from Standard;
    	    theI2:Integer from Standard); 
    ---C++: inline	  
    	---Purpose:  
    	--- Modifier   
	--- Sets the first index of the range  <theI1>
	--- Sets the second index of the range <theI2> 
	     
    Indices(me; 
    	    theI1:out Integer from Standard;
    	    theI2:out Integer from Standard);  
    ---C++: inline     
     	---Purpose:  
    	--- Selector   
	--- Returns the first index of the range  <theI1>
	--- Returns the second index of the range <theI2>  
	
    Contains(me; 
    	    theIndex:Integer from Standard) 
    	returns Boolean from Standard;  
    ---C++: inline	 
     	---Purpose:   
    	--- Query   
	--- Returns true if the range contains <theIndex>
	
    Dump(me);
    
     
    
fields 
    myFirst  :  Integer from Standard is protected;  
    myLast   :  Integer from Standard is protected;  

end IndexRange;
