-- File:	RWStepFEA_RWNode.cdl
-- Created:	Thu Dec 12 17:51:06 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWNode from RWStepFEA

    ---Purpose: Read & Write tool for Node

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    Node from StepFEA

is
    Create returns RWNode from RWStepFEA;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : Node from StepFEA);
	---Purpose: Reads Node

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: Node from StepFEA);
	---Purpose: Writes Node

    Share (me; ent : Node from StepFEA;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWNode;
