--Copyright:      Matra Datavision 1992,1993

-- File:          OSD_Chronometer.cdl
-- Created:       Tue 18 1992
-- Author:        Stephan GARNAUD (ARM)
--                <sga@sparc4>
-- Updated:       J.P. TIRAULT August 1993
--                All methods are static methods.
--                the "Show" method returns the consumed CPU time in a Real
--                variable.
--                J.P. TIRAULT October 15 1994
--                We measure both user and system cpu time.
--                
class Chronometer from OSD

 ---Purpose: This class measures CPU time (both user and system) consumed
 --          by current process or thread. The chronometer can be started
 --          and stopped multiple times, and measures cumulative time.
 --
 --          If only the thread is measured, calls to Stop() and Show()
 --          must occur from the same thread where Start() was called 
 --          (unless chronometer is stopped); otherwise measurement will 
 --          yield false values.

is

  Create (ThisThreadOnly: Boolean = Standard_False) returns Chronometer from OSD;
  ---Purpose: Initializes a stopped Chronometer.
  --
  --          If ThisThreadOnly is True, measured CPU time will account
  --          time of the current thread only; otherwise CPU of the 
  --          process (all threads, and completed children) is measured.
  --
  ---Level: Public

  Destroy ( me : out ) is virtual;
  ---C++: alias ~

  Reset (me : in out) is virtual;
  ---Purpose: Stops and Reinitializes the Chronometer.
  ---Level: Public

  Stop (me : in out) is virtual;
  ---Purpose: Stops the Chronometer. 
  ---Level: Public

  Start (me : in out) is virtual;
  ---Purpose: Starts (after Create or Reset) or restarts (after Stop)
  --          the chronometer.
  ---Level: Public

  Show (me : in out) is virtual;
  ---Purpose: Shows the current CPU user and system time on the 
  --          standard output stream <cout>.
  --          The chronometer can be running (laps Time) or stopped.
  ---Level: Public

  Show (me : in out; os : in out OStream from Standard) is virtual;
  ---Purpose: Shows the current CPU user and system time on the output 
  --          stream <os>.
  --          The chronometer can be running (laps Time) or stopped.
  ---Level: Public

  Show (me : in out; UserSeconds : in out Real from Standard) ;
  ---Purpose: Returns the current CPU user time in a variable.
  --          The chronometer can be running (laps Time) or stopped.
  ---Level: Public

  Show (me : in out; UserSeconds : in out Real from Standard;
                     SystemSeconds : in out Real from Standard) ;
  ---Purpose: Returns the current CPU user and system time in variables.
  --          The chronometer can be running (laps Time) or stopped.
  ---Level: Public

  GetProcessCPU (myclass; UserSeconds : out Real from Standard;
                          SystemSeconds : out Real from Standard);
  ---Purpose: Returns CPU time (user and system) consumed by the current
  --          process since its start, in seconds. The actual precision of 
  --          the measurement depends on granularity provided by the system,
  --          and is platform-specific.
  ---Level: Public
  
  GetThreadCPU (myclass; UserSeconds : out Real from Standard;
                         SystemSeconds : out Real from Standard);
  ---Purpose: Returns CPU time (user and system) consumed by the current
  --          thread since its start. Note that this measurement is
  --          platform-specific, as threads are implemented and managed 
  --          differently on different platforms and CPUs.
  ---Level: Advanced
  
fields

  Stopped    : Boolean is protected;
  ThreadOnly : Boolean;
  Start_user : Real;
  Start_sys  : Real;
  Cumul_user : Real;
  Cumul_sys  : Real;

end;


