-- Created on: 2002-12-12
-- Created by: data exchange team
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class Curve3dElementProperty from StepFEA
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity Curve3dElementProperty

uses
    HAsciiString from TCollection,
    HArray1OfCurveElementInterval from StepFEA,
    HArray1OfCurveElementEndOffset from StepFEA,
    HArray1OfCurveElementEndRelease from StepFEA

is
    Create returns Curve3dElementProperty from StepFEA;
	---Purpose: Empty constructor

    Init (me: mutable; aPropertyId: HAsciiString from TCollection;
                       aDescription: HAsciiString from TCollection;
                       aIntervalDefinitions: HArray1OfCurveElementInterval from StepFEA;
                       aEndOffsets: HArray1OfCurveElementEndOffset from StepFEA;
                       aEndReleases: HArray1OfCurveElementEndRelease from StepFEA);
	---Purpose: Initialize all fields (own and inherited)

    PropertyId (me) returns HAsciiString from TCollection;
	---Purpose: Returns field PropertyId
    SetPropertyId (me: mutable; PropertyId: HAsciiString from TCollection);
	---Purpose: Set field PropertyId

    Description (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Description
    SetDescription (me: mutable; Description: HAsciiString from TCollection);
	---Purpose: Set field Description

    IntervalDefinitions (me) returns HArray1OfCurveElementInterval from StepFEA;
	---Purpose: Returns field IntervalDefinitions
    SetIntervalDefinitions (me: mutable; IntervalDefinitions: HArray1OfCurveElementInterval from StepFEA);
	---Purpose: Set field IntervalDefinitions

    EndOffsets (me) returns HArray1OfCurveElementEndOffset from StepFEA;
	---Purpose: Returns field EndOffsets
    SetEndOffsets (me: mutable; EndOffsets: HArray1OfCurveElementEndOffset from StepFEA);
	---Purpose: Set field EndOffsets

    EndReleases (me) returns HArray1OfCurveElementEndRelease from StepFEA;
	---Purpose: Returns field EndReleases
    SetEndReleases (me: mutable; EndReleases: HArray1OfCurveElementEndRelease from StepFEA);
	---Purpose: Set field EndReleases

fields
    thePropertyId: HAsciiString from TCollection;
    theDescription: HAsciiString from TCollection;
    theIntervalDefinitions: HArray1OfCurveElementInterval from StepFEA;
    theEndOffsets: HArray1OfCurveElementEndOffset from StepFEA;
    theEndReleases: HArray1OfCurveElementEndRelease from StepFEA;

end Curve3dElementProperty;
