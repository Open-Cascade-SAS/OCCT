-- Created on: 1994-08-31
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class VertexInfo from Draft

	---Purpose: 

uses Pnt                       from gp,
     Edge                      from TopoDS,
     ListOfShape               from TopTools,
     ListOfReal                from TColStd,
     ListIteratorOfListOfShape from TopTools

raises DomainError  from Standard,
       NoMoreObject from Standard

is

    Create
    
    	returns VertexInfo from Draft;
	
	
    Add(me: in out; E: Edge from TopoDS)
    
    	is static;


    Geometry(me)
    
    	returns Pnt from gp
	is static;
	---C++: return const&


    Parameter(me: in out; E: Edge from TopoDS)
    
    	returns Real from Standard
	raises DomainError from Standard
	is static;


    InitEdgeIterator(me: in out)

    	is static;

    
    Edge(me)
    	returns Edge from TopoDS
	is static;
	---C++: return const&


    NextEdge(me: in out)
    
    	raises NoMoreObject from Standard
    	is static;


    MoreEdge(me)
    
    	returns Boolean from Standard
	is static;



    ChangeGeometry(me: in out)
    
    	returns Pnt from gp
	is static;
	---C++: return &


    ChangeParameter(me: in out; E: Edge from TopoDS)
    
    	returns Real from Standard
	is static;
	---C++: return &


fields

    myGeom    : Pnt  from gp;
    myEdges   : ListOfShape from TopTools;
    myParams  : ListOfReal  from TColStd;
    myItEd    : ListIteratorOfListOfShape from TopTools;

end VertexInfo;
