-- Created on: 1997-04-01
-- Created by: Christian CAILLET
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class MarkerMember  from StepVisual    inherits SelectInt  from StepData

    ---Purpose : Defines MarkerType as unique member of MarkerSelect
    --           Works with an EnumTool

uses CString, MarkerType from StepVisual

is

    Create returns mutable MarkerMember;

    HasName (me) returns Boolean  is redefined;
    -- returns True

    Name    (me) returns CString  is redefined;
    -- returns MARKER_TYPE

    SetName (me : mutable; name : CString)  returns Boolean  is redefined;
    -- does nothing and returns True

    EnumText (me) returns CString  is redefined;
    -- returns the string counterpart of a value

    SetEnumText (me : mutable; val : Integer; text : CString)  is redefined;
    -- considers text and interprets it to set val

    SetValue  (me : mutable; val : MarkerType from StepVisual);
    -- Sets directly the good value as enum

    Value     (me) returns MarkerType from StepVisual;

end MarkerMember;
