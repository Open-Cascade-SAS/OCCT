-- File:	IGESDefs_ToolAttributeDef.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolAttributeDef  from IGESDefs

    ---Purpose : Tool to work on a AttributeDef. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses AttributeDef from IGESDefs,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolAttributeDef;
    ---Purpose : Returns a ToolAttributeDef, ready to work


    ReadOwnParams (me; ent : mutable AttributeDef;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : AttributeDef;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : AttributeDef;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a AttributeDef <ent>, from
    --           its specific (own) parameters

    DirChecker (me; ent : AttributeDef) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : AttributeDef;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : AttributeDef; entto : mutable AttributeDef;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : AttributeDef;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolAttributeDef;
