-- Created on: 1993-08-16
-- Created by: Bruno DUMORTIER
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Chronometer from Draw inherits Drawable3D from Draw

	---Purpose: Class to store chronometer variables.

uses

    Timer from OSD,
    Display from Draw,
    Interpretor from Draw

is

    Create returns Chronometer from Draw;
    
    
    Timer(me : mutable) returns Timer from OSD
	---C++: return &
    is static;

    DrawOn(me; dis : in out Display);
	---Purpose: Does nothhing,
    
    Copy(me) returns Drawable3D from Draw
	---Purpose: For variable copy.
    is redefined;
	
    Dump(me; S : in out OStream)
	---Purpose: For variable dump.
    is redefined;

    Whatis(me;  I : in out Interpretor from Draw)
	---Purpose: For variable whatis command.
    is redefined;

fields

    myTimer : Timer from OSD;

end Chronometer;
