-- Created on: 1993-08-12
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class AncestorsTool from TopOpeBRepTool

	-- as AncestorsTool from TopOpeInter 
	--  (Shape from TopoDS,
	--   IndexedDataMapOfShapeListOfShape from TopTools)
	
	---Purpose: Describes the ancestors tool needed by 
	--          the class DSFiller from TopOpeInter.
	--          
	-- This class has been created because it is not possible
	-- to instantiate the argument TheAncestorsTool (of
	-- DSFiller from TopOpeInter) with a  package (TopExp)
	-- giving services as package methods.

uses

    Shape from TopoDS,
    ShapeEnum from TopAbs,
    IndexedDataMapOfShapeListOfShape from TopTools

is

    MakeAncestors(myclass;
    	    	  S  : Shape from TopoDS;
		  TS : ShapeEnum from TopAbs;
		  TA : ShapeEnum from TopAbs;
		  M  : in out IndexedDataMapOfShapeListOfShape from TopTools); 
		  
	---Purpose: same as package method TopExp::MapShapeListOfShapes()
		  
      		      
end AncestorsTool;
