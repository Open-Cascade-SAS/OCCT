-- Created on: 1994-01-24
-- Created by: Gilles DEBARBOUILLE
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class BooleanParameter from Dynamic

inherits
    Parameter from Dynamic     
    
	---Purpose: This class describes a parameter with a boolean 
	--          as value.

uses

   CString from Standard,
   OStream from Standard

is

    Create(aparameter : CString from Standard)
    
    ---Level: Advanced 
    
    ---Purpose: Creates a boolean parameter with <aparameter> as name.

    returns mutable BooleanParameter from Dynamic;
    
    Create(aparameter : CString from Standard; 
           avalue : Boolean from Standard) 

    ---Level: Advanced 
    
    ---Purpose: Creates a boolean parameter with <aparameter> and <avalue>
    --          respectively as name and value.

    returns mutable BooleanParameter from Dynamic;
    
    Create(aparameter , avalue : CString from Standard)
    
    ---Level: Advanced 
    
    ---Purpose: Creates a boolean parameter with <aparameter> as name 
    --          and <avalue> as value. <avalue> is a CString with two possible
    --          values which are : "Standard_True" and "Standard_False".

    returns mutable BooleanParameter from Dynamic;
    
    Value(me) returns Boolean from Standard
    
    ---Level: Public 
    
    ---Purpose: Returns the boolean value <thevalue>.
    
    is static;
    
    Value (me : mutable ; avalue : Boolean from Standard)
    
    ---Level: Advanced 
    
    --- Purpose: Sets the field <thevalue> with the boolean value <avalue>

    is static;
    
    Dump(me ; astream : in out OStream from Standard)
    
    ---Level: Internal 
    
    ---Purpose: Useful for debugging.
    
    is redefined;
    
fields

    thevalue : Boolean from Standard;

end BooleanParameter;
