-- Created on: 2008-01-20
-- Created by: Alexander A. BORODIN
-- Copyright (c) 2008-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


-- Updated:       


class SystemFont from OSD inherits TShared from MMgt

 ---Purpose: Structure for store of Font System Information

uses FontAspect,
     HAsciiString from TCollection
     

is
 Create returns SystemFont;
    ---Purpose: Creates empty font object
    ---Level: Public

 Create (
         FontName : HAsciiString;
         Aspect   : FontAspect;
         FilePath : HAsciiString )  returns SystemFont;
    ---Purpose: Creates Font object initialized with <FontName> as name
    ---         <FontAspect>.... TODO
    ---Level: Public

 Create (
         XLFD     : HAsciiString;
         FilePath : HAsciiString ) returns SystemFont;
    ---Purpose: TODO
    ---Level: Public
 
 FontName (me)
        returns HAsciiString;
    --- Purpose: Returns font family name
    ---Level: Public    
        
 FontPath (me)
        returns HAsciiString;
    --- Purpose: Returns font file path
    --- Level: Public

 FontAspect (me)
        returns FontAspect from OSD;
    --- Purpose: Returns font aspect
    --- Level: Public
    
 FontHeight (me)
        returns Integer from Standard;
    --- Purpose: Returns font height
    --- If returned value is equal -1 it means that font is resizable
    --- Level: Public

 IsValid( me )
        returns Boolean;

 fields
  MyFontName:           HAsciiString;  --Font family name
  MyFontAspect:         FontAspect;    
  MyFaceSize:           Integer;       --height of font
  MyFilePath:           HAsciiString;  --absolute path to font file
  MyVerification:       Boolean;       --indicator of font initialization errors. False if initialization is failed.

end SystemFont;
