-- Created on: 1994-09-05
-- Created by: Gilles DEBARBOUILLE
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class AbstractVariableInstance from Dynamic

	---Purpose: This class is the header class to define instances
	--          of variables.  There  are two kinds  of instances,
	--          These  are VariableInstance  which  addresses only
	--          one Variable and CompositVariableInstance which is
	--          able to address  more than one variable. This last
	--          class is useful for methods with a variable number
	--          of arguments.

inherits

    Variable from Dynamic
   

is

    Initialize;
    
    Variable(me : mutable ; avariable : Variable from Dynamic)
    
    ---Level: Public
    
    ---Purpose: This  deferred method must     be implemented in   the
    --          derived    classes for  setting    reference(s) to the
    --          corresponding variable(s)  which define the  signature
    --          of the method definition.
    
    is deferred;
 
    
end AbstractVariableInstance;
