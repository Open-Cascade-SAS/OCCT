-- Created on: 1997-12-24
-- Created by: Xuan PHAM PHU
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Edge3dInterferenceTool from TopOpeBRepDS

---Purpose: a tool computing edge / face complex transition,
--          Interferences of edge reference are given by
--          I = (T on face, G = point or vertex, S = edge)

uses
    Pnt2d from gp,
    Pnt from gp,
    Dir from gp,
    Shape from TopoDS, 
    SurfaceTransition from TopTrans,
    Interference from TopOpeBRepDS
is
	  
    Create returns Edge3dInterferenceTool from TopOpeBRepDS;

    InitPointVertex(me : in out; 
            	    IsVertex : Integer;
    	    	    VonOO    : Shape from TopoDS);
	
    Init(me : in out; 
         Eref : Shape from TopoDS; 
	 E : Shape from TopoDS;   
	 F : Shape from TopoDS;
         I : Interference from TopOpeBRepDS);
    
    Add(me : in out; 
        Eref : Shape from TopoDS; 
	E : Shape from TopoDS;   
	F : Shape from TopoDS;
        I : Interference from TopOpeBRepDS);

    Transition(me; I : mutable Interference from TopOpeBRepDS)
    is static;

fields
    
    myFaceOriented : Integer;
    myTool         : SurfaceTransition from TopTrans;
    myTole         : Real; 
    myrefdef       : Boolean;

    myIsVertex     : Integer; -- 0 : geometry is a point
                              -- 1 : geometry is a vertex of reference
                              -- 2 : geometry is a vertex of the other shape
                              -- 3 : geometry is a vertex on the 2 shapes
    myVonOO        : Shape; -- only if myisvertex = 2,3
    myP3d          : Pnt from gp;
    myTgtref       : Dir from gp;

end Edge3dInterferenceTool from TopOpeBRepDS;
