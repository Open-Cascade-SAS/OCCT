-- Created on: 1996-01-26
-- Created by: Christian CAILLET
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ContextWrite    from IFSelect

    ---Purpose : This class gathers various informations used by File Modifiers
    --           apart from the writer object, which is specific of the norm
    --           and of the physical format
    --           
    --           These informations are controlled by an object AppliedModifiers
    --           (if it is not defined, no modification is allowed on writing)
    --           
    --           Furthermore, in return, ContextModif can record Checks, either
    --           one for all, or one for each Entity. It supports trace too.

uses Transient, CString, AsciiString from TCollection,
     InterfaceModel, EntityIterator, Graph, HGraph,
     Protocol from Interface, Check, CheckIterator, GeneralModifier,
     AppliedModifiers

raises NoSuchObject

is

    Create (model : InterfaceModel; proto : Protocol;
    	    applieds : mutable AppliedModifiers;  filename : CString)
    	returns ContextWrite;
    ---Purpose : Prepares a ContextWrite with these informations :
    --           - the model which is to be written
    --           - the protocol to be used
    --           - the filename
    --           - an object AppliedModifiers to work. It gives a list of
    --             FileModifiers to be ran, and for each one it can give
    --             a restricted list of entities (in the model), else all
    --             the model is considered

    Create (hgraph : HGraph; proto : Protocol;
    	    applieds : mutable AppliedModifiers;  filename : CString)
    	returns ContextWrite;
    ---Purpose : Same as above but with an already computed Graph

    Model (me) returns InterfaceModel;
    ---Purpose : Returns the Model

    Protocol (me) returns Protocol;
    ---Purpose : Returns the Protocol;

    FileName (me) returns CString;
    ---Purpose : Returns the File Name

    AppliedModifiers (me) returns mutable AppliedModifiers;
    ---Purpose : Returns the object AppliedModifiers

    Graph (me : in out) returns Graph;
    ---Purpose : Returns the Graph, either given when created, else created
    --           the first time it is queried
    ---C++ : return const &


    	--  --    Control when running    --  --

    NbModifiers (me) returns Integer;
    ---Purpose : Returns the count of recorded File Modifiers

    SetModifier (me : in out; numod : Integer) returns Boolean;
    ---Purpose : Sets active the File Modifier n0 <numod>
    --           Then, it prepares the list of entities to consider, if any
    --           Returns False if <numod> out of range

    FileModifier (me) returns mutable GeneralModifier;
    ---Purpose : Returns the currently active File Modifier. Cast to be done
    --           Null if not properly set : must be test IsNull after casting

    IsForNone (me) returns Boolean;
    ---Purpose : Returns True if no modifier is currently set

    IsForAll  (me) returns Boolean;
    ---Purpose : Returns True if the current modifier is to be applied to
    --           the whole model. Else, a restricted list of selected entities
    --           is defined, it can be exploited by the File Modifier

    NbEntities (me) returns Integer;
    ---Purpose : Returns the total count of selected entities

    Start (me : in out);
    ---Purpose : Starts an iteration on selected items. It takes into account
    --           IsForAll/IsForNone, by really iterating on all selected items.

    More (me) returns Boolean;
    ---Purpose : Returns True until the iteration has finished

    Next (me : in out);
    ---Purpose : Advances the iteration

    Value (me) returns  Transient  raises NoSuchObject;
    ---Purpose : Returns the current selected entity in the model


    	-- --    Trace and Check    -- --

    AddCheck (me : in out; check : Check)  is static;
    ---Purpose : Adds a Check to the CheckList. If it is empty, nothing is done
    --           If it concerns an Entity from the Model (by SetEntity)
    --           to which another Check is attached, it is merged to it.
    --           Else, it is added or merged as to GlobalCheck.

    AddWarning (me : in out; start : Transient; mess : CString; orig : CString = "");
    ---Purpose : Adds a Warning Message for an Entity from the Model
    --           If <start> is not an Entity from the model (e.g. the
    --           model itself) this message is added to Global Check.

    AddFail    (me : in out; start : Transient; mess : CString; orig : CString = "");
    ---Purpose : Adds a Fail Message for an Entity from the Model
    --           If <start> is not an Entity from the model (e.g. the
    --           model itself) this message is added to Global Check.

    CCheck (me : in out; num : Integer = 0) returns Check;
    ---Purpose : Returns a Check given an Entity number (in the Model)
    --           by default a Global Check. Creates it the first time.
    --           It can then be acknowledged on the spot, in condition that the
    --           caller works by reference ("Interface_Check& check = ...")

    CCheck (me : in out; start : Transient) returns Check;
    ---Purpose : Returns a Check attached to an Entity from the Model
    --           It can then be acknowledged on the spot, in condition that the
    --           caller works by reference ("Interface_Check& check = ...")

    CheckList (me) returns CheckIterator  is static;
    ---Purpose : Returns the complete CheckList

fields

    themodel : InterfaceModel;
    theproto : Protocol;
    thefile  : AsciiString;
    theapply : AppliedModifiers;
    thehgraf : HGraph;
    thecheck : CheckIterator;
    thenumod : Integer;
    thenbent : Integer;
    thecurr  : Integer;
    themodif : GeneralModifier;

end ContextWrite;
