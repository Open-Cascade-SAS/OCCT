-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class TextLiteral from StepVisual 

inherits GeometricRepresentationItem from StepGeom

uses

	HAsciiString from TCollection, 
	Axis2Placement from StepGeom, 
	TextPath from StepVisual, 
	FontSelect from StepVisual
is

	Create returns mutable TextLiteral;
	---Purpose: Returns a TextLiteral


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aLiteral : mutable HAsciiString from TCollection;
	      aPlacement : Axis2Placement from StepGeom;
	      aAlignment : mutable HAsciiString from TCollection;
	      aPath : TextPath from StepVisual;
	      aFont : FontSelect from StepVisual) is virtual;

	-- Specific Methods for Field Data Access --

	SetLiteral(me : mutable; aLiteral : mutable HAsciiString);
	Literal (me) returns mutable HAsciiString;
	SetPlacement(me : mutable; aPlacement : Axis2Placement);
	Placement (me) returns Axis2Placement;
	SetAlignment(me : mutable; aAlignment : mutable HAsciiString);
	Alignment (me) returns mutable HAsciiString;
	SetPath(me : mutable; aPath : TextPath);
	Path (me) returns TextPath;
	SetFont(me : mutable; aFont : FontSelect);
	Font (me) returns FontSelect;

fields

	literal : HAsciiString from TCollection;
	placement : Axis2Placement from StepGeom; -- a SelectType
	alignment : HAsciiString from TCollection;
	path : TextPath from StepVisual; -- an Enumeration
	font : FontSelect from StepVisual; -- a SelectType

end TextLiteral;
