-- Created on: 1995-04-20
-- Created by: Tony GEORGIADES
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

--		Modified Tue Sep 19 1995 by Jean-Louis Frenkel
--		Modified Tue Jan 19 1999 by Louis Dusuzeau

package Resource
    ---Purpose: Resources management.
    --          A RESOURCE is a parameter saved on a file and used to
    --          initialize a variable.

uses
    TCollection,MMgt,SortTools,TColStd
is 

   enumeration FormatType is     
    	SJIS,
	EUC,
	ANSI,
	GB
   end FormatType ;
    	---Purpose:
    	-- List of non ASCII format types which may be
    	-- converted into the Unicode 16 bits format type.
    	-- Use the functions provided by the
    	-- Resource_Unicode class to convert a string
    	-- from one of these non ASCII format to Unicode, and vice versa.

   class DataMapOfAsciiStringAsciiString instantiates
    	 DataMap from TCollection(AsciiString from TCollection,
	    	    	    	 AsciiString from TCollection,
	    	    	    	 AsciiString from TCollection) ;

   class DataMapOfAsciiStringExtendedString instantiates
    	 DataMap from TCollection(AsciiString from TCollection,
	    	    	    	  ExtendedString from TCollection,
	    	    	    	  AsciiString from TCollection) ;
	 
   class QuickSortOfArray1 instantiates
    	 QuickSort from SortTools(AsciiString from TCollection,
    	    	    	    	  Array1OfAsciiString from TColStd,
	    	    	    	  LexicalCompare from Resource) ;
				  
---Class:
   class LexicalCompare ;
   
   class Manager;
   ---Purpose: Defines a resource structure and its management methods.

   class Unicode;

   exception NoSuchResource inherits NoSuchObject from Standard;

end Resource;
