-- File:	QAOCC_OCC749Prs.cdl
-- Created:	Fri Sep 20 16:32:13 2002
-- Author:	Michael KUZMITCHEV
--		<mkv@russox>
---Copyright:	 Matra Datavision 2002

class OCC749Prs from QAOCC inherits InteractiveObject from AIS

uses
    PresentationManager3d from PrsMgr,
    Presentation          from Prs3d,
    Selection             from SelectMgr,
    Color                 from Quantity
    
is
    Create( reflection : Boolean from Standard;
    	    color      : Color from Quantity;
    	    color1      : Color from Quantity )
     returns mutable OCC749Prs from QAOCC;

    Compute(me                   : mutable;
            aPresentationManager : PresentationManager3d from PrsMgr;
            aPresentation        : mutable Presentation from Prs3d;
    	    aMode                : Integer from Standard = 0) 
    is redefined virtual protected;

    ComputeSelection(me          : mutable;
    	    	     aSelection  : mutable Selection from SelectMgr;
    	    	     aMode       : Integer from Standard)
    is redefined virtual protected; 

    SetReflection( me : mutable; reflection : Boolean from Standard );
    
    SetColor( me : mutable; color  : Color from Quantity;
    	    	    	    color1 : Color from Quantity );

fields
    myReflection   : Boolean from Standard;
    myColor1       : Color from Quantity;
    myColor2       : Color from Quantity;
end OCC749Prs;
