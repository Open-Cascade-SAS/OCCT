-- File:	QAMARTEC.cdl
-- Created:	Fri Oct 11 16:58:05 2002
-- Author:	Michael KUZMITCHEV
--		<mkv@russox>
---Copyright:	 Matra Datavision 2002

package QAMARTEC
     uses Draw
is
    
    Commands(DI : in out Interpretor from Draw);
end;
