-- Created on: 1993-04-23
-- Created by: Laurent BUCHARD
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


package ApproxInt

uses 
     Standard,TCollection,math,gp,TColStd,TColgp,
     IntImp,IntSurf,
     AppParCurves,StdFail,Approx,MMgt
     
is


    generic class WLine; -- Only on curves with ->NbPoles, ->IsNull and  ->Pole  Methods
    deferred class SvSurfaces;     
    generic class PrmPrmSvSurfaces,TheInt2S;
    generic class ImpPrmSvSurfaces,TheZerImpFunc;
    generic class MultiLine;
    generic class MultiLineTool;
    generic class Approx,ThePrmPrmSvSurfaces,
                         TheImpPrmSvSurfaces,
                         TheMultiLine,
                         TheMultiLineTool,
			 TheComputeLine,
                         TheComputeLineBezier;

end ApproxInt;
