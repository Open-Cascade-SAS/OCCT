-- Created on: 1997-02-12
-- Created by: Laurent BOURESCHE
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SurfPointConstRadInv from BRepBlend

inherits SurfPointFuncInv from Blend 

    ---Purpose: This function  is used  to find a  solution on  a done
    --          point   of   the curve when   using  SurfRstConsRad or
    --          CSConstRad...          
    --          The vector <X>  used in Value, Values and  Derivatives
    --          methods  has  to   be the  vector   of the  parametric
    --          coordinates w, U,  V where w is  the parameter  on the
    --          guide line, U,V   are the parametric coordinates of  a
    --          point on the partner surface.

uses
    Pnt      from gp,
    Vector   from math,
    Matrix   from math,
    HSurface from Adaptor3d,
    HCurve   from Adaptor3d


is
    Create(S : HSurface from Adaptor3d; C : HCurve from Adaptor3d)
    returns SurfPointConstRadInv from BRepBlend;
    	
    Set(me: in out; R: Real from Standard; Choix: Integer from Standard)
    is static;

    NbEquations(me)
    ---Purpose: returns 3.
    returns Integer from Standard;

    Value(me: in out; X: Vector; F: out Vector)
    ---Purpose: computes the values <F> of the Functions for the 
    --          variable <X>.
    --          Returns True if the computation was done successfully, 
    --          False otherwise.
    returns Boolean from Standard;
    
    Derivatives(me: in out; X: Vector; D: out Matrix)
    ---Purpose: returns the values <D> of the derivatives for the 
    --          variable <X>.
    --          Returns True if the computation was done successfully, 
    --          False otherwise.
    returns Boolean from Standard;
    
    Values(me: in out; X: Vector; F: out Vector; D: out Matrix)
    ---Purpose: returns the values <F> of the functions and the derivatives
    --          <D> for the variable <X>.
    --          Returns True if the computation was done successfully, 
    --          False otherwise.
    returns Boolean from Standard;

    Set(me: in out; P : Pnt from gp);
    ---Purpose: Set the Point on which a solution has to be found.

    GetTolerance(me; Tolerance: out Vector from math; Tol: Real from Standard);
    ---Purpose: Returns in the vector Tolerance the parametric tolerance
    --          for each of the 3 variables;
    --          Tol is the tolerance used in 3d space.

    GetBounds(me; InfBound,SupBound: out Vector from math);
    ---Purpose: Returns in the vector InfBound the lowest values allowed
    --          for each of the 3 variables.
    --          Returns in the vector SupBound the greatest values allowed
    --          for each of the 3 variables.

    IsSolution(me: in out; Sol: Vector from math; Tol: Real from Standard)
    ---Purpose: Returns Standard_True if Sol is a zero of the function.
    --          Tol is the tolerance used in 3d space.
    returns Boolean from Standard;

fields

    surf  : HSurface from Adaptor3d;
    curv  : HCurve   from Adaptor3d;
    point : Pnt      from gp;
    ray   : Real     from Standard;
    choix : Integer  from Standard;

end SurfPointConstRadInv;
