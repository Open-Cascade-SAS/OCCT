-- Created on: 1991-03-27
-- Created by: Michel CHAUVAT
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



package LProp

    ---Purpose: Handles local properties of curves and surfaces.
    --          Given a curve and a parameter value the following computations
    --          are available :
    --          - point,
    --          - derivatives,
    --          - tangent,
    --          - normal,
    --          - curvature,
    --          - centre of curvature,
    --          - Locals curvature's extremas,
    --          - Points of inflection,
    --          Given a surface and 2 parameters the following computations
    --          are available :
    --          - for each parameter:
    --            - derivatives,
    --            - tangent line,
    --            - centre of curvature,
    --          - point,
    --          - normal line,
    --          - maximum and minimum curvatures,
    --          - principal directions of curvature,
    --          - mean curvature,
    --          - Gaussian curvature.


    ---Level : Public. 
    --  All methods of all  classes will be public.

uses Standard, gp, math, TCollection, TColStd, GeomAbs

is

    enumeration Status is Undecided , Undefined, Defined, Computed;
    enumeration CIType is Inflection, MinCur   , MaxCur;
    	---Purpose:
    	-- Identifies the type of a particular point on a curve:
    	-- - LProp_Inflection: a point of inflection
    	-- - LProp_MinCur: a minimum of curvature
    	-- - LProp_MaxCur: a maximum of curvature.
        
    exception BadContinuity inherits Failure;
    exception NotDefined    inherits Failure;
    
    deferred generic class CurveTool;
        ---Purpose: The template class used in CLProps.
    deferred generic class SurfaceTool;
        ---Purpose: The template class used in SLProps.
    
    generic class CLProps;
    	---Purpose: Computation of local properties of a curve.
    generic class SLProps;
    	---Purpose: Computation of local properties of a surface.

							    
    class CurAndInf;	
    	---Purpose: Stores the parameters of a curve 2d or 3d corresponding
	--          to the curvature's extremas and the inflection's points.
    
    class AnalyticCurInf;
    	---Purpose: Computes the locals extremas of curvature of a gp curve.

    private generic class FuncCurExt;
    private generic class FuncCurNul;
    generic class NumericCurInf, FCurExt, FCurNul;    	
    	---Purpose: Computes the locals extremas of curvature and the 
    	--          inflections of a bounded curve in 2d.

    private class SequenceOfCIType instantiates Sequence from TCollection 
						        (CIType  from  LProp); 
    
end LProp;    
