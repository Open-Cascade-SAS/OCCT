-- Created on: 1993-09-22
-- Created by: Didier PIFFAULT
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package BRepMesh

        ---Purpose: Instantiated   package for the   class of packages

        ---Level : Advanced.  
        --  All methods of all  classes will be advanced.


uses    Standard,
        gp,
        Bnd,
        TColStd,
        TColgp,
        GCPnts,
        BRepAdaptor,
        BRepTopAdaptor,
        TCollection,
        MMgt,
        TopoDS,
        TopAbs,
        TopExp,
        TopTools,
        Poly,
        Geom2d,
        GeomAbs,
        GeomAdaptor,
        TopLoc,
        SortTools,
        Plugin

is
      imported DegreeOfFreedom from BRepMesh;
      imported Status from BRepMesh;
      imported FactoryError from BRepMesh;
      imported Vertex from BRepMesh;
      imported Edge from BRepMesh;
      imported Triangle from BRepMesh;
      imported Circle from BRepMesh;
      imported DiscretRoot from BRepMesh; 
      imported DiscretFactory from BRepMesh;
      --
      pointer PDiscretRoot to DiscretRoot from BRepMesh;
      
      imported ShapeTool from BRepMesh;
      imported Collections from BRepMesh;
      imported Delaun from BRepMesh;
      imported PairOfIndex from BRepMesh;
      imported CircleInspector from BRepMesh;
      imported VertexInspector from BRepMesh;
      imported WireInterferenceChecker from BRepMesh;
      imported EdgeChecker from BRepMesh;
      imported FaceChecker from BRepMesh;

      primitive PluginEntryType;

      imported SelectorOfDataStructureOfDelaun from BRepMesh;
      imported DataStructureOfDelaun from BRepMesh;
      imported CircleTool from BRepMesh;
      imported VertexTool from BRepMesh;
      imported BiPoint from BRepMesh;
      imported FastDiscretFace from BRepMesh;
      imported FastDiscret from BRepMesh;
      imported FaceAttribute from BRepMesh;
      imported Classifier from BRepMesh;
      imported WireChecker from BRepMesh;
      imported IncrementalMesh from BRepMesh;
      imported GeomTool from BRepMesh;
      imported PairOfPolygon from BRepMesh;

end BRepMesh;
