-- Created on: 1995-12-15
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class Face from BRepCheck inherits Result from BRepCheck

	---Purpose: 

uses Shape  from TopoDS,
     Face   from TopoDS,
     Status from BRepCheck,
     DataMapOfShapeListOfShape from TopTools

is

    Create(F: Face from TopoDS)
    
    	returns mutable Face from BRepCheck;


    InContext(me: mutable; ContextShape: Shape from TopoDS);
    


    Minimum(me: mutable);
    

    
    Blind(me: mutable);
    
    
    
    IntersectWires(me: mutable; Update: Boolean from Standard = Standard_False)
    
    	returns Status from BRepCheck
	is static;


    ClassifyWires(me: mutable; Update: Boolean from Standard = Standard_False)
    
    	returns Status from BRepCheck
	is static;



    OrientationOfWires(me: mutable; 
    	    	    	Update: Boolean from Standard = Standard_False)
    
    	returns Status from BRepCheck
	is static;


    SetUnorientable(me: mutable)
    
    	is static;


    IsUnorientable(me)
    
    	returns Boolean from Standard
	is static;

    GeometricControls(me)
    
    	returns Boolean from Standard
	is static;


    GeometricControls(me: mutable; B: Boolean from Standard)
    
	is static;



fields

    myIntdone : Boolean                   from Standard;
    myIntres  : Status                    from BRepCheck;
    myImbdone : Boolean                   from Standard;
    myImbres  : Status                    from BRepCheck;
    myOridone : Boolean                   from Standard;
    myOrires  : Status                    from BRepCheck;
    myMapImb  : DataMapOfShapeListOfShape from TopTools;
    myGctrl   : Boolean from Standard;

end Face;
