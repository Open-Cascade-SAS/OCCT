-- Created on: 1991-03-21
-- Created by: Philippe DAUTRY
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Circ2d2TanRad

from GccAna

	---Purpose: This class implements the algorithms used to 
	--          create 2d circles tangent to 2 
	--          points/lines/circles and with a given radius.
    	--          For each construction methods arguments are:
    	--            - Two Qualified elements for tangency constraints.
    	--            (for example EnclosedCirc if we want the 
    	--            solution inside the argument EnclosedCirc).
    	--            - Two Reals. One (Radius) for the radius and the 
    	--            other (Tolerance) for the tolerance.
    	--          Tolerance is only used for the limit cases.
    	--          For example : 
    	--          We want to create a circle inside a circle C1 and 
    	--          inside a circle C2 with a radius Radius and a 
    	--          tolerance Tolerance.
    	--          If we do not use Tolerance it is impossible to 
    	--          find a solution in the following case : C2 is 
    	--          inside C1 and there is no intersection point 
    	--          between the two circles.
    	--          With Tolerance it gives a solution if the lowest 
    	--          distance between C1 and C2 is lower than or equal
    	--          Tolerance.



uses Pnt2d           from gp,
     Circ2d          from gp,
     QualifiedLin    from GccEnt,
     QualifiedCirc   from GccEnt,
     Array1OfReal    from TColStd,
     Array1OfInteger from TColStd,
     Array1OfCirc2d  from TColgp,
     Array1OfPnt2d   from TColgp,
     Position         from GccEnt,
     Array1OfPosition from GccEnt

raises NegativeValue     from Standard,
       OutOfRange        from Standard,
       BadQualifier      from GccEnt,
       NotDone           from StdFail

is

Create(Qualified1 : QualifiedCirc from GccEnt  ;
       Qualified2 : QualifiedCirc from GccEnt  ;
       Radius     : Real          from Standard;
       Tolerance  : Real          from Standard) returns Circ2d2TanRad
	---Purpose: This method implements the algorithms used to 
	--          create 2d circles TANgent to two 2d circle with a 
	--          radius of Radius.
raises NegativeValue, BadQualifier;
	---Purpose: It raises NegativeValue if Radius is lower than zero.

Create(Qualified1 : QualifiedCirc from GccEnt  ;
       Qualified2 : QualifiedLin  from GccEnt  ;
       Radius     : Real          from Standard;
       Tolerance  : Real          from Standard) returns Circ2d2TanRad
	---Purpose: This method implements the algorithms used to 
	--          create 2d circles TANgent to a 2d circle and a 2d line
	--          with a radius of Radius.
raises NegativeValue, BadQualifier;
	---Purpose: It raises NegativeValue if Radius is lower than zero.

Create(Qualified1 : QualifiedCirc from GccEnt  ;
       Point2     : Pnt2d         from gp      ;
       Radius     : Real          from Standard;
       Tolerance  : Real          from Standard) returns Circ2d2TanRad
	---Purpose: This method implements the algorithms used to 
	--          create 2d circles TANgent to a 2d circle and a point
	--          with a radius of Radius.
raises NegativeValue, BadQualifier;
	---Purpose: It raises NegativeValue if Radius is lower than zero.

Create(Qualified1 : QualifiedLin from GccEnt  ;
       Point2     : Pnt2d        from gp      ;
       Radius     : Real         from Standard;
       Tolerance  : Real         from Standard) returns Circ2d2TanRad
	---Purpose: This method implements the algorithms used to 
	--          create 2d circles TANgent to a 2d line and a point
	--          with a radius of Radius.
raises NegativeValue, BadQualifier;
	---Purpose: It raises NegativeValue if Radius is lower than zero.

Create(Qualified1 : QualifiedLin from GccEnt  ;
       Qualified2 : QualifiedLin from GccEnt  ;
       Radius     : Real         from Standard;
       Tolerance  : Real         from Standard) returns Circ2d2TanRad
	---Purpose: This method implements the algorithms used to 
	--          create 2d circles TANgent to two 2d lines
	--          with a radius of Radius.
raises NegativeValue, BadQualifier;
	---Purpose: It raises NegativeValue if Radius is lower than zero.

Create(Point1     : Pnt2d   from gp      ;
       Point2     : Pnt2d   from gp      ;
       Radius     : Real    from Standard;
       Tolerance  : Real    from Standard) returns Circ2d2TanRad
	---Purpose: This method implements the algorithms used to 
	--          create 2d circles passing through two points with a 
	--          radius of Radius.
raises NegativeValue;
	---Purpose: It raises NegativeValue if Radius is lower than zero.

-- -- ....................................................................

IsDone(me) returns Boolean from Standard
is static;
    	---Purpose: This method returns True if the algorithm succeeded.
    	-- Note: IsDone protects against a failure arising from a
    	-- more internal intersection algorithm, which has reached its numeric limits.
    
NbSolutions(me) returns Integer from Standard
    	---Purpose: This method returns the number of circles, representing solutions computed by this algorithm.
    	-- Exceptions
    	-- StdFail_NotDone if the construction fails. of solutions.
raises NotDone
is static;

ThisSolution(me                           ;  
    	     Index : Integer from Standard) returns Circ2d from gp
    ---Purpose: Returns the solution number Index.
    --          Be careful: the Index is only a way to get all the 
    --          solutions, but is not associated to those outside the context
    --          of the algorithm-object. Raises OutOfRange exception if Index is greater 
    --          than the number of solutions.
    --          It raises NotDone if the construction algorithm did not 
    --          succeed.

raises OutOfRange, NotDone
is static;
    

WhichQualifier(me                                  ;
    	       Index   :     Integer  from Standard;
	       Qualif1 : out Position from GccEnt  ;
	       Qualif2 : out Position from GccEnt  )
raises OutOfRange, NotDone
is static;
    ---Purpose: Returns the information about the qualifiers of
    --          the tangency arguments concerning the solution number Index.
    --          It returns the real qualifiers (the qualifiers given to the 
    --          constructor method in case of enclosed, enclosing and outside 
    --          and the qualifiers computedin case of unqualified).

Tangency1(me                                       ;
          Index         :     Integer from Standard;
          ParSol        : out Real    from Standard;
          ParArg        : out Real    from Standard;
          PntSol        : out Pnt2d   from gp       )
    ---Purpose: Returns information about the tangency point between the 
    -- result number Index and the first argument.
    -- ParSol is the intrinsic parameter of the point PntSol on the solution.
    -- ParArg is the intrinsic parameter of the point PntSol on the first
    -- argument. Raises OutOfRange if Index is greater than the number 
    --          of solutions.
    --          It raises NotDone if the construction algorithm did not succeed
raises OutOfRange, NotDone
is static;
    

Tangency2(me                                       ;
          Index         :     Integer from Standard;
          ParSol,ParArg : out Real    from Standard;
          PntSol        : out Pnt2d   from gp      )
    ---Purpose: Returns information about the tangency point between the 
    --          result number Index and the second argument.
    --          ParSol is the intrinsic parameter of the point PntSol on 
    --          the solution.
    --          ParArg is the intrinsic parameter of the point PntArg on 
    --          the second argument. Raises OutOfRange if Index is greater than the number 
    --          of solutions.
    --          It raises NotDone if the construction algorithm did not succeed.
raises OutOfRange, NotDone
is static;
   

IsTheSame1(me                           ;
           Index : Integer from Standard) returns Boolean from Standard
    ---Purpose: Returns True if the solution number Index is equal to 
    --          the first argument. Raises OutOfRange if Index is greater than the number 
    --          of solutions.
    --          It raises NotDone if the construction algorithm did not 
    --          succeed.
raises OutOfRange, NotDone
is static;
 

IsTheSame2(me                           ;
           Index : Integer from Standard) returns Boolean from Standard
    ---Purpose: Returns True if the solution number Index is equal to 
    --          the second argument. Raises OutOfRange if Index is greater than the number 
    --          of solutions.
    --          It raises NotDone if the construction algorithm did not  succeed.
raises OutOfRange, NotDone
is static;
  

fields

    WellDone : Boolean from Standard;
    ---Purpose: True if the algorithm succeeded.

    qualifier1 : Array1OfPosition from GccEnt;
    -- The qualifiers of the first argument.

    qualifier2 : Array1OfPosition from GccEnt;
    -- The qualifiers of the second argument.

    TheSame1 : Array1OfInteger from TColStd;
    ---Purpose: 1 if the solution and the first argument are the same 
    --          (2 circles).
    --          If R1 is the radius of the first argument and Rsol the radius 
    --          of the solution and dist the distance between the two centers,
    --          we consider the two circles are identical if R1+dist-Rsol is 
    --          less than Tolerance.
    --          0 in the other cases.

    TheSame2 : Array1OfInteger from TColStd;
    ---Purpose: 1 if the solution and the second argument are the same 
    --          (2 circles).
    --          If R2 is the radius of the second argument and Rsol the radius 
    --          of the solution and dist the distance between the two centers,
    --          we consider the two circles are identical if R2+dist-Rsol is 
    --          less than Tolerance.
    --          0 in the other cases.

    NbrSol   : Integer from Standard;
    ---Purpose: The number of possible solutions.

    cirsol   : Array1OfCirc2d from TColgp;
    ---Purpose: The solutions.

    pnttg1sol   : Array1OfPnt2d from TColgp;
    ---Purpose: The tangency point between the solution and the first 
    --          argument on the solution.

    pnttg2sol   : Array1OfPnt2d from TColgp;
    ---Purpose: The tangency point between the solution and the second 
    --          argument on the solution.

    par1sol   : Array1OfReal from TColStd;
    ---Purpose: The parameter of the tangency point between the solution 
    --          and the first argument on the solution.

    par2sol   : Array1OfReal from TColStd;
    ---Purpose: The parameter of the tangency point between the solution 
    --          and the second argument on the solution.

    pararg1   : Array1OfReal from TColStd;
    ---Purpose: The parameter of the tangency point between the solution 
    --          and the first argument on the first argument.

    pararg2   : Array1OfReal from TColStd;
    ---Purpose: The parameter of the tangency point between the solution 
    --          and the second argument on the second argument.

end Circ2d2TanRad;
