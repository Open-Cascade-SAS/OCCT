-- Created on: 1993-03-10
-- Created by: Philippe DAUTRY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



deferred class BoundedSurface from Geom inherits Surface from Geom


        ---Purpose : The root class for bounded surfaces in 3D space. A
    	-- bounded surface is defined by a rectangle in its 2D parametric space, i.e.
    	-- - its u parameter, which ranges between two finite
    	--   values u0 and u1, referred to as "First u
    	--   parameter" and "Last u parameter" respectively, and
    	-- - its v parameter, which ranges between two finite
    	--   values v0 and v1, referred to as "First v
    	--   parameter" and the "Last v parameter" respectively.
    	--   The surface is limited by four curves which are the
    	-- boundaries of the surface:
    	-- - its u0 and u1 isoparametric curves in the u parametric direction, and
    	-- - its v0 and v1 isoparametric curves in the v parametric direction.
    	-- A bounded surface is finite.
    	-- The common behavior of all bounded surfaces is
    	-- described by the Geom_Surface class.
    	-- The Geom package provides three concrete
    	-- implementations of bounded surfaces:
    	-- - Geom_BezierSurface,
    	-- - Geom_BSplineSurface, and
    	-- - Geom_RectangularTrimmedSurface.
    	--  The first two of these implement well known
    	-- mathematical definitions of complex surfaces, the third
    	-- trims a surface using four isoparametric curves, i.e. it
    	-- limits the variation of its parameters to a rectangle in
    	-- 2D parametric space.

is


end;



