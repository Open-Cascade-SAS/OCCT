-- Created on: 1999-06-10
-- Created by: Vladislav ROMASHKO
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package TFunction 
    --- Purpose: Function attributes separate data from
    -- algorithms. Each function contains the ID of a function driver.
uses  

    Standard, 
    TCollection,  
    TColStd,
    TDF, 
    TDataStd
 
is 
  
    enumeration ExecutionStatus is
    	ES_WrongDefinition,
	ES_NotExecuted,
	ES_Executing,
	ES_Succeeded,
	ES_Failed;

    deferred class Driver;         

    class DriverTable;   

    class Logbook;

    class DataMapOfGUIDDriver
    instantiates DataMap from TCollection(GUID   from Standard, 
	    	 		       	  Driver from TFunction, 
				          GUID   from Standard);
    class Array1OfDataMapOfGUIDDriver
    instantiates Array1 from TCollection(DataMapOfGUIDDriver from TFunction);
    class HArray1OfDataMapOfGUIDDriver
    instantiates HArray1 from TCollection(DataMapOfGUIDDriver from TFunction,
    	    	    	    	    	  Array1OfDataMapOfGUIDDriver from TFunction);

    class Function; 
    class GraphNode;
    class Scope;

    class IFunction;
    class Iterator;

    class DataMapOfLabelListOfLabel
    instantiates DataMap from TCollection(Label          from TDF, 
	    	 		       	  LabelList      from TDF, 
				          LabelMapHasher from TDF);     
    class DoubleMapOfIntegerLabel
    instantiates DoubleMap from TCollection(Integer from Standard,
    	    	    	    	    	    Label from TDF,
					    MapIntegerHasher from TColStd,
					    LabelMapHasher from TDF);

end TFunction;    
