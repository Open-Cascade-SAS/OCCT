-- Created on: 2001-09-10
-- Created by: Sergey KUUL
-- Copyright (c) 2001-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MapContainer from Transfer inherits TShared from MMgt

	---Purpose: 

uses

    DataMapOfTransientTransient from TColStd

is

    Create returns mutable MapContainer from Transfer;
     
    SetMapObjects(me : mutable; theMapObjects : in out DataMapOfTransientTransient from TColStd);
    	---Purposes:Set map already translated geometry objects.
	
    GetMapObjects(me: mutable) returns DataMapOfTransientTransient from TColStd;
    	---Purposes:Get map already translated geometry objects.
    	---C++:return &
fields

  myMapObj           : DataMapOfTransientTransient from TColStd;
  
end MapContainer;
