-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class CsgSelect from StepShape 

    -- inherits SelectType from StepData

	-- <CsgSelect> is an EXPRESS Select Type construct translation.
	-- it gathers : BooleanResult, CsgPrimitive

uses

	BooleanResult,
	CsgPrimitive
is

	Create returns CsgSelect;
	---Purpose : Returns a CsgSelect SelectType

    	SetTypeOfContent(me : in out; aTypeOfContent : Integer);

	TypeOfContent(me) returns Integer;
	--        1 -> BooleanResult
	--        2 -> CsgPrimitive
	--        0 else
	
	BooleanResult (me) returns any BooleanResult;
	---Purpose : returns Value as a BooleanResult (Null if another type)

    	SetBooleanResult (me : in out;aBooleanResult : BooleanResult from StepShape);
	
	CsgPrimitive (me) returns CsgPrimitive;
	---Purpose : returns Value as a CsgPrimitive (Null if another type)

    	SetCsgPrimitive (me : in out; aCsgPrimitive : CsgPrimitive from StepShape);
	
fields

    theBooleanResult : BooleanResult from StepShape;
    theCsgPrimitive  : CsgPrimitive  from StepShape;  -- a Select Type
    theTypeOfContent : Integer       from Standard;

end CsgSelect;

