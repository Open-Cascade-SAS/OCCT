-- Created by: NW,JPB,CAL
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Light from Visual3d inherits TShared

	---Version:

	---Purpose: This class defines and updates light sources.
	--	    There is no limit to the number of light sources defined.
	--	    Only the number of active sources is limited.
	--
	--	    TypeOfLightSource = TOLS_AMBIENT
	--				TOLS_DIRECTIONAL
	--				TOLS_POSITIONAL
	--				TOLS_SPOT
	--
	--	    Angle is a radian value.
	--	    Concentration, Attenuation are in the [0,1] interval.
	--

	---Keywords: Light, View, Context, Ambient, Directional, Positional,
	--	     Spot, Angle, Concentration, Attenuation, Color, Shading

	---Warning:
	---References:

uses

  Color  from Quantity,
  CLight from Graphic3d,
  Vector from Graphic3d,
  Vertex from Graphic3d,
  TypeOfLightSource from Visual3d

raises

  LightDefinitionError from Visual3d

is

	Create
		returns Light from Visual3d;
	---Level: Public
	---Purpose: Creates a light from default values.
	--	    Light sources are created in a visualiser
	--	    and are activated in one of its views.
	--
	--	    Type	= TOLS_AMBIENT
	--	    Color	= WHITE

	Create ( Color		: Color from Quantity )
		returns Light from Visual3d;
	---Level: Public
	---Purpose: Creates an AMBIENT light source.
	--	    Light sources are created in a visualiser
	--	    and are activated in one of its views.

    Create ( theColor       : Color from Quantity;
             theDirection   : Vector from Graphic3d;
             theHeadlight   : Boolean from Standard = Standard_False;
             theSmoothAngle : Real from Standard = 0.0;
             theIntensity   : Real from Standard = 1.0 )
    returns Light from Visual3d
    ---Level: Public
    ---Purpose: Creates a DIRECTIONAL light source.
    --      Light sources are created in a visualiser
    --      and are activated in one of its views.
    --  Warning: Raises LightDefinitionError if <Direction> is null.
    raises LightDefinitionError;

    Create ( theColor        : Color from Quantity;
             thePosition     : Vertex from Graphic3d;
             theFact1        : Real from Standard;
             theFact2        : Real from Standard;
             theSmoothRadius : Real from Standard = 0.0;
             theIntensity   : Real from Standard = 1.0 )
    returns Light from Visual3d
    ---Level: Public
    ---Purpose: Creates a POSITIONAL light source.
    --      Light sources are created in a visualiser
    --      and are activated in one of its views.
    --  Warning: Raises LightDefinitionError 
    --      if <Fact1> and <Fact2> are null.
    --      if <Fact1> is a negative value or greater than 1.0.
    --      if <Fact2> is a negative value or greater than 1.0.
    raises LightDefinitionError;

	Create ( Color		: Color from Quantity;
		 Position	: Vertex from Graphic3d;
		 Direction	: Vector from Graphic3d;
		 Concentration	: Real from Standard;
		 Fact1, Fact2	: Real from Standard;
		 AngleCone	: Real from Standard )
		returns Light from Visual3d
	---Level: Public
	---Purpose: Creates a SPOT light source.
	--	    Light sources are created in a visualiser
	--	    and are activated in one of its views.
	--	    <Concentration> specifies the intensity distribution of 
	--	    the light.
	--	    <AngleCone> specifies the angle (radians) of the cone 
	--	    created by the spot.
	-- 	    the global attenuation is equal :
	--	    1 / (Fact1 + Fact2 * (norm(ObjectPosition - LightPosition)))
	--  Warning: Raises LightDefinitionError
	--	    if <Direction> is null.
	--	    if <Concentration> is a negative value or greater than 1.0.
	--	    if <Fact1> and <Fact2> are null.
	--	    if <Fact1> is a negative value or greater than 1.0.
	--	    if <Fact2> is a negative value or greater than 1.0.
	--	    if <AngleCone> is a negative value or greater than PI/2.
	raises LightDefinitionError;

	---------------------------------------------------
	-- Category: Methods to modify the class definition
	---------------------------------------------------

	SetAngle ( me		: mutable;
		   AngleCone	: Real from Standard )
	---Level: Public
	---Purpose: Modifies the angle (radians) of the cone created by the spot.
	--	    Works only on TOLS_SPOT lights. 
	--  Category: Methods to modify the class definition
	--  Warning: Raises LightDefinitionError
	--	    if the type of the light is not TOLS_SPOT.
	--	    if <AngleCone> is a negative value or greater than PI/2.
	raises LightDefinitionError is static;

	SetAttenuation1 ( me	: mutable;
			  Fact1	: Real from Standard )
	---Level: Public
	---Purpose: Modifies the attenuation factor of the light.
	--	    Works only on the TOLS_POSITIONAL and TOLS_SPOT lights.
	--  Category: Methods to modify the class definition
	--  Warning: Raises LightDefinitionError
	--	    if the type of the light is not TOLS_SPOT or TOLS_POSITIONAL.
	--	    if <Fact1> is a negative value or greater than 1.0.
	raises LightDefinitionError is static;

	SetAttenuation2 ( me	: mutable;
			  Fact2	: Real from Standard )
	---Level: Public
	---Purpose: Modifies the attenuation factor of the light.
	--	    Works only on the TOLS_POSITIONAL and TOLS_SPOT lights.
	--  Category: Methods to modify the class definition
	--  Warning: Raises LightDefinitionError
	--	    if the type of the light is not TOLS_POSITIONAL or TOLS_SPOT.
	--	    if <Fact2> is a negative value or greater than 1.0..
	raises LightDefinitionError is static;

	SetColor ( me		: mutable;
		   Color	: Color from Quantity )
		is static;
	---Level: Public
	---Purpose: Modifies the colour of the light.
	---Category: Methods to modify the class definition

	SetConcentration ( me			: mutable;
			   Concentration	: Real from Standard )
	---Level: Public
	---Purpose: Modifies the intensity distribution of the light.
	--	    Works only on the TOLS_SPOT lights.
	--  Category: Methods to modify the class definition
	--  Warning: Raises LightDefinitionError
	--	    if the type of the light is not TOLS_SPOT.
	--	    if <Concentration> is a negative value or greater than 1.0.
	raises LightDefinitionError is static;

	SetDirection ( me		: mutable;
		       Direction	: Vector from Graphic3d )
	---Level: Public
	---Purpose: Modifies the light direction.
	--	    Works only on the TOLS_DIRECTIONAL and TOLS_SPOT lights.
	--	    Default z
	--  Category: Methods to modify the class definition
	--  Warning: Raises LightDefinitionError
	--	    if the type of the light is not TOLS_DIRECTIONAL
	--	    or TOLS_SPOT.
	--	    if <Direction> is null.
	raises LightDefinitionError is static;

	SetPosition ( me	: mutable;
		      Position	: Vertex from Graphic3d )
	---Level: Public
	---Purpose: Modifies the position of the light.
	--	    Works only on the TOLS_POSITIONAL and TOLS_SPOT lights.
	--  Category: Methods to modify the class definition
	--  Warning: Raises LightDefinitionError 
	--	    if the type of the light is not TOLS_POSITIONAL or TOLS_SPOT.
	raises LightDefinitionError is static;

    SetSmoothAngle ( me       : mutable;
                     theValue : Real from Standard )
    ---Level: Public
    ---Purpose: Modifies the smoothing angle (in radians) of
    --          DIRECTIONAL light source.
    --  Category: Methods to modify the class definition
    --  Warning: Raises LightDefinitionError
    --      if the type of the light is not TOLS_DIRECTIONAL
    --      if <Value> is negative or greater than PI / 2.
    raises LightDefinitionError is static;

    SetSmoothRadius ( me       : mutable;
                      theValue : Real from Standard )
    ---Level: Public
    ---Purpose: Modifies the smoothing radius of
    --          POSITIONAL light source.
    --  Category: Methods to modify the class definition
    --  Warning: Raises LightDefinitionError
    --      if the type of the light is not TOLS_POSITIONAL
    --      if <Value> is negative.
    raises LightDefinitionError is static;

    SetIntensity ( me       : mutable;
                   theValue : Real from Standard )
    ---Level: Public
    ---Purpose: Modifies the intensity of light source.
    --  Category: Methods to modify the class definition
    --  Warning: Raises LightDefinitionError
    --      if <Value> is negative or equal to zero.
    raises LightDefinitionError is static;

    Intensity ( me ) returns Real from Standard is static;
    ---Level: Public
    ---Purpose: returns the intensity of light source

    Smoothness ( me ) returns Real from Standard is static;
    ---Level: Public
    ---Purpose: returns the smoothness of light source

	----------------------------
	-- Category: Inquire methods
	----------------------------

  Headlight ( me )
  returns  Boolean  from  Standard  is  static;
  ---Level: Public
  ---Purpose:  Returns the headlight  state of the light <me>
  ---Category: Inquire methods

  SetHeadlight( me : mutable; theValue : Boolean from Standard ) is static;
  ---Level: Public
  ---Purpose: Setup headlight flag.

	Color ( me )
		returns Color from Quantity is static;
	---Level: Public
	---Purpose: Returns the colour of the light <me>.
	---Category: Inquire methods

	LightType ( me )
		returns TypeOfLightSource from Visual3d is static;
	---Level: Public
	---Purpose: Returns the light type of <me>.
	--
	--	    TypeOfLightSource = TOLS_AMBIENT
	--				TOLS_DIRECTIONAL
	--				TOLS_POSITIONAL
	--				TOLS_SPOT
	--
	---Category: Inquire methods

	Values ( me;
		 Color		: out Color from Quantity )
	---Level: Public
	---Purpose: Returns the definition of <me> if <me> is
	--	    a light source of the TOLS_AMBIENT type.
	--  Category: Inquire methods
	--  Warning: Raises LightDefinitionError 
	--	    if the type of the light is not TOLS_AMBIENT.
	raises LightDefinitionError is static;

	Values ( me;
		 Color		: out Color from Quantity;
		 Direction	: out Vector from Graphic3d )
	---Level: Public
	---Purpose: Returns the definition of <me> if <me> is
	--	    a light source of the TOLS_DIRECTIONAL type.
	--  Category: Inquire methods
	--  Warning: Raises LightDefinitionError 
	--	    if the type of the light is not TOLS_DIRECTIONAL.
	raises LightDefinitionError is static;

	Values ( me;
		 Color		: out Color from Quantity;
		 Position	: out Vertex from Graphic3d;
		 Fact1,Fact2	: out Real from Standard )
	---Level: Public
	---Purpose: Returns the definition of <me> if <me> is
	--	    a light source of the TOLS_POSITIONAL type.
	--  Category: Inquire methods
	--  Warning: Raises LightDefinitionError 
	--	    if the type of the light is not TOLS_POSITIONAL.
	raises LightDefinitionError is static;

	Values ( me;
		 Color		: out Color from Quantity;
		 Position	: out Vertex from Graphic3d;
		 Direction	: out Vector from Graphic3d;
		 Concentration	: out Real from Standard;
		 Fact1,Fact2	: out Real from Standard;
		 AngleCone	: out Real from Standard )
	---Level: Public
	---Purpose: Returns the definition of <me> if <me> is
	--	    a light source of the TOLS_SPOT type.
	--  Category: Inquire methods
	--  Warning: Raises LightDefinitionError 
	--	    if the type of the light is not TOLS_SPOT.
	raises LightDefinitionError is static;

  CLight ( me )
  returns CLight from Graphic3d
  is static;
  ---C++: return const &
  ---Level: Public
  ---Purpose: Returns the light defintion.
  ---Category: Inquire methods

	--------------------------
	-- Category: Class methods
	--------------------------

	IsValid ( myclass;
		  AAngle	: Real from Standard )
		returns Boolean from Standard
		is private;
	---Level: Internal
	---Purpose: Returns True if <AAngle> is a valid
	--	    spot light spread angle.
	---Category: Private methods

--

fields

  -- the associated C structure
  myCLight : CLight from Graphic3d;

friends

	class View from Visual3d

end Light;
