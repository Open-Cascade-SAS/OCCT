-- Created on: 1995-02-10
-- Created by: Mister rmi
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class DefaultMap from V2d

     ---Purpose:  Modifies class definition.
        
uses
    GenericColorMap, TypeMap, WidthMap, FontMap, MarkMap from Aspect
is

    ColorMap(myclass) 
    ---Purpose: Returns a indexed color map with the following color
    --          White, black, red, green, blue1 , yellow, sienna, orange2 
    --          lightgray,lightseagreen,gray60,gray70. The index are 1 to 12.
    returns GenericColorMap from Aspect;


    TypeMap(myclass)
    ---Purpose: Returns a indexed type map with the following line types
    --          SOLID, DASH, DOT, DOTDASH. The index are 1 to 4.
    returns TypeMap from Aspect;
    
    WidthMap(myclass)
    ---Purpose: Returns a indexed width map with the following width
    --          0.0001, 0.0006, 0.001, 0.003. The index are 1 to 4.
    returns WidthMap from Aspect;
    
    FontMap(myclass)
    ---Purpose: Returns a indexed font map with the following font
    --          "Courier-Bold" 0.01 0.0
    --          "Helvetica-Bold" 0.01 0.2
    --          "-adobe-helvetica-medium-r-normal--12-120-75-75-p-67-iso8859-1" 0.003 0.0
    --          The index are 1 to 2.
    returns FontMap from Aspect;
    

    MarkMap(myclass)
    ---Purpose: Returns a indexed font map with the following width
    --          Point,Plus,Star,O,X,O_Point,O_Plus,O_STAR,O_X
    --          BALL,RING1,RING2,RING3
    returns MarkMap from Aspect;
   
end DefaultMap from V2d;
