-- Created on: 1991-04-25
-- Created by: Arnaud BOUZY
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Segment3D from Draw inherits Drawable3D from Draw

	---Purpose: 

uses Pnt from gp,
    Color from Draw,
    Display from Draw

is

    Create(p1,p2 : Pnt; col : Color)
    returns mutable Segment3D;
    
    DrawOn(me; dis : in out Display);
    
    First(me) returns Pnt from gp
	---C++: return const&
    is static;

    First(me : mutable; P : Pnt from gp)
    is static;

    Last(me) returns Pnt from gp
	---C++: return const&
    is static;

    Last(me : mutable; P : Pnt from gp)
    is static;

fields

    myFirst : Pnt;
    myLast  : Pnt;
    myColor : Color;
    
end Segment3D;
