-- Created on: 1993-06-11
-- Created by: Jean-Louis FRENKEL
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ArrowAspect from Prs3d inherits BasicAspect from Prs3d
    	---Purpose: A framework for displaying arrows in representations
    	-- of dimensions and relations.
uses
    Length from Quantity,
    PlaneAngle from Quantity,
    NameOfColor from Quantity,
    Color       from Quantity,
    AspectLine3d from Graphic3d
    
raises
    InvalidAngle from Prs3d
    
is
    Create returns ArrowAspect from Prs3d;
    	---Purpose: Constructs an empty framework for displaying arrows
    	-- in representations of lengths. The lengths displayed
    	-- are either on their own or in chamfers, fillets,
    	-- diameters and radii.    

    Create (anAngle: PlaneAngle from Quantity; aLength: Length from Quantity)
    returns ArrowAspect from Prs3d;
    	--- Purpose: Constructs a framework to display an arrow with a
    	-- shaft of the length aLength and having a head with
    	-- sides at the angle anAngle from each other.   

    Create( theAspect: AspectLine3d from Graphic3d )
    returns ArrowAspect from Prs3d;
        
    SetAngle(me: mutable; anAngle: PlaneAngle from Quantity)
    	---Purpose: defines the angle of the arrows.
    raises InvalidAngle from Prs3d
    is static;
    
    Angle(me) returns PlaneAngle from Quantity
    	---Purpose: returns the current value of the angle used when drawing an arrow.
    is static;
    
    SetLength(me: mutable; aLength: Length from Quantity)
	---Purpose: defines the length of the arrows.
    is static;
    
    Length(me) returns Length from Quantity
	---Purpose: returns the current value of the length used when drawing an arrow.
    is static;

    SetColor(me: mutable; aColor:  Color  from  Quantity);

    SetColor(me: mutable; aColor:  NameOfColor  from  Quantity);

    Aspect(me) returns AspectLine3d  from  Graphic3d;

    SetAspect( me: mutable; theAspect: AspectLine3d from Graphic3d );

fields
	    myArrowAspect: AspectLine3d  from  Graphic3d;
	    myAngle: PlaneAngle from Quantity;
	    myLength: Length from Quantity;

end ArrowAspect from Prs3d;
