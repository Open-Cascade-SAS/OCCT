-- Created on: 1993-05-10
-- Created by: Christian CAILLET
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class GeneralModule  from IGESSolid     inherits  GeneralModule  from IGESData

    ---Purpose : Definition of General Services for IGESSolid (specific part)
    --           This Services comprise : Shared & Implied Lists, Copy, Check

uses OStream,
     Check, ShareTool, EntityIterator, CopyTool,
     IGESEntity, DirChecker

is

    Create returns mutable GeneralModule from IGESSolid;
    ---Purpose : Creates a GeneralModule from IGESSolid and puts it into GeneralLib

    OwnSharedCase  (me; CN : Integer; ent : IGESEntity;
    	    	    iter : in out EntityIterator);
    ---Purpose : Lists the Entities shared by a given IGESEntity <ent>, from
    --           its specific parameters : specific for each type

    DirChecker (me; CN : Integer; ent : IGESEntity) returns DirChecker;
    ---Purpose : Returns a DirChecker, specific for each type of Entity
    --           (identified by its Case Number) : this DirChecker defines
    --           constraints which must be respected by the DirectoryPart

    OwnCheckCase (me; CN : Integer; ent : IGESEntity; shares : ShareTool;
    	          ach    : in out Check);
    ---Purpose : Performs Specific Semantic Check for each type of Entity


    NewVoid (me; CN : Integer; entto : out mutable Transient)
    	returns Boolean;
    ---Purpose : Specific creation of a new void entity

    OwnCopyCase (me; CN : Integer;
    	         entfrom : IGESEntity; entto : mutable IGESEntity;
    	         TC : in out CopyTool);
    ---Purpose : Copies parameters which are specific of each Type of Entity

    CategoryNumber (me; CN : Integer; ent : Transient; shares : ShareTool)
    	returns Integer  is redefined;
    ---Purpose : Returns a category number which characterizes an entity
    --           Shape for all

end GeneralModule;
