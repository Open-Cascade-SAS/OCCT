-- Created by: NW,JPB,CAL
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class VertexC from Graphic3d inherits Vertex from Graphic3d

	---Version:

	---Purpose: This class allows the creation and update of a point
	--	    with a colour value.

	---Keywords: Vertex, Color, Coordinate, Point

	---Warning:
	---References:

uses

	Color	from Quantity
    	---Purpose: Returns the color of this point.
is

	Create
		returns VertexC from Graphic3d;
    	---Purpose: Constructs an empty point
        
	Create ( AX, AY ,AZ	: Real from Standard;
		 AColor		: Color from Quantity )
		returns VertexC from Graphic3d;
	---Level: Public
	---Purpose: Creates a point with coordinates <AX>, <AY>, <AZ> and
	--	    with colour <AColor>.

	Create ( APoint	: Vertex from Graphic3d;
		 AColor	: Color from Quantity )
		returns VertexC from Graphic3d;
	---Level: Public
	---Purpose: Creates a point situated in <APoint> and
	--	    for which the colour is <AColor>.

	---------------------------------------------------
	-- Category: Methods to modify the class definition
	---------------------------------------------------

	SetColor ( me		: in out;
		   ColorNew	: Color from Quantity )
		is static;
	---Level: Public
	---Purpose: Modifies the colour of the point <me>.
	---Category: Methods to modify the class definition

	----------------------------
	-- Category: Inquire methods
	----------------------------

	Color ( me )
		returns Color from Quantity
		is static;
	---Level: Public
	---Purpose: Returns the colour of the point <me>.
	---Category: Inquire methods

--

fields

--
-- Class	:	Graphic3d_VertexC
--
-- Purpose	:	Declaration of variables specific to points
--
-- Reminder	:	a point is defined by its coordinates and its colour
--

	-- the colour of a point
	MyColor		:	Color from Quantity;

end VertexC;
