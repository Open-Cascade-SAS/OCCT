-- Created on: 1998-03-26
-- Created by: # Andre LIEUTIER
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class FreeGtoCConstraint from Plate
---Purpose: define a G1, G2 or G3 constraint on the Plate using weaker
--          constraint than GtoCConstraint 
--          

uses 
 XY from gp, 
 XYZ from gp, 
 D1 from Plate, 
 D2 from Plate, 
 D3 from Plate, 
 PinpointConstraint from Plate,
 LinearScalarConstraint from Plate

is
    Create(point2d : XY ; D1S , D1T : D1 from Plate; 
    IncrementalLoad:  Real  =1.0; orientation:  Integer  =  0   ) returns FreeGtoCConstraint;
    -- G1 constraint:   
    -- D1S : first  derivative of  S, the surface we want to  correct 
    -- D1T : first derivative of the reference surface


    Create(point2d : XY from gp; D1S , D1T : D1 from Plate;
       D2S, D2T : D2 from Plate; 
    IncrementalLoad:  Real  =1.0; orientation:  Integer  =  0   ) returns FreeGtoCConstraint;
    -- G2 constraint:   
    -- D1S : first  derivative of  S, the surface we want to  correct 
    -- D1T : first derivative of the reference surface
    -- D2S : second derivative of  S, the surface we want to  correct 
    -- D2T : second derivative of the reference surface

    Create(point2d : XY from gp; D1S , D1T : D1 from Plate;
       D2S, D2T : D2 from Plate;
       D3S, D3T : D3 from Plate; 
    IncrementalLoad:  Real  =1.0; orientation:  Integer  =  0   ) returns FreeGtoCConstraint;
    -- G3 constraint:   
    -- D1S : first  derivative of  S, the surface we want to  correct 
    -- D1T : first derivative of the reference surface
    -- D2S : second derivative of  S, the surface we want to  correct 
    -- D2T : second derivative of the reference surface
    -- D3S : third derivative of  S, the surface we want to  correct 
    -- D3T : third derivative of the reference surface

    -- Accessors :
    nb_PPC(me) returns Integer;
    ---C++: inline 
    ---C++: return const &
          
    GetPPC(me;  Index:  Integer) returns PinpointConstraint;
    --	"C style" Index :  Index : 0 --> nb_PPC-1
    ---C++: inline 
    ---C++: return const &
          
    nb_LSC(me) returns Integer;
    ---C++: inline 
    ---C++: return const &

    LSC(me;  Index:  Integer) returns LinearScalarConstraint;
    --	"C   style" Index  :  Index  :  0 -->  nb_PPC-1
    ---C++: inline 
    ---C++: return const &


fields

    pnt2d : XY ;
    nb_PPConstraints : Integer;
    nb_LSConstraints : Integer;
    myPPC : PinpointConstraint[5]; 
    myLSC : LinearScalarConstraint[4];
    
end;

