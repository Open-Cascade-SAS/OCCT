-- Created on: 1997-11-06
-- Created by: Roman BORISOV
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

private  class PrjResolve from ProjLib 

	---Purpose: 

uses     
    Pnt2d     from gp,
    Surface from Adaptor3d, 
    Curve  from  Adaptor3d, 
    SurfacePtr from Adaptor3d, 
    CurvePtr  from Adaptor3d

raises   
    	DomainError from Standard, 
	ConstructionError,
    	NotDone     from StdFail

is
    Create (C: Curve  from  Adaptor3d; S: Surface from Adaptor3d;  Fix: Integer)
    	returns PrjResolve 
    	raises  ConstructionError;
    	
     
    Perform(me:  in  out;  t,  U,  V:  Real;  Tol,  Inf,  Sup:  Pnt2d;  FTol:  Real  from  Standard  =  -1;  StrictInside:  Boolean  from  Standard  =  Standard_False) 
---Purpose: Calculates the ort from  C(t)  to  S  with a close point.
    	--          The close point is defined by the parameter values
    	--          U0 and V0.
    	--          The function F(u,v)=distance(S(u,v),C(t)) has an
    	--          extremum when gradient(F)=0. The algorithm searchs
    	--          a zero near the close point.
    	raises  DomainError;
	    	-- if U0,V0 are outside the definition ranges of the 
	    	-- surface.
     
    
    IsDone (me)  returns Boolean
    	---Purpose: Returns True if the distance is found.
    	is static;
 
    Solution (me) returns Pnt2d  from  gp
    	---Purpose: Returns the point of the extremum distance.
    	raises  NotDone from StdFail
	    	-- if IsDone(me)=False.
    	is static;

fields
     
    myCurve    :  CurvePtr    from  Adaptor3d; 
    mySurface  :  SurfacePtr  from  Adaptor3d;	     
    myDone     :  Boolean     from  Standard;
    mySolution :  Pnt2d       from  gp; 
    myFix      :  Integer     from  Standard; 
     
end PrjResolve;
