-- Created on: 2021-03-15
-- Created by: Stephan GARNAUD (ARM)
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SharedMemory from OSD 

   ---Purpose: IPC Tools -Shared Memory
   --          This is a low level interface for communications.
   --          Using shared memory, processes can use a common area to
   --          communicate.
   --          You can create and delete a shared memory.

uses Error, AsciiString from TCollection
raises ConstructionError, NullObject, OSDError, ProgramError
   

is
  Create returns SharedMemory;
    ---Purpose: Allocates room for shared memory name.
    --          This is to be used with 'Open'.
    --          In this case, the process is a client of shared memory.
    ---Level: Advanced

  Create (Name : AsciiString ; size : Integer) returns SharedMemory
    ---Purpose: Instantiates SharedMemory object with parameters.
    --          A name to make sure shared memory is unique and a size in
    --          bytes for the size of shared memory.
    --
    --          Raises ConstructionError when the name contains characters 
    --          not in range of ' '...'~'.
    --          Raises ProgramError when the size given is negative or null.
    --          This is for a server process.
    --          
    ---Level: Advanced
    raises ConstructionError, ProgramError;

  Build (me : in out)  is static;
    ---Purpose: Creates a shared memory in the system
    --          This is for a server process.
    ---Level: Advanced

  Open (me : in out ; Name : AsciiString ; size : Integer)
    ---Purpose: Opens a shared memory
    --          Raises ConstructionError when the name contains characters 
    --          not in range of ' '...'~'.
    --          Raises ProgramError when the size given is negative or null.
    --          This is for a server process.
    --          
    ---Level: Advanced
    raises ConstructionError, ProgramError is static;

  Delete (me : in out)
    ---Purpose: Removes a shared memory access.
    --          This is used only by a server process !
    ---Level: Advanced
    raises ProgramError is static;

  GiveAddress (me) returns Address
    ---Purpose: Returns address of shared memory.
    --          Raises NullObject when the Shared Memory is not created.
    ---Level: Advanced
    raises NullObject is static;

  Failed (me) returns Boolean is static;
    ---Purpose: Returns TRUE if an error occurs
    ---Level: Advanced

  Reset (me : in out) is static;
    ---Purpose: Resets error counter to zero
    ---Level: Advanced
      
  Perror (me : in out)
    ---Purpose: Raises OSD_Error
    ---Level: Advanced
    raises OSDError is static;

 Error (me) returns Integer is static;
   ---Purpose: Returns error number if 'Failed' is TRUE.
    ---Level: Advanced

fields
   myId : Integer;     -- Shared memory ID
   myAddress    : Address;
   myName : AsciiString;   
   mySize : Integer;
   myError : Error;
end SharedMemory from OSD;

