-- File:	GeomToStep_MakeBSplineSurfaceWithKnots.cdl
-- Created:	Thu Aug  5 16:48:07 1993
-- Author:	Martine LANGLOIS
--		<mla@mastox>
---Copyright:	 Matra Datavision 1993

class MakeBSplineSurfaceWithKnots from GeomToStep  
    inherits Root from GeomToStep
    
    ---Purpose: This class implements the mapping between class
    --          BSplineSurface from Geom and the class
    --          BSplineSurfaceWithKnots from  
    --          StepGeom which describes a 
    --          bspline_Surface_with_knots from Prostep
  
uses BSplineSurface from Geom,
     BSplineSurfaceWithKnots from StepGeom
     
raises NotDone from StdFail
     
is 

Create ( Bsplin : BSplineSurface from Geom ) returns
    MakeBSplineSurfaceWithKnots;

Value (me) returns
    BSplineSurfaceWithKnots from StepGeom
    raises NotDone
    is static;
    ---C++: return const&

fields

    theBSplineSurfaceWithKnots :
    	BSplineSurfaceWithKnots from StepGeom;
    	-- The solution from StepGeom
    	
end MakeBSplineSurfaceWithKnots;


