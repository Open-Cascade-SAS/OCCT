-- Created on: 1992-03-27
-- Created by: Remi GILET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package GC

uses gp,
     gce,
     Geom,
     StdFail


    ---Level : Public. 
    --  All methods of all  classes will be public.


is

private deferred class Root;

---------------------------------------------------------------------------
--         Constructions of 3d geometrical elements from Geom.
---------------------------------------------------------------------------

class MakeLine;
    	---Purpose: Makes a Line from Geom.

class MakeCircle;
    	---Purpose: Makes a Circle from Geom.

class MakeHyperbola;
    	---Purpose: Makes an hyperbola from Geom.

class MakeEllipse;
    	---Purpose: Makes an ellipse from Geom.

class MakeSegment;
    	---Purpose: Makes a segment of Line from the 2 points <P1> and <P2>.

class MakeArcOfCircle;
    	---Purpose: Makes an arc of circle (TrimmedCurve from Geom).

class MakeArcOfEllipse;
    	---Purpose: Makes an arc of Ellipse (TrimmedCurve from Geom).

class MakeArcOfHyperbola;
    	---Purpose: Makes an arc of hyperbola (TrimmedCurve from Geom). 

class MakeArcOfParabola;
    	---Purpose: Makes an arc of parabola (TrimmedCurve from Geom).

---------------------------------------------------------------------------
--                   Constructions of planes from Geom.
---------------------------------------------------------------------------

class MakePlane;

---------------------------------------------------------------------------
--                  Construction of surfaces from Geom.
---------------------------------------------------------------------------

class MakeCylindricalSurface;
    ---Purpose: Makes a cylindricalSurface <Cyl> from Geom. 

class MakeConicalSurface;
    ---Purpose: Makes a ConicalSurface <Cone> from Geom.

class MakeTrimmedCylinder;
    ---Purpose: Makes a cylindricalSurface <Cyl> from Geom

class MakeTrimmedCone;
    ---Purpose: Makes a ConicalSurface <Cyl> from Geom

---------------------------------------------------------------------------
--               Constructions of Transformation from Geom.
---------------------------------------------------------------------------

class MakeTranslation;
    	---Purpose: Returns a translation transformation of vector <V>.

class MakeMirror;
    	---Purpose: Returns a symmetry transformation of center <P>.

class MakeRotation;
    	---Purpose: Returns a rotation transformation around the axis <A> 
    	--          and of angle <Angle>.

class MakeScale;
    	---Purpose: Returns a scaling transformation with the center point
    	--          <Point> and the scaling value <Scale>.

end GC;
