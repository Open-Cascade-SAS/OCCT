-- Created on: 1995-09-21
-- Created by: Philippe GIRODENGO
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class MeshExplorer from StlMesh 

	---Purpose: Provides  facilities to explore  the triangles  of
	--          each mesh domain.
	--          
uses  

    Mesh                   from StlMesh,
    SequenceOfMeshTriangle from StlMesh,
    SequenceOfXYZ          from TColgp

raises 

    OutOfRange   from Standard,
    NoMoreObject from Standard,
    NoSuchObject from Standard

is

    Create (M : Mesh)  returns MeshExplorer;
    

    Deflection (me) returns Real is static;
    	---Purpose: Returns the mesh deflection of the current domain.

    InitTriangle (me : in out; DomainIndex : Integer = 1)
    	---Purpose: Initializes the exploration  of the  triangles  of
    	--          the mesh domain of range <DomainIndex>.
    raises OutOfRange
    	---Purpose: Raised if <DomainIndex> is lower than 1 or greater
    	--          than the number of domains.
    is static;


    MoreTriangle (me) returns Boolean is static;
    	---C++: inline


    NextTriangle (me : in out) 
    raises NoMoreObject
    	---Purpose: Raised if there is no more triangle in the current
    	--          domain.
    is static;


    TriangleVertices (me; X1, Y1, Z1, X2, Y2, Z2, X3, Y3, Z3 : in out Real)
    raises NoSuchObject
    	---Purpose: Raised if there is no more triangle in the current
    	--          domain.
    is static;

   
    TriangleOrientation (me; Xn, Yn, Zn : in out Real)
    raises NoSuchObject
    	---Purpose: Raised if there is no more triangle in the current
    	--          domain.
    is static;



fields

    mesh            : Mesh;
    xn, yn, zn      : Real;
    v1, v2, v3      : Integer;
    domainIndex     : Integer;
    nbTriangles     : Integer;
    triangleIndex   : Integer;
    trianglesVertex : SequenceOfXYZ;
    trianglesdef    : SequenceOfMeshTriangle;

end MeshExplorer;







