-- Created on: 1993-06-03
-- Created by: fid
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package PColPGeom 

        ---Purpose : This package  is used to  instantiate of  several
        --         generic classes from  the package  PCollection with
        --         objects from the package PGeom.

uses PCollection, PGeom

is


    class HArray1OfCurve 
    	instantiates HArray1 from PCollection (Curve from PGeom);
    class HArray1OfBoundedCurve 
    	instantiates HArray1 from PCollection (BoundedCurve from PGeom);
    class HArray1OfBezierCurve 
    	instantiates HArray1 from PCollection (BezierCurve from PGeom);
    class HArray1OfBSplineCurve 
    	instantiates HArray1 from PCollection (BSplineCurve from PGeom);
    class HArray1OfSurface 
    	instantiates HArray1 from PCollection (Surface from PGeom);
    class HArray1OfBoundedSurface 
    	instantiates HArray1 from PCollection (BoundedSurface from PGeom);



    class HArray2OfSurface 
    	instantiates HArray2 from PCollection (Surface from PGeom);
    class HArray2OfBoundedSurface 
    	instantiates HArray2 from PCollection (BoundedSurface from PGeom);
    class HArray2OfBezierSurface 
    	instantiates HArray2 from PCollection (BezierSurface from PGeom);
    class HArray2OfBSplineSurface 
    	instantiates HArray2 from PCollection (BSplineSurface from PGeom);



--    class HSequenceOfCurve  
--    	instantiates HSequence from PCollection (Curve from PGeom);
--    class HSequenceOfBoundedCurve  
--    	instantiates HSequence from PCollection (BoundedCurve from PGeom);
--    class HSequenceOfSurface 
--    	instantiates HSequence from PCollection (Surface from PGeom);
--    class HSequenceOfBoundedSurface 
--    	instantiates HSequence from PCollection (BoundedSurface from PGeom);


end PColPGeom;
