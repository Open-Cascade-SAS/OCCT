-- File:	IGESDefs_ToolAssociativityDef.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolAssociativityDef  from IGESDefs

    ---Purpose : Tool to work on a AssociativityDef. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses AssociativityDef from IGESDefs,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolAssociativityDef;
    ---Purpose : Returns a ToolAssociativityDef, ready to work


    ReadOwnParams (me; ent : mutable AssociativityDef;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : AssociativityDef;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : AssociativityDef;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a AssociativityDef <ent>, from
    --           its specific (own) parameters

    DirChecker (me; ent : AssociativityDef) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : AssociativityDef;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : AssociativityDef; entto : mutable AssociativityDef;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : AssociativityDef;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolAssociativityDef;
