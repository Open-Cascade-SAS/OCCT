-- Created on: 2008-12-10
-- Created by: Pavel TELKOV
-- Copyright (c) 2008-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Datum from PXCAFDoc inherits  Attribute from PDF

	---Purpose: 
uses
    HAsciiString  from PCollection
is
    Create returns mutable Datum from PXCAFDoc;

    Create (theName : HAsciiString from PCollection;
    	    theDescr: HAsciiString from PCollection;
            theId   : HAsciiString from PCollection)
    returns mutable Datum from PXCAFDoc;
    
    GetName (me) returns HAsciiString from PCollection;

    GetDescription (me) returns HAsciiString from PCollection;

    GetIdentification (me) returns HAsciiString from PCollection;
    
    Set (me : mutable; theName : HAsciiString from PCollection;
    	    	       theDescr: HAsciiString from PCollection;
    	    	       theId   : HAsciiString from PCollection);
    
fields

    myName : HAsciiString from PCollection;
    myDescr: HAsciiString from PCollection;
    myId   : HAsciiString from PCollection;

end Datum from PXCAFDoc;
