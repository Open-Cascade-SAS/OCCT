-- File:	AIS_Circle.cdl
-- Created:	Tue Jan 21 11:45:01 1997
-- Author:	Prestataire Christiane ARMAND
--		<car@chamalox.paris1.matra-dtv.fr>
--   GG  :  GER61351 17/11/1999 Change SetColor() with a compatible Quantity_Color instead
--				       the restricted NameOfColor.
---Copyright:	 Matra Datavision 1997

class Circle from AIS inherits InteractiveObject from AIS

	---Purpose: Constructs circle datums to be used in construction of
    	-- composite shapes.

uses 
    Circle                from Geom,
    Point                 from Geom,
    Presentation          from Prs3d,
    PresentationManager3d from PrsMgr,
    NameOfColor           from Quantity,
    Color			  from Quantity,
    Selection             from SelectMgr,
    Projector             from Prs3d,
    Transformation        from Geom,
    PresentationManager2d from PrsMgr,
    GraphicObject         from Graphic2d,    
    Line                  from AIS,
    KindOfInteractive from AIS
    

is
    Create(aCircle : Circle from Geom) 
    returns mutable Circle from AIS;
    	---Purpose: Initializes this algorithm for constructing AIS circle
    	-- datums initializes the circle aCircle
    Create(aCircle : Circle from Geom;
    	   aUStart : Real from Standard;
    	   aUEnd   : Real from Standard;
	   aSens   : Boolean from Standard = Standard_True) 
    returns mutable Circle from AIS;
    	---Purpose: Initializes this algorithm for constructing AIS circle datums.    
    	-- Initializes the circle aCircle, the arc
    	--   starting point UStart, the arc ending point UEnd,
    	--   and the direction aSens.

    Compute(me            : mutable;
    	    aPresentationManager: PresentationManager3d from PrsMgr;
    	    aPresentation : mutable Presentation from Prs3d;
    	    aMode         : Integer from Standard = 0) 
    is redefined static  private;
    
    Compute(me:mutable;
    	        aProjector: Projector from Prs3d;
                aPresentation: mutable Presentation from Prs3d)
    is redefined static private;     

    Compute(me:mutable;
    	    aPresentationManager: PresentationManager2d from PrsMgr;
            aPresentation: mutable GraphicObject from Graphic2d;
            aMode: Integer from Standard = 0)
    is redefined static private;	

    Compute(me            : mutable;
            aProjector    : Projector from Prs3d;
            aTrsf         : Transformation from Geom;
            aPresentation : mutable Presentation from Prs3d)
    is redefined;
	 ---Purpose: computes the presentation according to a point of view
    	 --          given by <aProjector>.
	 --          To be Used when the associated degenerated Presentations
	 --          have been transformed by <aTrsf> which is not a Pure
	 --          Translation. The HLR Prs can't be deducted automatically
	 --          WARNING :<aTrsf> must be applied
	 --           to the object to display before computation  !!!

-- Methods from SelectableObject

    ComputeSelection(me         : mutable;
    	    	     aSelection : mutable Selection from SelectMgr;
    	    	     aMode      : Integer from Standard)is private;

 
-- Methods from InteractiveObject

  
  Signature(me) returns Integer from Standard is redefined;
	 ---C++: inline
	 ---Purpose: Returns index 6 by default.
  
  Type(me) returns KindOfInteractive from AIS is redefined;
	 ---C++: inline
	 ---Purpose: Indicates that the type of Interactive Object is a datum.
  
  Circle(me) returns any Circle from Geom;
	 ---C++: inline
	 ---C++: return const & 
	 ---Purpose: Returns the circle component defined in SetCircle.
   
  Parameters(me; u1,u2 : in out Real from Standard);
	 ---C++: inline
	 ---Purpose:
	 -- Constructs instances of the starting point and the end
	 -- point parameters, u1 and u2.
 
  SetCircle(me:mutable;aCircle : Circle from Geom);
 	 ---C++: inline
	 ---Purpose: Allows you to provide settings for the circle datum aCircle.
  
  SetFirstParam(me:mutable;u:Real);
	 ---C++: inline
	 ---Purpose: Allows you to set the parameter u for the starting point of an arc.
  
  SetLastParam(me:mutable;u:Real);
	 ---C++: inline
	 ---Purpose: Allows you to provide the parameter u for the end point of an arc.

    SetColor(me :mutable; aColor : NameOfColor from Quantity)
    is redefined static;
    	--- Purpose: Assigns the color aColor to the solid line boundary of the circle datum.
    SetColor(me :mutable; aColor : Color from Quantity)
    is redefined static;
         
    SetWidth(me:mutable; aValue:Real from Standard)
    is redefined static; 
    	---Purpose: Assigns the width aValue to the solid line boundary of the circle datum.
    UnsetColor(me:mutable)
    is redefined static; 
    	---Purpose: Removes color from the solid line boundary of the circle datum.    
    UnsetWidth(me:mutable)    
    is redefined static; 
    	---Purpose: Removes width settings from the solid line boundary of the circle datum.


    ComputeCircle(me: mutable;
                  aPresentation : mutable Presentation from Prs3d)
    is private;
     
    ComputeArc(me: mutable;
               aPresentation : mutable Presentation from Prs3d)
    is private;

    ComputeCircleSelection(me: mutable;
                           aSelection : mutable Selection from SelectMgr)
    is private;
     
    ComputeArcSelection(me: mutable;
                        aSelection : mutable Selection from SelectMgr)
    is private;

fields

    myComponent   : Circle  from Geom;
    myUStart      : Real    from Standard;
    myUEnd        : Real    from Standard;
    myCircleIsArc : Boolean from Standard;
    mySens        : Boolean from Standard;
    
end Circle ;
