-- Created on: 2008-12-28
-- Created by: Roman Lygin
-- Copyright (c) 2008-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

--            roman.lygin@gmail.com

generic class CurveCache from Extrema
    (Curve as any; -- Adaptor3d_Curve or Adaptor2d_Curve2d
     Pnt as any;   -- gp_Pnt or gp_Pnt2d
     ArrayOfPnt as Transient from Standard) -- TColgp_HArray1OfPnt or TColgp_HArray1OfPnt2d
inherits Transient from Standard

    ---Purpose:

uses
    Array1OfReal  from TColStd,
    HArray1OfReal from TColStd

raises NotDone from StdFail

is

    Create returns mutable CurveCache from Extrema;

    Create (theC: Curve; theUFirst, theULast: Real; theNbSamples: Integer;
        theToCalculate: Boolean)returns mutable CurveCache from Extrema;

    Create (theC: Curve; theUFirst, theULast: Real;
    	    IntervalsCN: Array1OfReal from TColStd;
	    StartIndex, EndIndex: Integer;
	    Coeff: Real)
    returns mutable CurveCache from Extrema;

    SetCurve (me: mutable; theC: Curve; theNbSamples: Integer;
        theToCalculate: Boolean);
    ---Purpose: Sets the \a theRank-th curve (1 or 2) and its parameters.
    --          Caches sample points for further reuse in Perform().

    SetCurve (me: mutable; theC: Curve;
        theUFirst, theULast: Real; theNbSamples: Integer; theToCalculate: Boolean);
        ---Purpose:

    SetRange (me: mutable; Uinf, Usup: Real; theToCalculate: Boolean);
    ---Purpose:

    CalculatePoints (me: mutable);
    ---Purpose: Calculates points along the curve and stores
    --          them in internal array for further reuse in Perform().

    IsValid (me) returns Boolean;
    ---C++: inline
    ---Purpose: Returns True if the points array has already been calculated
    --          for specified curve and range

    Parameters (me) returns HArray1OfReal from TColStd
        raises  NotDone from StdFail;
    ---C++: inline
    ---C++: return const &
    ---Purpose: Raises StdFail_NotDone if points have not yet been calculated.

    Points (me) returns ArrayOfPnt
        raises  NotDone from StdFail;
    ---C++: inline
    ---C++: return const &
    ---Purpose: Raises StdFail_NotDone if points have not yet been calculated.

    CurvePtr (me) returns Address from Standard;
    ---C++: inline
    ---Purpose:

    NbSamples (me) returns Integer;
    ---C++: inline
    ---Purpose:

    FirstParameter (me) returns Real;
    ---C++: inline
    ---Purpose:

    LastParameter (me) returns Real;
    ---C++: inline
    ---Purpose:

    TrimFirstParameter (me) returns Real;
    ---C++: inline
    ---Purpose: For bounded curves returns FirstParameter(), for unbounded - -1e-10.

    TrimLastParameter (me) returns Real;
    ---C++: inline
    ---Purpose: For bounded curves returns LastParameter(), for unbounded - 1e-10.

fields

    myC           : Address from Standard;
    myFirst       : Real;
    myLast        : Real;
    myTrimFirst   : Real;
    myTrimLast    : Real;
    myNbSamples   : Integer;
    myParamArray  : HArray1OfReal from TColStd;
    myPntArray    : ArrayOfPnt;
    myIsArrayValid: Boolean;

end;
