-- File:	ProjLib_ProjectedCurve.cdl
-- Created:	Wed Aug 25 15:07:07 1993
-- Author:	Bruno DUMORTIER
--		<dub@topsn3>
---Copyright:	 Matra Datavision 1993


class ProjectedCurve from ProjLib inherits Curve2d from Adaptor2d 
    


uses

     Projector       from ProjLib,
     Shape           from GeomAbs,
     CurveType       from GeomAbs,
     Vec2d           from gp,
     Pnt2d           from gp,
     Circ2d          from gp,
     Elips2d         from gp,
     Hypr2d          from gp,
     Parab2d         from gp,
     Lin2d           from gp,
     HCurve          from Adaptor3d,
     HCurve2d        from Adaptor2d,
     HSurface        from Adaptor3d,
     BezierCurve     from Geom2d,
     BSplineCurve    from Geom2d,
     Array1OfReal    from TColStd
     
     
raises
    
    OutOfRange          from Standard,
    NoSuchObject        from Standard,
    DomainError         from Standard,
    NotImplemented      from Standard
    
 
is

    Create returns ProjectedCurve;
    
    Create(S : HSurface from Adaptor3d) 
    returns ProjectedCurve;
    
    Create(S : HSurface from Adaptor3d; 
    	   C : HCurve   from Adaptor3d) 
    returns ProjectedCurve; 
      
    Create(S   : HSurface from Adaptor3d; 
    	   C   : HCurve   from Adaptor3d;
    	   Tol : Real     from Standard) 
    returns ProjectedCurve; 
      
    
    Load(me : in out ; Tolerance : Real) 
    ---Purpose: Changes the tolerance used to project
    --          the curve on the surface
    is static;
    
    Load(me : in out; S : HSurface from Adaptor3d)
	---Purpose: Changes the Surface.
    is static;
    
    Load(me : in out; C : HCurve from Adaptor3d)
	---Purpose: Changes the Curve.
    is static;
    
    GetSurface(me) returns HSurface from Adaptor3d
	---C++: return const &
    is static;

    GetCurve(me) returns  HCurve from Adaptor3d 
	---C++: return const &
    is static;
    
    GetTolerance(me) returns Real from Standard
	---Purpose: returns the tolerance reached if an approximation
	--          is Done.
    is static;

    --
    --     Global methods - Apply to the whole curve.
    --     
    
    FirstParameter(me) returns Real
    is redefined static;

    LastParameter(me) returns Real
    is redefined static;
    
    Continuity(me) returns Shape from GeomAbs
    is redefined static;
    
    NbIntervals(me ; S : Shape from GeomAbs) returns Integer
	---Purpose: If necessary,  breaks the  curve in  intervals  of
	--          continuity  <S>.    And  returns   the number   of
	--          intervals.
    is redefined static;
    
    Intervals(me; T : in out Array1OfReal from TColStd; 
    	          S : Shape from GeomAbs)
	---Purpose: Stores in <T> the  parameters bounding the intervals
	--          of continuity <S>.
	--          
	--          The array must provide  enough room to  accomodate
	--          for the parameters. i.e. T.Length() > NbIntervals()
    raises
    	OutOfRange from Standard 
    is redefined static;
    
    Trim(me; First, Last, Tol : Real) returns HCurve2d from Adaptor2d
	---Purpose: Returns    a  curve equivalent   of  <me>  between
	--          parameters <First>  and <Last>. <Tol>  is used  to
	--          test for 3d points confusion.
    raises
    	OutOfRange from Standard
	---Purpose: If <First> >= <Last> 
    is redefined static;
    
    IsClosed(me) returns Boolean
    is redefined static;
     
    IsPeriodic(me) returns Boolean
    is redefined static;
    
    Period(me) returns Real
    raises
    	DomainError from Standard -- if the curve is not periodic
    is redefined static;
     
    Value(me; U : Real) returns Pnt2d from gp
         --- Purpose : Computes the point of parameter U on the curve.
    is redefined static;
    
    D0 (me; U : Real; P : out Pnt2d from gp)
         --- Purpose : Computes the point of parameter U on the curve.
    is redefined static;
    
    D1 (me; U : Real; P : out Pnt2d from gp ; V : out Vec2d from gp)
         --- Purpose : Computes the point of parameter U on the curve with its
         --  first derivative.
     raises 
    	DomainError from Standard
        --- Purpose : Raised if the continuity of the current interval
        --  is not C1.
    is redefined static;
    
    D2 (me; U : Real; P : out Pnt2d from gp; V1, V2 : out Vec2d from gp)
        --- Purpose :
        --  Returns the point P of parameter U, the first and second
        --  derivatives V1 and V2.
     raises 
    	DomainError from Standard
        --- Purpose : Raised if the continuity of the current interval
        --  is not C2.
     is redefined static;

    D3 (me; U : Real; P : out Pnt2d from gp; V1, V2, V3 : out Vec2d from gp)
        --- Purpose :
        --  Returns the point P of parameter U, the first, the second 
        --  and the third derivative.
     raises 
    	DomainError from Standard
        --- Purpose : Raised if the continuity of the current interval
        --  is not C3.
     is redefined static;
        
    DN (me; U : Real; N : Integer)   returns Vec2d from gp
        --- Purpose :
        --  The returned vector gives the value of the derivative for the 
        --  order of derivation N.
     raises  
    	DomainError from Standard,
        --- Purpose : Raised if the continuity of the current interval
        --  is not CN.
        OutOfRange from Standard
        --- Purpose : Raised if N < 1.            
     is redefined static;

    Resolution(me; R3d : Real) returns Real
         ---Purpose :  Returns the parametric  resolution corresponding
         --         to the real space resolution <R3d>.
    is redefined static;   
        
    GetType(me) returns CurveType from GeomAbs
	---Purpose: Returns  the  type of the   curve  in the  current
	--          interval :   Line,   Circle,   Ellipse, Hyperbola,
	--          Parabola, BezierCurve, BSplineCurve, OtherCurve.
    is redefined static;

    --
    --     The following methods must  be called when GetType returned
    --     the corresponding type.
    --     

     Line(me) returns Lin2d from gp
     raises 
    	NoSuchObject from Standard
     is redefined static;
     
     Circle(me) returns Circ2d from gp
     raises 
    	NoSuchObject from Standard
     is redefined static;
     
     Ellipse(me) returns Elips2d from gp
     raises 
    	NoSuchObject from Standard
     is redefined static;
     
     Hyperbola(me) returns  Hypr2d from gp
     raises 
    	NoSuchObject from Standard
     is redefined static;
     
     Parabola(me) returns Parab2d from gp
     raises 
    	NoSuchObject from Standard
     is redefined static;
     
     Degree(me) returns Integer
     raises 
    	NoSuchObject from Standard
     is redefined static;
     
     IsRational(me) returns Boolean
     raises 
    	NoSuchObject from Standard
     is redefined static;
     
     NbPoles(me) returns Integer
     raises 
    	NoSuchObject from Standard
     is redefined static;
     
    
     NbKnots(me) returns Integer
     raises 
    	NoSuchObject from Standard
     is redefined static;
     
     


     Bezier(me) returns BezierCurve from Geom2d
     raises 
    	NoSuchObject from Standard
     is redefined static;
     ---Purpose:  Warning ! This will  NOT make a copy  of the -- Bezier Curve -
     --         If you want to modify -- the Curve  please make a copy
     --         yourself --  Also it will  NOT trim the surface  to --
     --         myFirst/Last.
    
     BSpline(me) returns BSplineCurve from Geom2d
     raises 
    	NoSuchObject from Standard
     is redefined static;
      ---Purpose:  Warning ! This will NOT make a copy of the BSpline Curve - If
      --         you want to  modify the   Curve  please make a   copy
      --         yourself Also it   will  NOT  trim   the surface   to
      --         myFirst/Last.
     
    
fields

     myTolerance : Real ;
     mySurface   : HSurface   from Adaptor3d ;
     myCurve     : HCurve     from Adaptor3d ;
     myResult    : Projector  from ProjLib ;
     
end ProjectedCurve;
