-- Created on: 2000-11-21
-- Created by: Peter KURNEV
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class VEInterference from BOPTools 
    inherits ShapeShapeInterference from BOPTools  
     
    	---Purpose:  
    	--  class for storing info about an Verex/Edge interference
	--- 

is 
    Create  
    	returns  VEInterference from BOPTools; 
    	---Purpose: 
    	--- Empty constructor  
    	---
    Create  (anIndex1, anIndex2:  Integer from Standard; 
    	    aT: Real from Standard)
    	returns  VEInterference from BOPTools;  
    	---Purpose:   
    	--- Constructor  
    	--- anIndex1,  
    	--- anIndex2 see BOPTools_ShapeShapeInterference for details      
    	--- aT -  values of parameter on the edge    
    	---
    SetParameter  (me:out; aT: Real from Standard); 
    	---Purpose:  
    	--- Modifier   
    	---
    Parameter     (me) 
	returns Real from Standard;   
    	---Purpose:  
    	--- Selector  
    	---
    
fields
    myParameter:  Real from Standard;  

end VEInterference;
