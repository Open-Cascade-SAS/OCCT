-- File:	StepElement_UniformSurfaceSection.cdl
-- Created:	Thu Dec 12 17:29:05 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class UniformSurfaceSection from StepElement
inherits SurfaceSection from StepElement

    ---Purpose: Representation of STEP entity UniformSurfaceSection

uses
    MeasureOrUnspecifiedValue from StepElement

is
    Create returns UniformSurfaceSection from StepElement;
	---Purpose: Empty constructor

    Init (me: mutable; aSurfaceSection_Offset: MeasureOrUnspecifiedValue from StepElement;
                       aSurfaceSection_NonStructuralMass: MeasureOrUnspecifiedValue from StepElement;
                       aSurfaceSection_NonStructuralMassOffset: MeasureOrUnspecifiedValue from StepElement;
                       aThickness: Real;
                       aBendingThickness: MeasureOrUnspecifiedValue from StepElement;
                       aShearThickness: MeasureOrUnspecifiedValue from StepElement);
	---Purpose: Initialize all fields (own and inherited)

    Thickness (me) returns Real;
	---Purpose: Returns field Thickness
    SetThickness (me: mutable; Thickness: Real);
	---Purpose: Set field Thickness

    BendingThickness (me) returns MeasureOrUnspecifiedValue from StepElement;
	---Purpose: Returns field BendingThickness
    SetBendingThickness (me: mutable; BendingThickness: MeasureOrUnspecifiedValue from StepElement);
	---Purpose: Set field BendingThickness

    ShearThickness (me) returns MeasureOrUnspecifiedValue from StepElement;
	---Purpose: Returns field ShearThickness
    SetShearThickness (me: mutable; ShearThickness: MeasureOrUnspecifiedValue from StepElement);
	---Purpose: Set field ShearThickness

fields
    theThickness: Real;
    theBendingThickness: MeasureOrUnspecifiedValue from StepElement;
    theShearThickness: MeasureOrUnspecifiedValue from StepElement;

end UniformSurfaceSection;
