-- Created on: 1993-06-14
-- Created by: Martine LANGLOIS
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MakeAxis2Placement3d from GeomToStep inherits Root from GeomToStep

    ---Purpose: This class implements the mapping between classes 
    --          Axis2Placement from Geom and Ax2, Ax3 from gp, and the class
    --          Axis2Placement3d from StepGeom which describes an
    --          axis2_placement_3d from Prostep. 
   
uses Ax2 from gp,
     Ax3 from gp,
     Trsf from gp,
     Axis2Placement from Geom,
     Axis2Placement3d from StepGeom
     
raises NotDone from StdFail
     
is 

Create returns MakeAxis2Placement3d;
-- creates an identity (original axis)

Create ( A : Ax2 from gp ) returns MakeAxis2Placement3d;

Create ( A : Ax3 from gp ) returns MakeAxis2Placement3d;

Create ( T : Trsf from gp) returns MakeAxis2Placement3d;

Create ( A : Axis2Placement from Geom ) returns MakeAxis2Placement3d;

Value (me) returns Axis2Placement3d from StepGeom
    raises NotDone
    is static;
    ---C++: return const&

fields

    theAxis2Placement3d : Axis2Placement3d from StepGeom;
    	-- TheOP solution from StepGeom
    	
end MakeAxis2Placement3d;


