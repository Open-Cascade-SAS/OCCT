-- Created on: 2001-07-25
-- Created by: Julia DOROVSKIKH
-- Copyright (c) 2001-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DocumentStorageDriver from XmlDrivers inherits DocumentStorageDriver from XmlLDrivers

uses
    ExtendedString              from TCollection,
    ADriverTable		from XmlMDF, 
    Element                     from XmlObjMgt,
    MessageDriver               from CDM

is
    Create (theCopyright: ExtendedString from TCollection)
    	returns DocumentStorageDriver from XmlDrivers;
    -- Constructor

    AttributeDrivers  (me : mutable; theMsgDriver: MessageDriver from CDM)
	returns ADriverTable from XmlMDF
	is redefined virtual;

    WriteShapeSection (me:mutable; thePDoc  : out Element from XmlObjMgt)  
        returns Boolean from Standard
        is redefined virtual; 
    
end DocumentStorageDriver;
