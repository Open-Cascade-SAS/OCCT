-- Created on: 1992-08-26
-- Created by: Jean Louis FRENKEL
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package Prs3d

      ---Purpose: The Prs3d package provides the following services
  -- -   a presentation object (the context for all
  --   modifications to the display, its presentation will be
  --   displayed in every view of an active viewer)
  -- -   an attribute manager governing how objects such
  --   as color, width, and type of line are displayed;
  --   these are generic objects, whereas those in
  --   StdPrs are specific geometries and topologies.
  -- -   generic   algorithms providing default settings for
  --   objects such as points, curves, surfaces and shapes
  -- -   a root object which provides the abstract
  --   framework for the DsgPrs definitions at work in
  --   display of dimensions, relations and trihedra.
    
uses
  Graphic3d,
  Aspect,
  Quantity,
  MMgt,
  Standard,
  Adaptor3d,
  BRepAdaptor,
  Geom,
  CPnts,
  GCPnts,
  TopAbs,
  TopLoc,
  TopoDS,
  TopTools,
  TopExp,
  HLRAlgo,
  TCollection,
  TColgp,
  Bnd,
  gp,
  Poly,
  TColStd
is  
  exception InvalidAngle inherits RangeError from Standard;

  enumeration TypeOfLinePicking is TOLP_Point,
                                   TOLP_Segment
  end TypeOfLinePicking;
        
  enumeration TypeOfHLR is TOH_NotSet,
                           TOH_PolyAlgo,
                           TOH_Algo;
  ---Purpose: Declares types of hidden line removal algorithm.
  --          TOH_Algo enables using of exact HLR algorithm.
  --          TOH_PolyAlgo enables using of polygonal HLR algorithm.
  --          TOH_NotSet is used by Prs3d_Drawer class, it means that the drawer should return the global value.
  --          For more details see Prs3d_Drawer class, AIS_Shape::Compute() method and
  --          HLRAlgo package from TKHLR toolkit.
  
  enumeration DimensionTextHorizontalPosition is DTHP_Left, DTHP_Right, DTHP_Center, DTHP_Fit;
  ---Purpose: Specifies options for positioning dimension value label in horizontal direction.
  -- DTHP_Left   - value label located at left side on dimension extension.
  -- DTHP_Right  - value label located at right side on dimension extension.
  -- DTHP_Center - value label located at center of dimension line.
  -- DTHP_Fit    - value label located automatically at left side if does not fits
  --               the dimension space, otherwise the value label is placed at center.

  enumeration DimensionTextVerticalPosition is DTVP_Above, DTVP_Below, DTVP_Center;
  ---Purpose: Specifies options for positioning dimension value label in vertical direction
  -- with respect to dimension (extension) line.
  -- DTVP_Above - text label is located above the dimension or extension line.
  -- DTVP_Below - text label is located below the dimension or extension line.
  -- DTVP_Center - the text label middle-point is in line with dimension or extension line.

  enumeration DimensionArrowOrientation is DAO_Internal, DAO_External, DAO_Fit;
  ---Purpose: Specifies dimension arrow location and orientation.
  -- DAO_Internal - arrows "inside", pointing outwards.
  -- DAO_External - arrows "outside", pointing inwards.
  -- DAO_Fit      - arrows oriented inside if value label with arrowtips fit the dimension line,
  --                otherwise - externally

  enumeration VertexDrawMode is VDM_Isolated, VDM_All, VDM_Inherited;
  ---Purpose: Describes supported modes of visualization of the shape's vertices:
  -- VDM_Isolated  - only isolated vertices (not belonging to a face) are displayed.
  -- VDM_All       - all vertices of the shape are displayed.
  -- VDM_Inherited - the global settings are inherited and applied to the shape's presentation.

  class Presentation;

  ---Category: Aspect classes.

  deferred class BasicAspect;	
  class PointAspect;
  class LineAspect;
  class ShadingAspect;
  class TextAspect;
  class IsoAspect;
  class ArrowAspect;
  class PlaneAspect;
  class DimensionAspect;
  class DatumAspect;
  imported DimensionUnits;

  imported transient class Drawer;

  class Projector;

  class PlaneSet;

  deferred class Root;

  ---Category: Basis construction elements.

  class Text;

        ---Category: Class signatures.

  class ShapeTool;

  class Arrow;
  ---Purpose: draws an arrow at a given location, with respect
  --          to a given direction.

  imported NListOfSequenceOfPnt; 
  imported NListIteratorListOfSequenceOfPnt;
  imported Point;
  imported WFShape;
  
  MatchSegment(X,Y,Z: Length from Quantity;
              aDistance: Length from Quantity;
              p1,p2: Pnt from gp;
              dist: out Length from Quantity)
  returns Boolean from Standard;

  GetDeflection (theShape  : Shape from TopoDS;
                 theDrawer : Drawer from Prs3d)
  returns Real from Standard;
  ---Purpose: Computes the absolute deflection value depending on
  -- the type of deflection in theDrawer:
  -- <ul>
  -- <li><b>Aspect_TOD_RELATIVE</b>: the absolute deflection is computed using the relative
  --   deviation coefficient from theDrawer and the shape's bounding box;</li>
  -- <li><b>Aspect_TOD_ABSOLUTE</b>: the maximal chordial deviation from theDrawer is returned.</li>
  -- </ul>
  -- This function should always be used to compute the deflection value for building
  -- discrete representations of the shape (triangualtion, wireframe) to avoid incosistencies
  -- between different representations of the shape and undesirable visual artifacts.
end Prs3d;
