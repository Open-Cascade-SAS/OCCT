-- Created on: 1995-03-13
-- Created by: Christian CAILLET
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package XSControl

    ---Purpose : This package provides complements to IFSelect & Co for
    --           control of a session

uses Standard , MMgt, TCollection , TColStd, Dico,
     Interface, Transfer, IFSelect, Message, MoniTool,
     TopoDS,    TopTools, TopAbs ,   Geom, Geom2d, gp

is

    deferred class Controller;
    class TransferReader;
    class TransferWriter;

    class WorkSession;
    class SelectForTransfer;
    class SignTransferStatus;
    class ConnectedShapes;

    class Reader;
    class Writer;

    class Functions;
    class FuncShape;
    class Utils;
    class Vars;

    Session (pilot : SessionPilot from IFSelect) returns WorkSession from XSControl;
    ---Purpose : Returns the WorkSession of a SessionPilot, but casts it as
    --           from XSControl : it then gives access to Control & Transfers

    Vars    (pilot : SessionPilot from IFSelect) returns Vars from XSControl;
    ---Purpose : Returns the Vars of a SessionPilot, it is brought by Session
    --           it provides access to external variables

end XSControl;
