-- Created on: 1998-11-25
-- Created by: Julia GERASIMOVA
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Aij from GeomPlate

	---Purpose: A structure containing indexes of two normals and its cross product

uses
    Vec from gp
is
    Create returns Aij from GeomPlate;
    
    Create( anInd1 : Integer from Standard;
    	    anInd2 : Integer from Standard;
	    aVec   : Vec from gp )
    returns Aij from GeomPlate;

fields

    Ind1 : Integer from Standard;
    Ind2 : Integer from Standard;
    Vec  : Vec from gp;

friends
    class BuildAveragePlane from GeomPlate

end Aij;
