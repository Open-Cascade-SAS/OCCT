-- File:	RWStepBasic_RWAction.cdl
-- Created:	Fri Nov 26 16:26:28 1999 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0
-- Copyright:	Matra Datavision 1999

class RWAction from RWStepBasic

    ---Purpose: Read & Write tool for Action

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    Action from StepBasic

is
    Create returns RWAction from RWStepBasic;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : Action from StepBasic);
	---Purpose: Reads Action

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: Action from StepBasic);
	---Purpose: Writes Action

    Share (me; ent : Action from StepBasic;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWAction;
