-- Created on: 1993-07-06
-- Created by: Yves FRICAUD
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package MAT2d 

	---Purpose : Package of computation of Bisector locus on a
        --           Set of geometrys from Geom2d.

uses
    GeomAbs,
    MMgt,
    gp,
    Geom2d,
    TColStd,
    TCollection,
    TColgp,
    TColGeom2d,
    MAT,
    Bisector

is

    deferred class SketchExplorer;

    class Tool2d;

    class Mat2d;

    class Connexion;

    class MiniPath;

    class Circuit;

    class CutCurve;   

    class SequenceOfConnexion instantiates Sequence  from TCollection
    	    	    	    	    	    	     (Connexion from  MAT2d); 

    class DataMapOfIntegerSequenceOfConnexion instantiates DataMap 
                   from TCollection (Integer              from Standard,
				     SequenceOfConnexion  from MAT2d,
				     MapIntegerHasher     from TColStd);
                                         
    class Array2OfConnexion  instantiates Array2 from TCollection
   	    	    	    	    	    	     (Connexion from  MAT2d); 
               

    class DataMapOfIntegerBisec  instantiates DataMap from TCollection 
    	                                   (Integer          from Standard,
					    Bisec            from Bisector,
					    MapIntegerHasher from TColStd); 
					    
    class DataMapOfIntegerPnt2d  instantiates DataMap from TCollection 
    	                                   (Integer          from Standard,
					    Pnt2d            from gp,
					    MapIntegerHasher from TColStd);  
	    
    class DataMapOfIntegerVec2d  instantiates DataMap from TCollection 
    	                                   (Integer          from Standard,
					    Vec2d            from gp,
					    MapIntegerHasher from TColStd); 

    class SequenceOfSequenceOfCurve  instantiates Sequence from TCollection 
    	                                    (SequenceOfCurve from TColGeom2d); 
					    
    class SequenceOfSequenceOfGeometry instantiates Sequence from TCollection
    	                                (SequenceOfGeometry from  TColGeom2d); 

    class DataMapOfIntegerConnexion instantiates DataMap from TCollection 
    	                                   (Integer          from Standard,
					    Connexion        from MAT2d,
					    MapIntegerHasher from TColStd);

    class BiInt;
	
    class MapBiIntHasher;
    
    class DataMapOfBiIntSequenceOfInteger instantiates DataMap 
         from TCollection (BiInt               from MAT2d,
			   SequenceOfInteger   from TColStd,
			   MapBiIntHasher      from MAT2d);
        
    class DataMapOfBiIntInteger instantiates DataMap 
         from TCollection (BiInt               from MAT2d,
			   Integer             from Standard,
			   MapBiIntHasher      from MAT2d);
end MAT2d;



