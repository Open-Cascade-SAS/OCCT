-- Created on: 2002-02-01
-- Created by: QA Admin
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package QADraw
    uses Draw
is
    
    CommonCommands(DI : in out Interpretor from Draw);
    ---Purpose: Define specicial commands for AIS.

    AdditionalCommands(DI : in out Interpretor from Draw);
    
    Factory (DI : out Interpretor from Draw);
    ---Purpose: Loads all QA Draw commands. Used for plugin.

end;
    
