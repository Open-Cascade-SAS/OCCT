-- Created on: 2007-08-17
-- Created by: Sergey ZARITCHNY
-- Copyright (c) 2007-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class HDataMapOfStringInteger from TDataStd inherits TShared from MMgt 

	---Purpose: Extension of TColStd_DataMapOfStringInteger class  
    	--    	    to be manipulated by handle. 

uses
    DataMapOfStringInteger from TColStd 
    
is
    Create( NbBuckets: Integer from Standard = 1 )  
    returns mutable HDataMapOfStringInteger from TDataStd;    
     
    Create( theOther:  DataMapOfStringInteger from TColStd)  
    returns mutable HDataMapOfStringInteger from TDataStd;
     
    Map( me ) returns DataMapOfStringInteger from TColStd
	---C++: return const &
        ---C++: inline      
    is static;	    	
	  
    ChangeMap( me: mutable ) returns DataMapOfStringInteger from TColStd 
    	---C++: return &
        ---C++: inline 
    is static; 	    	
 
fields
    
    myMap : DataMapOfStringInteger from TColStd ;  
   
end HDataMapOfStringInteger;
