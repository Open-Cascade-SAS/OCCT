-- Created on: 1994-04-05
-- Created by: Yves FRICAUD
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



private class FunctionH from Bisector 

inherits FunctionWithDerivative from math
     
             --                                  2           2 
	---Purpose: H(v) = (T1  .P2(v) - P1) * ||T(v)||  -
	--                                  2         2
	--                 (T(v).P2(v) - P1) * ||T1|| 
	
uses 
    Curve from Geom2d,
    Pnt2d from gp, 
    Vec2d from gp  

is

    Create (C2 : Curve from Geom2d ;
            P1 : Pnt2d from gp     ;
            T1   : Vec2d from gp   ) 
    returns FunctionH from Bisector;
    
    Value(me : in out; X : Real; F : out Real) 
    	---Purpose: Computes the values of the Functions for the variable <X>.
    returns Boolean;
    
    Derivative(me : in out; X : Real; D : out Real) 
    returns Boolean;

    Values(me : in out ; X  : Real; F  : out Real; D  : out Real)    
    	---Purpose: Returns the values of the functions and the derivatives
    	--          for the variable <X>.
    returns Boolean;

fields
    
    curve2 : Curve from Geom2d;
    p1     : Pnt2d from gp;
    t1     : Vec2d from gp;
    
end FunctionH;
