-- Created on: 1993-01-09
-- Created by: CKY / Contract Toubro-Larsen ( Arun MENON )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class GroupWithoutBackP from IGESBasic  inherits Group

        ---Purpose: defines GroupWithoutBackP, Type <402> Form <7>
        --          in package IGESBasic
        --          this class defines a Group without back pointers
        --          
        --          It inherits from Group

uses

        Transient        ,
        HArray1OfIGESEntity from IGESData

raises OutOfRange

is

        Create returns mutable GroupWithoutBackP;

        -- Specific Methods pertaining to the class : see Group

--
-- Class    : IGESBasic_GroupWithoutBackP
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class GroupWithoutBackP.
--
-- Reminder : A GroupWithoutBackP instance is defined by :
--            - an array of Entities
--            See Group

end GroupWithoutBackP;
