-- Created on: 1998-03-23
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class C2DF from TopOpeBRepTool

uses

    Curve from Geom2d,
    Face from TopoDS

is

    Create returns C2DF from TopOpeBRepTool;    
    Create(PC : Curve from Geom2d; f2d,l2d,tol : Real; F : Face from TopoDS) 
    returns C2DF from TopOpeBRepTool;
    SetPC(me : in out;PC : Curve from Geom2d; f2d,l2d,tol : Real);
    SetFace(me : in out; F : Face from TopoDS);
    PC(me; f2d,l2d,tol : out Real) returns Curve from Geom2d;
    ---C++: return const &
    Face(me) returns Face from TopoDS;
    ---C++: return const &
    IsPC(me;PC:Curve from Geom2d) returns Boolean;
    IsFace(me;F:Face from TopoDS) returns Boolean;
    
fields
    
    myPC : Curve from Geom2d;
    myf2d,myl2d,mytol : Real;
    myFace : Face from TopoDS;
    
end C2DF;
