-- Created on: 1996-10-11
-- Created by: Philippe MANGIN
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

private class Newton from FairCurve inherits NewtonMinimum from  math

	---Purpose: Algorithme of Optimization used to make "FairCurve"

uses 
    Vector from math, 
    MultipleVarFunctionWithHessian from math

is
    Create(theFunction: in MultipleVarFunctionWithHessian;
    	   theSpatialTolerance:  Real = 1.0e-7;
           theCriteriumTolerance: Real=1.0e-7;
	   theNbIterations: Integer=40; 
           theConvexity: Real=1.0e-6; 
           theWithSingularity:  Boolean = Standard_True)
    ---Purpose:
    -- The tolerance  required on  the  solution is given  by Tolerance.  
    -- Iteration are  stopped if (!WithSingularity)  and H(F(Xi)) is not definite
    -- positive  (if the smaller eigenvalue of H < Convexity)
    -- or IsConverged() returns True for 2 successives Iterations.
    -- Warning: This constructor do not computation 
    returns  Newton;   
	   
    IsConverged(me)
    	---Purpose: 
        -- This method is  called    at the end  of   each
    	-- iteration to  check the convergence :
    	-- || Xi+1 - Xi || < SpatialTolerance/100 Or
    	-- || Xi+1 - Xi || < SpatialTolerance and
    	-- |F(Xi+1) - F(Xi)| < CriteriumTolerance * |F(xi)|
    	-- It can be redefined in a sub-class to implement a specific test.
   
    returns Boolean is redefined;    

fields
    mySpTol : Real;
end Newton;

