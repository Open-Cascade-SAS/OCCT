-- Created on: 1991-03-27
-- Created by: Michel CHAUVAT
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package LProp

    ---Purpose: Handles local properties of curves and surfaces.
    --          Given a curve and a parameter value the following computations
    --          are available :
    --          - point,
    --          - derivatives,
    --          - tangent,
    --          - normal,
    --          - curvature,
    --          - centre of curvature,
    --          - Locals curvature's extremas,
    --          - Points of inflection,
    --          Given a surface and 2 parameters the following computations
    --          are available :
    --          - for each parameter:
    --            - derivatives,
    --            - tangent line,
    --            - centre of curvature,
    --          - point,
    --          - normal line,
    --          - maximum and minimum curvatures,
    --          - principal directions of curvature,
    --          - mean curvature,
    --          - Gaussian curvature.


    ---Level : Public. 
    --  All methods of all  classes will be public.

uses Standard, gp, math, TCollection, TColStd, GeomAbs

is

    enumeration Status is Undecided , Undefined, Defined, Computed;
    enumeration CIType is Inflection, MinCur   , MaxCur;
    	---Purpose:
    	-- Identifies the type of a particular point on a curve:
    	-- - LProp_Inflection: a point of inflection
    	-- - LProp_MinCur: a minimum of curvature
    	-- - LProp_MaxCur: a maximum of curvature.
        
    exception BadContinuity inherits Failure;
    exception NotDefined    inherits Failure;
    
    generic class CLProps;

    generic class SLProps;

    class CurAndInf;	

    class AnalyticCurInf;

    private class SequenceOfCIType instantiates Sequence from TCollection 
						        (CIType  from  LProp); 
    
end LProp;    
