-- Created on: 1993-06-11
-- Created by: Martine LANGLOIS
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class MakeCartesianPoint from GeomToStep inherits Root from GeomToStep

    ---Purpose: This class implements the mapping between classes 
    --          CartesianPoint from Geom and Pnt from gp, and the class
    --          CartesianPoint from StepGeom which describes a point from
    --          Prostep. 
  
uses Pnt from gp,
     Pnt2d from gp,
     CartesianPoint from Geom,
     CartesianPoint from Geom2d,
     CartesianPoint from StepGeom
     
raises NotDone from StdFail
     
is 

Create ( P : Pnt from gp ) returns MakeCartesianPoint;

Create ( P : Pnt2d from gp ) returns MakeCartesianPoint;

Create ( P : CartesianPoint from Geom ) returns MakeCartesianPoint;

Create ( P : CartesianPoint from Geom2d ) returns MakeCartesianPoint;

Value (me) returns CartesianPoint from StepGeom
    raises NotDone
    is static;
    ---C++: return const&
    
fields

    theCartesianPoint : CartesianPoint from StepGeom;
    	-- The solution from StepGeom
    	
end MakeCartesianPoint;


