-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SurfaceStyleElementSelect from StepVisual inherits SelectType from StepData

	-- <SurfaceStyleElementSelect> is an EXPRESS Select Type construct translation.
	-- it gathers : SurfaceStyleFillArea, SurfaceStyleBoundary, SurfaceStyleSilhouette, SurfaceStyleSegmentationCurve, SurfaceStyleControlGrid, SurfaceStyleParameterLine
	-- Rev4 : only remain SurfaceStyleFillArea, SurfaceStyleBoundary, SurfaceStyleParameterLine

uses

	SurfaceStyleFillArea,
	SurfaceStyleBoundary,
--	SurfaceStyleSilhouette,
--	SurfaceStyleSegmentationCurve,
--	SurfaceStyleControlGrid,
	SurfaceStyleParameterLine
is

	Create returns SurfaceStyleElementSelect;
	---Purpose : Returns a SurfaceStyleElementSelect SelectType

	CaseNum (me; ent : Transient) returns Integer;
	---Purpose: Recognizes a SurfaceStyleElementSelect Kind Entity that is :
	--        1 -> SurfaceStyleFillArea
	--        2 -> SurfaceStyleBoundary
	--        3 -> SurfaceStyleParameterLine
	--        4 -> SurfaceStyleSilhouette
	--        5 -> SurfaceStyleSegmentationCurve
	--        6 -> SurfaceStyleControlGrid
	--        0 else

	SurfaceStyleFillArea (me) returns any SurfaceStyleFillArea;
	---Purpose : returns Value as a SurfaceStyleFillArea (Null if another type)

	SurfaceStyleBoundary (me) returns any SurfaceStyleBoundary;
	---Purpose : returns Value as a SurfaceStyleBoundary (Null if another type)

	SurfaceStyleParameterLine (me) returns any SurfaceStyleParameterLine;
	---Purpose : returns Value as a SurfaceStyleParameterLine (Null if another type)


end SurfaceStyleElementSelect;

