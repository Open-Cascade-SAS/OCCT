-- Created on: 1991-12-13
-- Created by: Christophe MARION
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Intervals from Intrv
	---Purpose: The class  Intervals is a  sorted  sequence of non
	--          overlapping  Real Intervals.

uses
    Integer            from Standard,
    Interval           from Intrv,
    SequenceOfInterval from Intrv

raises
    OutOfRange

is
    Create returns Intervals from Intrv;
	---Purpose: Creates a void sequence of intervals.

    Create(Int : Interval from Intrv) returns Intervals from Intrv;
	---Purpose: Creates a sequence of one interval.
	
    Create(Int : Intervals from Intrv) returns Intervals from Intrv;
	---Purpose: Creates   by   copying  an   existing  sequence of
	--          intervals.
	
    Intersect(me : in out; Tool : Interval from Intrv)
	---Purpose: Intersects the intervals with the interval <Tool>.
    is static;

    Intersect(me : in out; Tool : Intervals from Intrv)
	---Purpose: Intersects the intervals with the intervals in the
	--          sequence  <Tool>.
    is static;

    Subtract(me : in out; Tool : Interval from Intrv)
    is static;

    Subtract(me : in out; Tool : Intervals from Intrv)
    is static;

    Unite(me : in out; Tool : Interval from Intrv)
    is static;

    Unite(me : in out; Tool : Intervals from Intrv)
    is static;

    XUnite(me : in out; Tool : Interval from Intrv)
    is static;

    XUnite(me : in out; Tool : Intervals from Intrv)
    is static;

    NbIntervals(me) returns Integer from Standard
    	---C++: inline
    is static;

    Value(me; Index : Integer from Standard) 
    returns Interval from Intrv
    	---C++: inline
    	---C++: return const &
    raises OutOfRange from Standard
    is static;
    
fields
    myInter : SequenceOfInterval from Intrv;

end Intervals;
