-- Created on: 2005-12-21
-- Created by: Julia GERASIMOVA
-- Copyright (c) 2005-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ComputeKronrodPointsAndWeights from math 

uses 
 
    Vector from math, 
    HArray1OfReal from TColStd

is 
    Create(Number : Integer from Standard) 
    returns ComputeKronrodPointsAndWeights; 

    IsDone(me) 
    returns Boolean from Standard;

    Points(me) 
    returns Vector from math;

    Weights(me)
    returns Vector from math;

fields 
 
    myPoints  : HArray1OfReal from TColStd;
    myWeights : HArray1OfReal from TColStd; 
    myIsDone  : Boolean from Standard;
     
end ComputeKronrodPointsAndWeights;
