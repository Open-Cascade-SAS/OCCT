-- Created on: 1993-07-06
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Curve3D from BRep inherits GCurve from BRep

	---Purpose: Representation of a curve by a 3D curve.

uses
    Pnt                 from gp,
    Location            from TopLoc,
    Curve               from Geom,
    CurveRepresentation from BRep

is

    Create(C : Curve    from Geom;
    	   L : Location from TopLoc) 
    returns mutable Curve3D from BRep;

    D0(me; U : Real; P : out Pnt from gp);
	---Purpose: Computes the point at parameter U.

    IsCurve3D(me) returns Boolean
	 ---Purpose: Returns True.
    is redefined;
	
    Curve3D(me) returns any Curve from Geom
	---C++: return const &
    is redefined;

    Curve3D(me : mutable; C : Curve from Geom)
    is redefined;
	
    Copy(me) returns mutable CurveRepresentation from BRep;
	---Purpose: Return a copy of this representation.

fields
    
    myCurve : Curve from Geom;

end Curve3D;
