-- Created on: 1996-03-07
-- Created by: Jean-Louis Frenkel
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


deferred class View from Viewer inherits TShared from MMgt
    	---Purpose: This class defines a view.        
uses
    Length from Quantity,Factor from Quantity
raises
    BadValue from Viewer
is 
    Initialize;

    Update(me)
    	---Purpose: Clears the window and redraws all primitives.
    is deferred;

  
    SetImmediateUpdate(me: mutable; onoff: Boolean from Standard)
    	---Purpose: sets the immediate update mode and returns the previous one.
    returns Boolean from Standard;
    
    ImmediateUpdate(me)
    	---Purpose: 
    is static protected;
    
    WindowFit(me: mutable ; Xmin, Ymin, Xmax, Ymax : Integer)
    	---Purpose: Centres the defined pixel window defined by the
    	-- minimum and maximum pixels Xmin, Ymin, Xmax,
    	-- Ymax so that it occupies the largest possible space
    	-- while maintaining the initial height/width ratio.
    	-- Exceptions
    	-- Viewer_BadValue if the size of the defined
    	-- projection window is equal to 0.
    raises BadValue from Viewer
    is deferred;

    Place (me:mutable; x,y: Integer from Standard;
                      aZoomFactor: Factor from Quantity = 1)
    	---Purpose: Sets the center of the object space defined by x, y
    	-- and the zoom factor aZoomFactor. The view is updated.
    is deferred;

fields

    myImmediateUpdate: Boolean from Standard is protected;


end View from Viewer;
