-- Created on: 1992-04-07
-- Created by: Christian CAILLET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



deferred class IGESEntity  from IGESData  inherits TShared

    ---Purpose : defines root of IGES Entity definition, including Directory
    --           Part, lists of (optionnal) Properties and Associativities

uses CString, Type,   HAsciiString from TCollection, OStream, GTrsf,
     EntityList,      EntityIterator,
     IGESType,   DefSwitch, DefType,      DefList,
     LineFontEntity,  LevelListEntity,    ViewKindEntity,
     TransfEntity,    LabelDisplayEntity, ColorEntity

raises InterfaceError

is

    Initialize;
    ---Purpose : prepares lists of optionnal data, set values to defaults

    Clear (me : mutable) is private;
    ---Purpose : Clears specific IGES data

    	-- --   Queries on Componants (Directory Part, optional lists)   -- --

    IGESType (me) returns IGESType;
    ---Purpose : gives IGES typing info (includes "Type" and "Form" data)

    TypeNumber (me) returns Integer;
    ---Purpose : gives IGES Type Number (often coupled with Form Number)

    FormNumber (me) returns Integer;
    ---Purpose : Returns the form number for that
    --           type of an IGES entity. The default form number is 0.


    DirFieldEntity (me; fieldnum : Integer) returns IGESEntity;
    ---Purpose : Returns the Entity which has been recorded for a given
    --           Field Number, i.e. without any cast. Maps with :
    --           3 : Structure   4 : LineFont     5 : LevelList     6 : View
    --           7 : Transf(ormation Matrix)      8 : LabelDisplay
    --           13 : Color.  Other values give a null handle
    --           It can then be of any kind, while specific items have a Type

    HasStructure (me) returns Boolean;
    ---Purpose : returns True if an IGESEntity is defined with a Structure
    --           (it is normally reserved for certain classes, such as Macros)

    Structure (me) returns IGESEntity;
    ---Purpose : Returns Structure (used by some types of IGES Entities only)
    --           Returns a Null Handle if Structure is not defined

    DefLineFont (me) returns DefType  is virtual;
    ---Purpose : Returns the definition status of LineFont

    RankLineFont (me) returns Integer;
    ---Purpose : Returns LineFont definition as an Integer (if defined as Rank)
    --           If LineFont is defined as an Entity, returns a negative value

    LineFont (me) returns LineFontEntity;
    ---Purpose : Returns LineFont as an Entity (if defined as Reference)
    --           Returns a Null Handle if DefLineFont is not "DefReference"

    DefLevel (me) returns DefList  is virtual;
    ---Purpose : Returns the definition status of Level

    Level (me) returns Integer;
    ---Purpose : Returns the level the entity
    --           belongs to. Returns -1 if the entity belongs to more than one  level.
        
    LevelList (me) returns LevelListEntity;
    ---Purpose : Returns LevelList if Level is
    --           defined as a list. Returns a null handle if DefLevel is not DefSeveral.

    DefView (me) returns DefList  is virtual;
    ---Purpose : Returns the definition status of
    --           the view. This can be: none, one or several.

    View (me) returns ViewKindEntity;
    ---Purpose : Returns the view of this IGES entity.
    --           This view can be a single view or a list of views.
    --           Warning A null handle is returned if the view is not defined.

    SingleView (me) returns ViewKindEntity;
    ---Purpose : Returns the view as a single view
    --           if it was defined as such and not as a list of views.
    --           Warning A null handle is returned if DefView does not have the value DefOne.

    ViewList (me) returns ViewKindEntity;
    ---Purpose : Returns the view of this IGES entity as a list.
    --           Warning A null handle is returned if the
    --           definition status does not have the value DefSeveral.

    HasTransf (me) returns Boolean;
    ---Purpose : Returns True if a Transformation Matrix is defined

    Transf (me) returns TransfEntity;
    ---Purpose : Returns the Transformation Matrix (under IGES definition)
    --           Returns a Null Handle if there is none
    --           for a more complete use, see Location & CompoundLocation

    HasLabelDisplay (me) returns Boolean;
    ---Purpose : Returns True if a LabelDisplay mode is defined for this entity

    LabelDisplay (me) returns LabelDisplayEntity;
    ---Purpose : Returns the Label Display
    --           Associativity Entity if there is one. Returns a null handle if there is none.

    BlankStatus (me) returns Integer;
    ---Purpose : gives Blank Status (0 visible, 1 blanked)

    SubordinateStatus (me) returns Integer;
    ---Purpose : gives Subordinate Switch (0-1-2-3)

    UseFlag (me) returns Integer;
    ---Purpose : gives Entity's Use Flag (0 to 5)

    HierarchyStatus (me) returns Integer;
    ---Purpose : gives Hierarchy status (0-1-2)

    LineWeightNumber (me) returns Integer;
    ---Purpose : Returns the LineWeight Number (0  not defined), see also LineWeight

    LineWeight (me) returns Real;
    ---Purpose : Returns the true Line Weight, computed from LineWeightNumber and
    --           Global Parameter in the Model by call to SetLineWeight

    DefColor (me) returns DefType  is virtual;
    ---Purpose : Returns the definition status of Color.

    RankColor (me) returns Integer;
    ---Purpose : Returns the color definition as
    --           an integer value if the color was defined as a rank.
    --           Warning A negative value is returned if the color was defined as an entity.

    Color (me) returns ColorEntity;
    ---Purpose : Returns the IGES entity which
-- describes the color of the entity.
-- Returns a null handle if this entity was defined as an integer.

    CResValues (me; res1,res2 : CString) returns Boolean;
    ---Purpose : returns "reserved" alphanumeric values res1 and res2
    --           res1 and res2 have to be reserved as Character[9 at least]
    --           (remark : their content is changed)
    --           returned values are ended by null character in 9th
    --           returned Boolean is False if res1 and res2 are blank, true else

    HasShortLabel (me) returns Boolean;
    ---Purpose : Returns true if a short label is defined.
    --           A short label is a non-blank 8-character string.

    ShortLabel (me) returns HAsciiString from TCollection;
    ---Purpose : Returns the label value for this IGES entity as a string.
    --           Warning If the label is blank, this string is null.

    HasSubScriptNumber (me) returns Boolean  is virtual;
    ---Purpose : Returns true if a subscript number is defined.
    --           A subscript number is an integer used to identify a label.

    SubScriptNumber (me) returns Integer;
    ---Purpose : Returns the integer subscript number used to identify this IGES entity.
    -- Warning 0 is returned if no subscript number is defined for this IGES entity.
        
    InitTypeAndForm (me : mutable; typenum,formnum : Integer)  is protected;
    ---Purpose : Initializes Type and Form Numbers to new values. Reserved for
    --           special uses

    InitDirFieldEntity (me : mutable; fieldnum : Integer; ent : IGESEntity);
    ---Purpose : Initializes a directory field as an Entiy of any kind
    --           See DirFieldEntity for more details

    InitTransf (me : mutable; ent : TransfEntity);
    ---Purpose : Initializes Transf, or erases it if <ent> is given Null

    InitView (me : mutable; ent : ViewKindEntity);
    ---Purpose : Initializes View, or erases it if <ent> is given Null

    InitLineFont (me : mutable; ent : LineFontEntity; rank : Integer = 0);
    ---Purpose : Initializes LineFont : if <ent> is not Null, it gives LineFont,
    --           else <rank> gives or erases (if zero) RankLineFont

    InitLevel (me : mutable; ent : LevelListEntity; val : Integer = 0);
    ---Purpose : Initializes Level : if <ent> is not Null, it gives LevelList,
    --           else <val> gives or erases (if zero) unique Level

    InitColor (me : mutable; ent : ColorEntity; rank : Integer = 0);
    ---Purpose : Initializes Color data : if <ent> is not Null, it gives Color,
    --           else <rank> gives or erases (if zero) RankColor

    InitStatus (me : mutable; blank, subordinate, useflag, hierarchy : Integer);
    ---Purpose : Initializes the Status of Directory Part

    SetLabel (me  : mutable; label : HAsciiString from TCollection;
              sub : Integer = -1);
    ---Purpose : Sets a new Label to an IGES Entity
    --           If <sub> is given, it sets value of SubScriptNumber
    --           else, SubScriptNumber is erased

    InitMisc (me : mutable; str : IGESEntity; lab : LabelDisplayEntity;
    	    	    	    weightnum : Integer);
    ---Purpose : Initializes various data (those not yet seen above), or erases
    --           them if they are given as Null (Zero for <weightnum>) :
    --           <str> for Structure, <lab> for LabelDisplay, and
    --           <weightnum> for WeightNumber

    	-- --    Complements (with a basic sense)    -- -- 

    HasOneParent (me) returns Boolean;
    ---Purpose : Returns True if an entity has one and only one parent, defined
    --           by a SingleParentEntity Type Associativity (explicit sharing).
    --           Thus, implicit sharing remains defined at model level
    --           (see class ToolLocation)

    UniqueParent (me) returns IGESEntity  raises InterfaceError;
    ---Purpose : Returns the Unique Parent (in the sense given by HasOneParent)
    --           Error if there is none or several

    Location (me) returns GTrsf;
    ---Purpose : Returns Location given by Transf in Directory Part (see above)
    --           It must be considered for local definition : if the Entity is
    --           set in a "Parent", that one can add its one Location, but this
    --           is not taken in account here : see CompoundLocation for that.
    --           If no Transf is defined, returns Identity
    --           If Transf is itself compound, gives the final result

    VectorLocation (me) returns GTrsf;
    ---Purpose : Returns Location considered for Vectors, i.e. without its
    --           Translation Part. As Location, it gives local definition.

    CompoundLocation (me) returns GTrsf;
    ---Purpose : Returns Location by taking in account a Parent which has its
    --           own Location : that one will be combined to that of <me>
    --           The Parent is considered only if HasOneParent is True,
    --           else it is ignored and CompoundLocation = Location

    HasName (me) returns Boolean;
    ---Purpose : says if a Name is defined, as Short Label or as Name Property
    --           (Property is looked first, else ShortLabel is considered)

    NameValue (me) returns HAsciiString from TCollection;
    ---Purpose : returns Name value as a String (Property Name or ShortLabel)
    --           if SubNumber is defined, it is concatenated after ShortLabel
    --           as follows label(number). Ignored with a Property Name

    	-- --    Optionnal lists of Associativities and Properties    -- --

    ArePresentAssociativities (me) returns Boolean;
    ---Purpose : Returns True if the Entity is defined with an Associativity
    --           list, even empty (that is, file contains its length 0)
    --           Else, the file contained NO idencation at all about this list.

    NbAssociativities (me) returns Integer;
    ---Purpose : gives number of recorded associativities (0  no list defined)

    Associativities (me) returns EntityIterator;
    ---Purpose : Returns the Associativity List under the form of an EntityIterator.

    NbTypedAssociativities (me; atype : Type) returns Integer;
    ---Purpose : gives how many Associativities have a given type

    TypedAssociativity (me; atype : Type)
    	returns mutable IGESEntity    raises InterfaceError;
    ---Purpose : returns the Associativity of a given Type (if only one exists)
    --           Error if none or more than one

    AddAssociativity (me : mutable; ent : IGESEntity) is private;
    ---Purpose : Adds an Associativity in the list (called by Associate only)

    RemoveAssociativity (me : mutable; ent : IGESEntity) is private;
    ---Purpose : Removes an Associativity from the list (called by Dissociate)

    LoadAssociativities (me : mutable; list : EntityList) is protected;
    ---Purpose : Loads a complete, already loaded, List of Asociativities
    --           (used during Read or Copy Operations)

    ClearAssociativities (me : mutable) is private;
    ---Purpose : Removes all associativities in once

    Associate (me ; ent : mutable IGESEntity);
    ---Purpose : Sets "me" in the Associativity list of another Entity

    Dissociate (me ; ent : mutable IGESEntity);
    ---Purpose : Resets "me" from the Associativity list of another Entity


    ArePresentProperties (me) returns Boolean;
    ---Purpose : Returns True if the Entity is defined with a Property list,
    --           even empty (that is, file contains its length 0)
    --           Else, the file contained NO idencation at all about this list

    NbProperties (me) returns Integer;
    ---Purpose : Gives number of recorded properties (0  no list defined)

    Properties (me) returns EntityIterator;
    ---Purpose : Returns Property List under the form of an EntityIterator

    NbTypedProperties (me; atype : Type) returns Integer;
    ---Purpose : gives how many Properties have a given type

    TypedProperty (me; atype : Type; anum : Integer = 0)
    	returns mutable IGESEntity    raises InterfaceError;
    ---Purpose : returns the Property of a given Type 
    --           Error if none or more than one

    AddProperty (me : mutable; ent : IGESEntity);
    ---Purpose : Adds a Property in the list

    RemoveProperty (me : mutable; ent : IGESEntity);
    ---Purpose : Removes a Property from the list

    LoadProperties (me : mutable; list : EntityList) is protected;
    ---Purpose : Loads a complete, already loaded, List of Properties
    --           (used during Read or Copy Operations)

    ClearProperties (me : mutable) is protected;
    ---Purpose : Removes all properties in once

    	-- --    General actions    -- --

    SetLineWeight (me : mutable; defw,maxw : Real; gradw : Integer);
    ---Purpose : computes and sets "true" line weight according IGES rules from
    --           global data MaxLineWeight (maxv) and LineWeightGrad (gradw),
    --           or sets it to defw (Default) if LineWeightNumber is null

fields
--  Entities are recorded as any, this allows special uses (with user defs)

    theType        : Integer;
    theForm        : Integer;
    theStructure   : IGESEntity;      -- used by some Entities
    theDefLineFont : DefSwitch;
    theLineFont    : IGESEntity;      -- LineFont  if Def if "Reference"
    theDefLevel    : Integer;         -- >0 (One level) =0 (None) <0 (Several)
    theLevelList   : IGESEntity;      -- LevelList  if Def is "Several"
    theView        : IGESEntity;      -- Simple View, List of Views, Null,other
    theTransf      : IGESEntity;      -- Transformation Matrix or Null
    theLabDisplay  : IGESEntity;      -- LabelDisplay .. or Null
    theStatusNum   : Integer;  -- for BlankSt,SubordinateSt,UseFlag,Hierarchy
    theLWeightNum  : Integer;         -- recorded LineWeightNumber (can be 0)
    theLWeightVal  : Real;            -- LineWeight computed from global data
    theDefColor    : DefSwitch;
    theColor       : IGESEntity;      -- ColorEntity if DefColor is "Reference"
    theRes1        : Character[9];    -- reserved for future use
    theRes2        : Character[9];
    theShortLabel  : HAsciiString from TCollection;  -- .. or Null if blank
    theSubScriptN  : Integer;         -- <0 blank, =0 given 0, >0 defined


    theAssocs : EntityList;     -- Associativity list
    theProps  : EntityList;     -- Property list

friends

    class ReadWriteModule from IGESData , class GeneralModule from IGESData ,
    class IGESReaderTool  from IGESData , class DirChecker    from IGESData

end IGESEntity;
