-- Created on: 1997-07-28
-- Created by: Pierre CHALAMET
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class TextureEnv from Graphic3d

inherits TextureRoot from Graphic3d

  ---Purpose: This class provides environment texture usable only in Visual3d_ContextView

uses

  NameOfTextureEnv from Graphic3d,
  AsciiString      from TCollection

raises

  OutOfRange from Standard

is

  Create (theFileName : AsciiString from TCollection) returns  mutable TextureEnv from Graphic3d;
  ---Purpose: Creates an environment texture from a file.

  Create (theName : NameOfTextureEnv from Graphic3d) returns mutable TextureEnv from Graphic3d;
  ---Purpose: Creates an environment texture from a predefined texture name set.

  Name (me) returns NameOfTextureEnv from Graphic3d;
  ---Purpose:
  -- Returns the name of the predefined textures or NOT_ENV_UNKNOWN
  -- when the name is given as a filename.
  ---Level: Public

  NumberOfTextures (myclass) returns Integer from Standard;
  ---Purpose:
  -- Returns the number of predefined textures.
  ---Level: Public

  TextureName (myclass; theRank: Integer from Standard)
  returns AsciiString from TCollection
  raises OutOfRange from Standard;
  ---Purpose:
  -- Returns the name of the predefined texture of rank <aRank>
  ---Trigger: when <aRank> is < 1 or > NumberOfTextures.
  ---Level: Public

fields

  myName : NameOfTextureEnv from Graphic3d;

end TextureEnv;
