-- File:	StepRepr_ShapeRepresentationRelationship.cdl
-- Created:	Tue Jun 30 18:07:23 1998
-- Author:	Christian CAILLET
--		<cky@heliox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1998


class ShapeRepresentationRelationship  from StepRepr    inherits RepresentationRelationship  from StepRepr

uses
     HAsciiString from TCollection

is

    Create returns mutable ShapeRepresentationRelationship;

end ShapeRepresentationRelationship;
