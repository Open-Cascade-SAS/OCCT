-- Created on: 1991-11-04
-- Created by: NW,JPB,CAL
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Modified:    1/08/97 ; PCT : Ajout texture mapping
--              16/01/98 ; FMN : Ajout Hiddenline
--              0312/99  ; GG : BUC60488 Why the field DistinguishModeActive
--                      field is not accessible properly ?
--                      workaround : Move the Material fields at end.
--              22/03/04 ; OCC4895 SAN High-level interface for controlling polygon offsets

class AspectFillArea3d from Graphic3d inherits AspectFillArea from Aspect

        ---Version:

        ---Purpose: This class permits the creation and updating of
        --          a graphic attribute context for opaque 3d
        --          primitives (polygons, triangles, quadrilaterals)
        --  Keywords: Face, FillArea, Triangle, Quadrangle, Polygon,
        --           TriangleMesh, QuadrangleMesh, Edge, Border, Interior,
        --           Color, Type, Width, Style, Hatch, Material,
        --           BackFaceRemoval, DistinguishMode

        ---Warning:
        ---References:

uses

        Color                 from Quantity,
        Ratio                 from Quantity,

        TypeOfLine            from Aspect,    
        InteriorStyle         from Aspect,

        MaterialAspect        from Graphic3d,
        TextureMap            from Graphic3d,

        ShaderProgram_Handle  from Graphic3d

is

        Create
                returns mutable AspectFillArea3d from Graphic3d;
        ---Level: Public
        ---Purpose: Creates a context table for fill area primitives
        --          defined with the following default values:
        --
        --          InteriorStyle       : IS_EMPTY
        --          InteriorColor       : NOC_CYAN1
        --          EdgeColor           : NOC_WHITE
        --          EdgeLineType        : TOL_SOLID
        --          EdgeWidth           : 1.0
        --          FrontMaterial       : NOM_BRASS
        --          BackMaterial        : NOM_BRASS
        --
        --          Display of back-facing filled polygons.
        --          No distinction between external and internal
        --          faces of FillAreas.
        --          The edges are not drawn.
        --          Polygon offset parameters: mode = Aspect_POM_None, factor = 1., units = 0.


        Create ( Interior       : InteriorStyle from Aspect;
                 InteriorColor  : Color from Quantity;
                 EdgeColor      : Color from Quantity;
                 EdgeLineType   : TypeOfLine from Aspect;
                 EdgeWidth      : Real from Standard;
                 FrontMaterial  : MaterialAspect from Graphic3d;
                 BackMaterial   : MaterialAspect from Graphic3d )
                returns mutable AspectFillArea3d from Graphic3d;

        ---Level: Public
        ---Purpose: Creates a context table for fill area primitives
        --          defined with the specified values.
        --
        --          Display of back-facing filled polygons.
        --          No distinction between external and internal
        --          faces of FillAreas.
        --          The edges are not drawn.
        --          Polygon offset parameters: mode = Aspect_POM_None, factor = 1., units = 0.
    	-- Warning
    	-- EdgeWidth is the "line width scale factor".   The
    	-- nominal line width is 1 pixel.   The width of the line is
    	-- determined by applying the line width scale factor to
    	-- this nominal line width.   The supported line widths
    	-- vary by 1-pixel units.

        ---------------------------------------------------
        -- Category: Methods to modify the class definition
        ---------------------------------------------------

        AllowBackFace ( me      : mutable )
                is static;
        ---Purpose: Allows the display of back-facing filled
        --          polygons.

        SetBackMaterial ( me            : mutable;
                          AMaterial     : MaterialAspect from Graphic3d )
                is static;
        ---Level: Public
        ---Purpose: Modifies the surface material of internal faces
        ---Category: Methods to modify the class definition

        SetDistinguishOn ( me   : mutable )
                is static;
        ---Level: Public
        ---Purpose: Allows distinction between external and internal
        --          faces of FillAreas.
        ---Category: Methods to modify the class definition

        SetDistinguishOff ( me  : mutable )
                is static;
        ---Level: Public
        ---Purpose: Forbids distinction between external and internal
        --          faces of FillAreas.
        ---Category: Methods to modify the class definition

        SetEdgeOn ( me  : mutable )
                is static;
        ---Level: Public
        ---Purpose: The edges of FillAreas are drawn.
        ---Category: Methods to modify the class definition

        SetEdgeOff ( me : mutable )
                is static;
        ---Level: Public
        ---Purpose: The edges of FillAreas are not drawn.
        ---Category: Methods to modify the class definition

        SetFrontMaterial ( me           : mutable;
                           AMaterial    : MaterialAspect from Graphic3d )
                is static;
        ---Level: Public
        ---Purpose: Modifies the surface material of external faces
        ---Category: Methods to modify the class definition

        SuppressBackFace ( me   : mutable )
                is static;
        ---Level: Public
        ---Purpose: Suppress the display of back-facing filled
        --          polygons.
        --          A back-facing polygon is defined as a polygon whose
        --          vertices are in a clockwise order with respect
        --          to screen coordinates.
        ---Category: Methods to modify the class definition

 
        SetTextureMap(me  :  mutable; 
                      ATexture  :  TextureMap  from Graphic3d);
 
        SetTextureMapOn(me  :  mutable);
        SetTextureMapOff(me :  mutable);

        -- 22-03-04 OCC4895 SAN High-level interface for controlling polygon offsets
        SetPolygonOffsets ( me : mutable;
                            aMode   : Integer from Standard;
                            aFactor : ShortReal from Standard = 1.0;
                            aUnits  : ShortReal from Standard = 0.0 );
        ---Level: Public
        ---Purpose: Sets up OpenGL polygon offsets mechanism.
        --          <aMode> parameter can contain various combinations of 
        --          Aspect_PolygonOffsetMode enumeration elements (Aspect_POM_None means
        --          that polygon offsets are not changed).
        --          If <aMode> is different from Aspect_POM_Off and Aspect_POM_None, then <aFactor> and <aUnits> 
        --          arguments are used by graphic renderer to calculate a depth offset value:
        --          
        --          offset = <aFactor> * m + <aUnits> * r, where
        --          m - maximum depth slope for the polygon currently being displayed,
        --          r - minimum window coordinates depth resolution (implementation-specific)
        --
        --          Deafult settings for OCC 3D viewer: mode = Aspect_POM_Fill, factor = 1., units = 0.
        --
        --          Negative offset values move polygons closer to the viewport,
        --          while positive values shift polygons away.
        --          Consult OpenGL reference for details (glPolygonOffset function description).
        ---Category: Methods to modify the class definition

        SetShaderProgram ( me  :  mutable; 
                           theProgram  :  ShaderProgram_Handle from Graphic3d );
        ---Level: Public
        ---Purpose: Sets up OpenGL/GLSL shader program.
        ---Category: Methods to modify the class definition

        ----------------------------
        -- Category: Inquire methods
        ----------------------------

        BackFace ( me )
                returns Boolean from Standard
                is static;
        ---Level: Public
        ---Purpose: Returns the Back Face Removal status.
        --          Standard_True if SuppressBackFace is activated.
        ---Category: Inquire methods

        Distinguish ( me )
                returns Boolean from Standard
                is static;
        ---Level: Public
        ---Purpose: Returns the Distinguish Mode status.
        ---Category: Inquire methods

        Edge ( me )
                returns Boolean from Standard
                is static;
        ---Level: Public
        ---Purpose: Returns Standard_True if the edges are drawn and
        --          Standard_False if the edges are not drawn.
        ---Category: Inquire methods

        BackMaterial ( me )
                returns MaterialAspect from Graphic3d
                is static;
        ---Level: Public
        ---Purpose: Returns the surface material of internal faces
        ---Category: Inquire methods

        FrontMaterial ( me )
                returns MaterialAspect from Graphic3d
                is static;
        ---Level: Public
        ---Purpose: Returns the surface material of external faces
        ---Category: Inquire methods

 
        TextureMap(me) 
            returns  TextureMap  from  Graphic3d; 
             
        TextureMapState(me) 
            returns  Boolean  from  Standard;

        -- 22-03-04 OCC4895 SAN High-level interface for controlling polygon offsets
        PolygonOffsets ( me;
                         aMode   : out Integer from Standard;
                         aFactor : out ShortReal from Standard;
                         aUnits  : out ShortReal from Standard );
        ---Level: Public
        ---Purpose: Returns current polygon offsets settings.
        ---Category: Inquire methods

        ShaderProgram ( me )
        returns ShaderProgram_Handle from Graphic3d;
        ---C++: return const &

--

fields

--
-- Class        :       Graphic3d_AspectFillArea3d
--
-- Purpose      :       Declaration of variables specific to
--                      the context of drawing 3d faces
--
-- Reminder     :       A context for drawing 3d faces inherits a context
--                      defined by :
--                      - the interior style of the face
--                      - the edge style of the face
--                      - the colour
--                      It also possesses a definition of the materials for the
--                      internal and external faces.
--
--


        -- flag to distinguish between internal and external faces
        DistinguishModeActive   :       Boolean from Standard;

        -- flag to draw the edges or not
        EdgeModeActive          :       Boolean from Standard;

        -- display flag for reversed polygons.
        BackFaceRemovalActive   :       Boolean from Standard;

        MyTextureMap            :       TextureMap  from  Graphic3d; 
        MyTextureMapState       :       Boolean  from  Standard;

        -- the material
        MyFrontMaterial         :       MaterialAspect from Graphic3d;
        MyBackMaterial          :       MaterialAspect from Graphic3d;

        -- 22-03-04 OCC4895 SAN High-level interface for controlling polygon offsets
        -- polygon offsets
        MyPolygonOffsetMode     :       Integer from Standard;
        MyPolygonOffsetFactor   :       ShortReal from Standard;
        MyPolygonOffsetUnits    :       ShortReal from Standard;

        MyShaderProgram         :       ShaderProgram_Handle  from  Graphic3d;

end AspectFillArea3d;
