-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SelectorOfDataStructureOfDelaun from BRepMesh

  ---Purpose: Describes a selector and  an Iterator on a
  --          selector of components of a Mesh.

  uses    Integer from Standard,
          Box from Bnd,
          MapOfInteger from BRepMesh,
          DataStructureOfDelaun from BRepMesh,
          Vertex from BRepMesh,
          Edge from BRepMesh,
          Triangle from BRepMesh

is          Create returns SelectorOfDataStructureOfDelaun from BRepMesh;

            Create      (theMesh     : DataStructureOfDelaun from BRepMesh)
            returns SelectorOfDataStructureOfDelaun from BRepMesh;

            Initialize   (me          : in out;
                          theMesh     :DataStructureOfDelaun from BRepMesh) 
            is static;


            NeighboursOf(me          : in out;
                         theNode     : in Vertex from BRepMesh) 
              is static;

            NeighboursOfNode(me          : in out;
                             indexNode   : in Integer from Standard) 
              is static;


            NeighboursOf(me          : in out;
                         theLink     : in Edge from BRepMesh) 
              is static;

            NeighboursOfLink(me          : in out;
                             indexLink   : in Integer from Standard) 
              is static;


            NeighboursOf(me          : in out;
                         theElem     : in Triangle from BRepMesh) 
              is static;

            NeighboursOfElement(me        : in out;
                                indexElem : in Integer from Standard) 
            ---Purpose: All Neighbours  Of the Element. By
            --          edge or by vertices.
              is static;


            NeighboursByEdgeOf (me        : in out;
                                theElem   : in Triangle from BRepMesh) 
              ---Purpose: Neighbours by edge Of the Element.
              is static;


            NeighboursOf(me          : in out;
                         theSelector : in SelectorOfDataStructureOfDelaun from BRepMesh) 
                ---Purpose: Adds a level of Neighbours by edge
                --          to the selector <theSelector>.
                is static;


            AddNeighbours(me       : in out)
              ---Purpose: Adds a level of Neighbours by edge
              --          to the selector <me>.
              is static;


            Nodes       (me) 
              ---C++: return const &
              returns  MapOfInteger from BRepMesh is static;

            Links       (me) 
              ---C++: return const &
              returns  MapOfInteger from BRepMesh is static;

            Elements    (me) 
              ---C++: return const &
              returns  MapOfInteger from BRepMesh is static;

            FrontierLinks(me) 
              ---Purpose: Gives the  list  of links  incices
              --          frontier  of  the  selector  <me>.
              ---C++: return const &
              returns  MapOfInteger from BRepMesh is static;


              fields  myMesh      :DataStructureOfDelaun from BRepMesh;
                      myNodes     : MapOfInteger from BRepMesh;
                      myLinks     : MapOfInteger from BRepMesh;
                      myElements  : MapOfInteger from BRepMesh;
                      myFrontier  : MapOfInteger from BRepMesh;

end SelectorOfDataStructureOfDelaun;
