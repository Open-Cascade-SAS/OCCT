-- Created on: 1996-04-09
-- Created by: Joelle CHAUVET
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Node from AdvApp2Var
    ---Purpose :
    -- used to store constraints on a (Ui,Vj) point
    --

uses
    XY,Pnt           from gp,
    HArray2OfPnt     from TColgp,
    HArray2OfReal    from TColStd
    
	 
is
    Create returns Node;    
    Create(iu,iv : Integer) returns Node;   
    Create(UV : XY from gp; iu,iv : Integer) returns Node;    
    Create(Other : Node) returns Node is private;    
    Coord(me) returns XY from gp;    
    SetCoord(me : in out; x1,x2 : Real);    
    UOrder(me) returns Integer;
    VOrder(me) returns Integer;
    SetPoint(me : in out; iu,iv : Integer; Cte : Pnt from gp);    
    Point(me; iu,iv : Integer) returns Pnt from gp;    
    SetError(me : in out; iu,iv : Integer; error : Real);    
    Error(me; iu,iv : Integer) returns Real;     
    
    
fields

    myCoord            : XY               from gp;
    myOrdInU, myOrdInV : Integer;
    myTruePoints       : HArray2OfPnt     from TColgp;
    myErrors           : HArray2OfReal    from TColStd;
    
end Node;







