-- Created on: 1992-11-18
-- Created by: Christian CAILLET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class SelectDiff  from IFSelect  inherits SelectControl

    ---Purpose : A SelectDiff keeps the entities from a Selection, the Main
    --           Input, which are not listed by the Second Input

uses AsciiString from TCollection, EntityIterator, Graph

is

    Create returns mutable SelectDiff;
    ---Purpose : Creates an empty SelectDiff


    RootResult (me; G : Graph) returns EntityIterator;
    ---Purpose : Returns the list of selected entities : they are the Entities
    --           gotten from the Main Input but not from the Diff Input

    HasUniqueResult (me) returns Boolean  is redefined protected;
    ---Purpose : Returns always True, because RootResult gives a Unique list


    Label (me) returns AsciiString from TCollection;
    ---Purpose : Returns a text defining the criterium : "Difference"

end SelectDiff;
