-- Created on: 1995-12-04
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class RWViewVolume from RWStepVisual

	---Purpose : Read & Write Module for ViewVolume

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     ViewVolume from StepVisual,
     EntityIterator from Interface

is

	Create returns RWViewVolume;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable ViewVolume from StepVisual);

	WriteStep (me; SW : in out StepWriter; ent : ViewVolume from StepVisual);

	Share(me; ent : ViewVolume from StepVisual; iter : in out EntityIterator);

end RWViewVolume;
