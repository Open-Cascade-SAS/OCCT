-- Created on: 1999-04-15
-- Created by: Denis PASCAL
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DocumentRetrievalDriver from MDocStd inherits RetrievalDriver from PCDM

	---Purpose: retrieval driver of a standard document

uses Document         from TDocStd,
     Document         from PDocStd,  
     RRelocationTable from MDF,
     Document         from PCDM, 
     Document         from CDM,  
     MessageDriver    from CDM,
     ExtendedString   from TCollection,
     ARDriverTable    from MDF

is


    Create
    returns mutable DocumentRetrievalDriver from MDocStd;    

    Paste (me : mutable; PDOC   : Document from PDocStd;
                         TDOC   : Document from TDocStd;
			 aReloc : RRelocationTable from MDF);
    
    ---Purpose: deferred methods of RetrievalDriver from PCDM
    --          =============================================

    Make (me : mutable; aPCDM: Document from PCDM; aCDM : mutable Document from CDM); 

    ---Purpose: virtual methods (may be redefined by specialized application)
    --          =============================================================

    SchemaName(me) returns ExtendedString from  TCollection
    is virtual;

    CreateDocument (me: mutable) returns Document from CDM  
    ---Purpose: returns an empty TDocStd_Document. may be redefined;
    is virtual;
    
    AttributeDrivers(me : mutable; theMessageDriver : MessageDriver from CDM) 
    returns ARDriverTable from MDF
    is virtual;
    
fields

    myDrivers : ARDriverTable  from MDF;

end DocumentRetrievalDriver;
