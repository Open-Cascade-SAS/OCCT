-- Created on: 1996-12-05
-- Created by: Jean-Pierre COMBE/Odile Olivier
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class PerpendicularRelation from AIS inherits Relation from AIS
    	---Purpose: A framework to display constraints of perpendicularity
    	-- between two or more interactive datums. These
    	-- datums can be edges or faces.
uses Shape                 from TopoDS,
     Presentation          from Prs3d,
     PresentationManager3d from PrsMgr,
     Selection             from SelectMgr,
     Pnt                   from gp,
     Dir                   from gp,
     Projector             from Prs3d,
    Transformation        from Geom,
     PresentationManager2d from PrsMgr,
     GraphicObject         from Graphic2d,     
     Plane                 from Geom

is
    Create (aFShape     : Shape          from TopoDS;
    	    aSShape     : Shape          from TopoDS;
	    aPlane      : Plane          from Geom)
	---Purpose:  Constructs an object to display constraints of
    	-- perpendicularity on shapes.
    	-- This object is defined by a first shape aFShape, a
    	-- second shape aSShape, and a plane aPlane.
    	-- aPlane is the plane of reference to show and test the
    	-- perpendicular relation between two shapes, at least
    	-- one of which has a revolved surface.
    returns mutable PerpendicularRelation from AIS;

    Create (aFShape     : Shape          from TopoDS;
    	    aSShape     : Shape          from TopoDS)
	---Purpose:  Constructs an object to display constraints of
    	-- perpendicularity on shapes.
    	-- This object is defined by a first shape aFShape and a
    	-- second shape aSShape.
    returns mutable PerpendicularRelation from AIS;

-- -- Methods from PresentableObject

    Compute(me            : mutable;
    	    aPresentationManager: PresentationManager3d from PrsMgr;
    	    aPresentation : mutable Presentation from Prs3d;
    	    aMode         : Integer from Standard= 0) 
    is redefined static private;
    
    Compute(me:mutable;
    	        aProjector: Projector from Prs3d;
                aPresentation: mutable Presentation from Prs3d)
    is redefined static private;     

    Compute(me:mutable;
    	    aPresentationManager: PresentationManager2d from PrsMgr;
            aPresentation: mutable GraphicObject from Graphic2d;
            aMode: Integer from Standard = 0)
    is redefined static private;	    

    Compute(me            : mutable;
    	    aProjector    : Projector from Prs3d;
    	    aTrsf         : Transformation from Geom;
	    aPresentation : mutable Presentation from Prs3d)
    is redefined;
    	---Purpose: computes the presentation according to a point of view
    	--          given by <aProjector>. 
    	--          To be Used when the associated degenerated Presentations 
    	--          have been transformed by <aTrsf> which is not a Pure
    	--          Translation. The HLR Prs can't be deducted automatically
    	--          WARNING :<aTrsf> must be applied
    	--           to the object to display before computation  !!!

-- Methods from SelectableObject

    ComputeSelection(me         : mutable;
    	    	     aSelection : mutable Selection from SelectMgr;
    	    	     aMode      : Integer from Standard)is private;


--
--     Computation private methods
--

    ComputeTwoFacesPerpendicular(me: mutable;
    	    	    	         aPresentation : mutable Presentation from Prs3d)
    is private;
    
    ComputeTwoEdgesPerpendicular(me: mutable;
    	    	    	         aPresentation : mutable Presentation from Prs3d)
    is private;
    

fields

    myFAttach     : Pnt from gp;
    mySAttach     : Pnt from gp;
    
end PerpendicularRelation;


