-- Created on: 1998-06-04
-- Created by: Philippe NOUAILLE
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ChAsymInv from BlendFunc 

inherits FuncInv from Blend

uses Vector   from math,
     Matrix   from math,
     HCurve2d from Adaptor2d,
     HCurve   from Adaptor3d,
     HSurface from Adaptor3d

is
    Create(S1,S2: HSurface from Adaptor3d; C: HCurve from Adaptor3d)
    
    	returns ChAsymInv from BlendFunc;
	
    Set(me: in out; OnFirst: Boolean from Standard;
    	            COnSurf: HCurve2d from Adaptor2d)

    	;


    GetTolerance(me; Tolerance: out Vector from math; Tol: Real from Standard)
    
    	;


    GetBounds(me; InfBound,SupBound: out Vector from math)
    
    	;


    IsSolution(me: in out; Sol: Vector from math; Tol: Real from Standard)
    
    	returns Boolean from Standard
    
    	;


    NbEquations(me)
    	---Purpose: returns the number of equations of the function.
    	returns Integer from Standard
    	is redefined static ;

    ComputeValues(me   : in out;
                  X    : Vector from math;
                  DegF : Integer from Standard;
		  DegL : Integer from Standard)
    ---Purpose: computes the values <F> of the derivatives for the 
    --          variable <X> between DegF and DegL.
    --          Returns True if the computation was done successfully, 
    --          False otherwise.
    returns Boolean from Standard
    is static;

    Value(me: in out; X: Vector; F: out Vector)
    	---Purpose: computes the values <F> of the Functions for the 
    	--          variable <X>.
    	--          Returns True if the computation was done successfully, 
    	--          False otherwise.

    	returns Boolean from Standard
    	is redefined static ;
    
    
    Derivatives(me: in out; X: Vector; D: out Matrix)
    	---Purpose: returns the values <D> of the derivatives for the 
    	--          variable <X>.
    	--          Returns True if the computation was done successfully, 
    	--          False otherwise.

    returns Boolean from Standard
    is redefined static	;
    
    
    Values(me: in out; X: Vector; F: out Vector; D: out Matrix)
    	---Purpose: returns the values <F> of the functions and the derivatives
    	--          <D> for the variable <X>.
    	--          Returns True if the computation was done successfully, 
    	--          False otherwise.

    returns Boolean from Standard
    	is redefined static ;

-- methodes hors template (en plus du create)

    Set(me: in out; 
        Dist1 : Real from Standard;
	Angle : Real from Standard;
        Choix : Integer from Standard)

    is static;


fields

    surf1 : HSurface from Adaptor3d;
    surf2 : HSurface from Adaptor3d;
    dist1 : Real from Standard;
    angle : Real from Standard;
    tgang : Real from Standard;
    curv  : HCurve from Adaptor3d;
    csurf : HCurve2d from Adaptor2d;
    choix : Integer from Standard;
    first : Boolean from Standard;

    FX       : Vector  from math;
    DX       : Matrix  from math;
    
end ChAsymInv;
