-- Created on: 1993-01-28
-- Created by: Gilles DEBARBOUILLE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class InterpretedMethod from Dynamic

inherits

    MethodDefinition from Dynamic

	---Purpose: This class derived from Method, describes an  
	--          interpreted method. The additional field is the 
	--          name of the file to be interpreted.

uses

    CString from Standard,
    HAsciiString from TCollection,
    AsciiString  from TCollection

is

    Create(aname , afile : CString from Standard) returns mutable InterpretedMethod from Dynamic;
    
    ---Level: Public 
    
    ---Purpose: Creates a new  InterpretedMethod with <aname> as  name
    --          and <afile> as file name to be interpreted.
    
    Function(me : mutable ; afile : CString from Standard)
    
    ---Level: Public 
    
    ---Purpose: Sets the the   name of the  file to  be interpreted to
    --          <afile>.
    
    is static;
    
    Function(me) returns AsciiString from TCollection
    
    ---Level: Public 
    
    ---Purpose: Returns the name of the file to be interpreted.
    
    is static;
    
fields

    thefunction : HAsciiString from TCollection;

end InterpretedMethod;
