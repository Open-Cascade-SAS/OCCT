-- Created on: 1994-01-10
-- Created by: Yves FRICAUD
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PointOnBis from Bisector 

	---Purpose: 
    
uses 
    Pnt2d from gp

is
    Create returns PointOnBis from Bisector;
    
    Create ( Param1, Param2, ParamBis, Distance : Real; Point : Pnt2d) 
    returns PointOnBis from Bisector; 
    
    ParamOnC1 (me : in out; Param : Real)
    is static;
    
    ParamOnC2 (me : in out; Param : Real)
    is static;
    
    ParamOnBis (me : in out; Param : Real)
    is static;
    
    Distance (me : in out; Distance : Real)
    is static;
    
    IsInfinite (me : in out; Infinite : Boolean)
    is static;

    Point (me : in out ; P :Pnt2d)
    is static;
    
    ParamOnC1 (me) returns Real
    is static;
    
    ParamOnC2 (me) returns Real
    is static;

    ParamOnBis (me) returns Real
    is static;
        
    Distance (me) returns Real
    is static;
    
    Point (me) returns Pnt2d
    is static;
    
    IsInfinite (me) returns Boolean 
    is static;
    
    Dump (me) is static;
    
fields

    param1   : Real;
    param2   : Real;
    paramBis : Real;
    distance : Real;
    infinite : Boolean;	
    point    : Pnt2d from gp;
    
end PointOnBis;
