-- Created on: 1992-02-04
-- Created by: Laurent PAINNOT
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

generic class SingleTab from math (Item as any)
uses Address from Standard
is

    Create(LowerIndex, UpperIndex: Integer)
       returns SingleTab;    	
    
    Create(Tab : Item; LowerIndex, UpperIndex: Integer)
       returns SingleTab;    	
    
    Init(me : in out;  InitValue: Item) is static;

    Create(Other: SingleTab)
    	returns SingleTab;
	
    Copy(me; Other : in out SingleTab)
    	---C++: inline
    is static;

    SetLower(me: in out; LowerIndex : Integer)
    is static;
    
    Value(me; Index: Integer)
    	---C++: alias operator()
    	---C++: return &
    	---C++: inline
       returns Item
    is static;


    Free(me: in out)
    	---C++: alias ~

    is static;

fields

Addr        : Address;
Buf         : Item[512];
isAllocated : Boolean;
First       : Integer;
Last        : Integer;

end;

