-- Created on: 2008-12-10
-- Created by: Pavel TELKOV
-- Copyright (c) 2008-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Material from PXCAFDoc inherits  Attribute from PDF

	---Purpose: 
uses
    Real          from Standard,
    HAsciiString  from PCollection
is
    Create returns mutable Material from PXCAFDoc;

    Create (theName       : HAsciiString from PCollection;
    	    theDescr      : HAsciiString from PCollection;
	    theDensity    : Real         from Standard;
    	    theDensName   : HAsciiString from PCollection;
    	    theDensValType: HAsciiString from PCollection)
    returns mutable Material from PXCAFDoc;
    
    GetName (me) returns HAsciiString from PCollection;

    GetDescription (me) returns HAsciiString from PCollection;

    GetDensity (me) returns Real from Standard;

    GetDensName (me) returns HAsciiString from PCollection;

    GetDensValType (me) returns HAsciiString from PCollection;

    Set (me : mutable; theName       : HAsciiString from PCollection;
                       theDescr      : HAsciiString from PCollection;
                       theDensity    : Real         from Standard;
                       theDensName   : HAsciiString from PCollection;
                       theDensValType: HAsciiString from PCollection);
    
fields

    myName        : HAsciiString from PCollection;
    myDescr       : HAsciiString from PCollection;
    myDensity     : Real from Standard;
    myDensName    : HAsciiString from PCollection;
    myDensValType : HAsciiString from PCollection;

end Material from PXCAFDoc;
