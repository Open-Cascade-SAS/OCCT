-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class TrimmedCurve from StepGeom 

inherits BoundedCurve from StepGeom 

uses

	Curve from StepGeom, 
	HArray1OfTrimmingSelect from StepGeom, 
	Boolean from Standard, 
	TrimmingPreference from StepGeom, 
	TrimmingSelect from StepGeom, 
	HAsciiString from TCollection
is

	Create returns mutable TrimmedCurve;
	---Purpose: Returns a TrimmedCurve


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aBasisCurve : mutable Curve from StepGeom;
	      aTrim1 : mutable HArray1OfTrimmingSelect from StepGeom;
	      aTrim2 : mutable HArray1OfTrimmingSelect from StepGeom;
	      aSenseAgreement : Boolean from Standard;
	      aMasterRepresentation : TrimmingPreference from StepGeom) is virtual;

	-- Specific Methods for Field Data Access --

	SetBasisCurve(me : mutable; aBasisCurve : mutable Curve);
	BasisCurve (me) returns mutable Curve;
	SetTrim1(me : mutable; aTrim1 : mutable HArray1OfTrimmingSelect);
	Trim1 (me) returns mutable HArray1OfTrimmingSelect;
	Trim1Value (me; num : Integer) returns TrimmingSelect;
	NbTrim1 (me) returns Integer;
	SetTrim2(me : mutable; aTrim2 : mutable HArray1OfTrimmingSelect);
	Trim2 (me) returns mutable HArray1OfTrimmingSelect;
	Trim2Value (me; num : Integer) returns TrimmingSelect;
	NbTrim2 (me) returns Integer;
	SetSenseAgreement(me : mutable; aSenseAgreement : Boolean);
	SenseAgreement (me) returns Boolean;
	SetMasterRepresentation(me : mutable; aMasterRepresentation : TrimmingPreference);
	MasterRepresentation (me) returns TrimmingPreference;

fields

	basisCurve : Curve from StepGeom;
	trim1 : HArray1OfTrimmingSelect from StepGeom; -- a SelectType
	trim2 : HArray1OfTrimmingSelect from StepGeom; -- a SelectType
	senseAgreement : Boolean from Standard;
	masterRepresentation : TrimmingPreference from StepGeom; -- an Enumeration

end TrimmedCurve;
