-- Created on: 1996-12-25
-- Created by: Alexander BRIVIN
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Cylinder from Vrml 

	---Purpose: defines a Cylinder node of VRML specifying geometry shapes.
    	-- This  node  represents  a  simple  capped  cylinder  centred  around the  y-axis. 
    	-- By  default ,  the  cylinder  is  centred  at  (0,0,0) 
	-- and  has  size  of  -1  to  +1  in  the  all  three  dimensions. 
	-- The  cylinder  has  three  parts: 
	-- the  sides,  the  top  (y=+1)  and  the  bottom (y=-1)

uses
 
    CylinderParts from Vrml

is

    Create ( aParts  : CylinderParts from Vrml  = Vrml_CylinderALL;
    	     aRadius : Real          from Standard = 1;
	     aHeight : Real          from Standard = 2 )
        returns Cylinder from Vrml;

    SetParts ( me : in out; aParts : CylinderParts from Vrml );
    Parts ( me  )  returns CylinderParts from Vrml;
    
    SetRadius ( me : in out; aRadius : Real from Standard );
    Radius ( me )  returns Real  from  Standard;
  
    SetHeight ( me : in out; aHeight : Real from Standard );
    Height ( me )  returns Real  from  Standard;

    Print  ( me;  anOStream: in out OStream from Standard) returns OStream from Standard;
    ---C++:  return  & 

fields

    myParts  : CylinderParts from Vrml; -- Visible parts of cylinder
    myRadius : Real from Standard;      -- Radius in x and z dimensions
    myHeight : Real from Standard;      -- Size in y dimension
    
end Cylinder;
