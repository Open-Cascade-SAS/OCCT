-- File:        ContextDependentShapeRepresentation.cdl
-- Created:     Mon Dec  4 12:02:23 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWContextDependentShapeRepresentation from RWStepShape

	---Purpose : Read & Write Module for ContextDependentShapeRepresentation

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     ContextDependentShapeRepresentation from StepShape,
     EntityIterator from Interface

is

    Create returns RWContextDependentShapeRepresentation;

    ReadStep (me; data : StepReaderData; num : Integer; ach : in out Check;
                  ent : mutable ContextDependentShapeRepresentation from StepShape);

    WriteStep (me; SW : in out StepWriter; ent : ContextDependentShapeRepresentation from StepShape);

    Share(me; ent : ContextDependentShapeRepresentation from StepShape; iter : in out EntityIterator);

end RWContextDependentShapeRepresentation;
