-- Created on: 1999-09-13
-- Created by: data exchange team
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class FixSmallFace from ShapeFix inherits Root from ShapeFix

	---Purpose: 

uses
    Shape from TopoDS,
    Face from TopoDS,
    Edge from TopoDS,
    Compound from TopoDS,
    CheckSmallFace from ShapeAnalysis
    
is
    Create returns FixSmallFace;
    ---Purpose :
    Init(me: mutable; S : Shape from TopoDS); 
    ---Purpose :
    
    Perform(me:mutable);	
    ---Purpose :
    -- Fixing case of spot face
    FixSpotFace (me: mutable) returns Shape from TopoDS;
    ---Purpose : Fixing case of spot face, if tol = -1 used local tolerance.
    ReplaceVerticesInCaseOfSpot(me; F : in out Face from TopoDS; tol : Real) returns Boolean;
    ---Purpose : Compute average vertex and replacing vertices by new one.

     RemoveFacesInCaseOfSpot(me; F :  Face from TopoDS) returns Boolean;
    ---Purpose : Remove spot face from compound
    --
    
     -- Fixing case of strip face   
     FixStripFace(me: mutable; wasdone: Boolean = Standard_False) returns Shape from TopoDS;
    ---Purpose : Fixing case of strip face, if tol = -1 used local tolerance

    ReplaceInCaseOfStrip(me;F : in out Face from TopoDS; E1 : in out  Edge from TopoDS; E2 : in out  Edge from TopoDS;tol : Real) returns Boolean;
    ---Purpose : Replace veretces and edges.
    --
    RemoveFacesInCaseOfStrip(me; F :  Face from TopoDS) returns Boolean;
    ---Purpose : Remove strip face from compound.
    
    ComputeSharedEdgeForStripFace(me; F :  Face from TopoDS; E1 : Edge from TopoDS; E2 : Edge from TopoDS; 
    F1 :  Face from TopoDS;     tol : Real ) 
    returns Edge from TopoDS;
    ---Purpose : Compute average edge for strip face

     -- Fixing case split
    
    FixSplitFace(me: mutable; S: Shape from TopoDS) returns Shape from TopoDS;
    ---Purpose : 
    --
    
    SplitFaces(me: mutable) returns Shape from TopoDS;
    ---Purpose : Split faces by splitting vertices
    --
    
    SplitOneFace(me: mutable; F : in out Face from TopoDS;theSplittedFaces: in out Compound from TopoDS) returns Boolean;
    ---Purpose : Compute data for face splitting.
    --
    
    RemoveSmallFaces(me:mutable) returns Shape from TopoDS;
    ---Purpose : Remove small faces from compound.
  
    --Fixes after removing
    FixFace(me: mutable; F: Face from TopoDS) returns Face from TopoDS;
    FixShape(me: mutable) returns Shape from TopoDS;

    Shape(me : mutable) returns Shape from TopoDS;
    
    FixPinFace (me: mutable;F : in out Face from TopoDS) returns Boolean;

fields

    myShape    : Shape from TopoDS;
    myResult   : Shape from TopoDS;
    myStatus   : Integer; -- error status
    myAnalyzer : CheckSmallFace from ShapeAnalysis;




end FixSmallFace;
