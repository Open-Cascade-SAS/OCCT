-- Created on: 2001-09-11
-- Created by: Julia DOROVSKIKH
-- Copyright (c) 2001-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


package XmlMXCAFDoc

        ---Purpose: Storage and Retrieval drivers for modelling attributes.
        --          Transient attributes are defined in package XCAFDoc

uses TopLoc,
     XmlMDF,
     XmlObjMgt,
     TDF,
     CDM,
     TopTools

is
    class AreaDriver;

    class CentroidDriver;

    class ColorDriver;

    class GraphNodeDriver;

    class LocationDriver;

    class VolumeDriver;

    class DatumDriver;
    class DimTolDriver;
    class MaterialDriver;

    class ColorToolDriver;
    class DocumentToolDriver;
    class LayerToolDriver;
    class ShapeToolDriver;
    class DimTolToolDriver;
    class MaterialToolDriver;

    AddDrivers (aDriverTable : ADriverTable  from XmlMDF;
                anMsgDrv     : MessageDriver from CDM);
        ---Purpose: Adds the attribute drivers to <aDriverTable>.

end XmlMXCAFDoc;
