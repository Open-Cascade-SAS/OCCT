-- Created on: 1998-06-03
-- Created by: data exchange team
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ShellSewing from ShapeUpgrade 

    ---Purpose: This class provides a tool for applying sewing algorithm from
    --          BRepAlgo: it takes a shape, calls sewing for each shell, 
    --          and then replaces sewed shells with use of ShapeBuild_ReShape

uses 
    Shape from TopoDS,
    IndexedMapOfShape from TopTools,
    ReShape from ShapeBuild

is

    Create returns ShellSewing;
    ---Purpose: Creates a ShellSewing, empty

    ApplySewing (me: in out; shape: Shape from TopoDS; tol: Real = 0.0)
    	returns Shape from TopoDS;
    ---Purpose: Builds a new shape from a former one, by calling Sewing from
    --          BRepOffsetAPI. Rebuilt solids are oriented to be "not infinite"
    --           
    --          If <tol> is not given (i.e. value 0. by default), it is
    --          computed as the mean tolerance recorded in <shape>
    --           
    --          If no shell has been sewed, this method returns the input
    --          shape

    Init (me: in out; shape: Shape from TopoDS) is private;

    Prepare (me: in out; tol: Real) returns Integer is private;
    
    Apply (me: in out; shape: Shape from TopoDS; tol: Real) 
    returns Shape from TopoDS is private;
    
fields

    myShells: IndexedMapOfShape from TopTools;
    myReShape: ReShape from ShapeBuild;

end ShellSewing;
