-- Created by: Tanya COOL
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Repere from Prs2d inherits Dimension from Prs2d

 ---Purpose: Constructs the repere

uses

	Drawer		       from Graphic2d,
	GraphicObject	   from Graphic2d,
	Pnt2d              from gp,
	ExtendedString     from TCollection,
	Array1OfShortReal  from TShort,
    	ArrowSide          from Prs2d,
	TypeOfArrow        from Prs2d,
    	FStream            from Aspect 

is
	Create( aGO           : GraphicObject  from Graphic2d;
	        aPnt1         : Pnt2d          from gp;
            	aPnt2         : Pnt2d          from gp;
		aLenBase      : Real           from Standard; 
		aText         : ExtendedString from TCollection;
       	    	aTxtScale     : Real           from Standard = 1.0;
            	aDrawArrow    : Boolean        from Standard = Standard_False; 
            	anArrAngle    : Real           from Standard = 10.0;
		anArrLength   : Real           from Standard = 10.0;
            	anArrType     : TypeOfArrow    from Prs2d    = Prs2d_TOA_OPENED;
		anArrow       : ArrowSide      from Prs2d    = Prs2d_AS_BOTHAR;
		IsRevArrow    : Boolean        from Standard = Standard_False ) 

	returns mutable Repere from Prs2d;
    	---Level: Public
    	---Purpose: Creates repere 

	-------------------------------------------------
	-- Category: Draw and Pick
	-------------------------------------------------

	Draw( me : mutable; aDrawer: Drawer from Graphic2d ) is static protected;
	---Level: Internal
	---Purpose: Draws the repere <me>.

    	DrawElement( me : mutable; aDrawer: Drawer from Graphic2d;
            	     anIndex: Integer from Standard)
            is redefined protected;
    	---Level: Internal
    	---Purpose: 

    	DrawVertex( me : mutable; aDrawer: Drawer from Graphic2d;
                    anIndex: Integer from Standard)
            is redefined protected;
    	---Level: Internal
    	---Purpose: 

    	Pick( me : mutable; X, Y: ShortReal from Standard;
       	      aPrecision: ShortReal from Standard;
	      aDrawer: Drawer from Graphic2d ) 
    	returns Boolean from Standard is static protected;
	---Level: Internal
	---Purpose: Returns Standard_True if the repere <me> is picked,
	--	    Standard_False if not.

	Save( me; aFStream: in out FStream from Aspect ) is virtual;
													
    	CalcTxtPos(me:mutable; theFromAbs: 
    	    	    Boolean from Standard) 
    	---C++: inline
    	is redefined protected;

fields 
 
    myXVert        : Array1OfShortReal from TShort;
    myYVert        : Array1OfShortReal from TShort;
    myObtuse       : Boolean           from Standard;
    myDrawArrow    : Boolean           from Standard;

end Repere from Prs2d;
