-- Created on: 2005-05-17
-- Created by: Eugeny NAPALKOV <eugeny.napalkov@opencascade.com>
-- Copyright (c) 2005-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ColorToolDriver from BinMXCAFDoc inherits ADriver from BinMDF

uses
    MessageDriver    from CDM,
    SRelocationTable from BinObjMgt,
    RRelocationTable from BinObjMgt,
    Persistent       from BinObjMgt,
    Attribute        from TDF

is
    Create (theMsgDriver:MessageDriver from CDM)
    returns ColorToolDriver from BinMXCAFDoc;

    NewEmpty (me)  returns Attribute from TDF
    is redefined;

    Paste(me; theSource     : Persistent from BinObjMgt;
              theTarget     : Attribute from TDF;
              theRelocTable : out RRelocationTable from BinObjMgt)
    returns Boolean from Standard is redefined;

    Paste(me; theSource     : Attribute from TDF;
              theTarget     : in out Persistent from BinObjMgt;
              theRelocTable : out SRelocationTable from BinObjMgt)
    is redefined;

end;

