-- File:	Contap_ArcTool.cdl
-- Created:	Wed May 12 09:09:34 1993
-- Author:	Jacques GOUSSARD
--		<jag@topsn2>
---Copyright:	 Matra Datavision 1993



deferred generic class ArcTool from Contap
    (TheArc as any )


    ---Purpose: Template class for a tool on the restriction of
    --          a surface.
    -- It is possible to implement this class with an instantiation
    -- of the class CurveTool from Adaptor3d.


uses Pnt2d from gp,
     Vec2d from gp

is

    Value(myclass; A: TheArc; X: Real from Standard)
    
	---Purpose: Returns the value in the parametric space
	--          of the surface S, of the point of parameter X
	--          on the arc A.

    	returns Pnt2d from gp;


    D1(myclass; A: TheArc; X: Real from Standard;
                P      : out Pnt2d from gp;
                D2D    : out Vec2d from gp);
    
	---Purpose: Returns the value and the first derivatives in
	--          the parametric space of the surface S of the point
	--          at parameter X on the arc A.


    Resolution(myclass; A: TheArc; Tol3d: Real from Standard)

        ---Purpose :  Returns the parametric resolution corresponding
        --         to the space resolution Tol3d.

    	returns Real from Standard;


end ArcTool;


