-- Created on: 2000-09-29
-- Created by: Pavel TELKOV
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class GraphNode from PXCAFDoc inherits Attribute from PDF

	---Purpose: 

uses
    Attribute         from PDF,
    GUID              from Standard,
    GraphNodeSequence from PXCAFDoc

is
    Create returns mutable GraphNode from PXCAFDoc;
    
    SetFather (me : mutable;F : GraphNode from PXCAFDoc)
    returns Integer from Standard;

    SetChild (me : mutable;Ch : GraphNode from PXCAFDoc)
    returns Integer from Standard;
    
    GetFather (me ; Findex : Integer from Standard)
    returns GraphNode from PXCAFDoc;
	
    GetChild (me ; Chindex : Integer from Standard)
    returns GraphNode from PXCAFDoc;
    
    FatherIndex (me ; F : GraphNode from PXCAFDoc)
    returns Integer from Standard;
    
    ChildIndex (me ; Ch : GraphNode from PXCAFDoc)
    returns Integer from Standard;

    NbFathers (me) returns Integer from Standard;

    NbChildren (me) returns Integer from Standard;

    SetGraphID(me : mutable; GUID : GUID from Standard);

    GetGraphID(me) returns GUID from Standard;

fields

	myFathers  : GraphNodeSequence from PXCAFDoc;
	myChildren : GraphNodeSequence from PXCAFDoc;
    	myGraphID  : GUID              from Standard;
	
end GraphNode;
