-- File:	GeomFill_DraftTrihedron.cdl
-- Created:	Tue Apr 14 09:48:24 1998
-- Author:	 Stephanie HUMEAU
--		<shu@sun17>
---Copyright:	 Matra Datavision 1998

----------------------------------------------------
-- Triedre de Frenet pour une surface de depouille
----------------------------------------------------

class  DraftTrihedron  from  GeomFill   
inherits  TrihedronLaw  from  GeomFill 

uses  
    Shape  from  GeomAbs, 
    Array1OfReal   from TColStd, 
    Vec  from  gp  

raises
    OutOfRange,  ConstructionError

is 
    Create (BiNormal :  Vec from gp;   
    	    Angle  :  Real )   
    returns  DraftTrihedron  from  GeomFill;  
     
    SetAngle(me  :  mutable; Angle  :  Real) 
    is  static; 

    Copy(me)  returns  TrihedronLaw  from  GeomFill          
     is  redefined;
     
  
    D0( me : mutable;  
        Param  : Real; 
        Tangent    : out  Vec  from  gp; 
        Normal     : out  Vec  from  gp;  
        BiNormal   : out  Vec  from  gp)        
    returns Boolean  is  redefined;    
      
  ---Purpose: compute Triedrhon and derivative Trihedron on curve at
  --          parameter <Param>
  --  Warning : It used  only for C1 or C2 aproximation
    D1( me : mutable;
        Param: Real;       
        Tangent    : out  Vec  from  gp;  
        DTangent   : out  Vec  from  gp; 
        Normal     : out  Vec  from  gp; 
        DNormal    : out  Vec  from  gp;                 
        BiNormal   : out  Vec  from  gp; 
        DBiNormal  : out  Vec  from  gp)
    returns Boolean  is  redefined; 

    ---Purpose: compute Trihedron on curve          
    --          first and seconde  derivatives.         
    --  Warning : It used only for C2 aproximation   
    D2( me : mutable;
        Param: Real;       
        Tangent    : out  Vec  from  gp;  
        DTangent   : out  Vec  from  gp; 
        D2Tangent  : out  Vec  from  gp; 
        Normal     : out  Vec  from  gp; 
        DNormal    : out  Vec  from  gp;                 
        D2Normal   : out  Vec  from  gp; 
        BiNormal   : out  Vec  from  gp; 
        DBiNormal  : out  Vec  from  gp; 
        D2BiNormal : out  Vec  from  gp)    
    returns Boolean  is  redefined;  

-- 
--  =================== Management  of  continuity  ===================
--                 
   NbIntervals(me; S : Shape from GeomAbs) 
	---Purpose: Returns  the number  of  intervals for  continuity
	--          <S>. 
        --          May be one if Continuity(me) >= <S>
   returns Integer  is  redefined;

   Intervals(me; T : in out Array1OfReal from TColStd; 
    	         S : Shape from GeomAbs)
	---Purpose: Stores in <T> the  parameters bounding the intervals
	--          of continuity <S>.
	--          
	--          The array must provide  enough room to  accomodate
	--          for the parameters. i.e. T.Length() > NbIntervals()
    raises
    	OutOfRange from Standard 
    is redefined;    
    
--  =====================  To help   computation of  Tolerance ============	 
    GetAverageLaw(me  :  mutable;
      ATangent    : out  Vec  from  gp; 
      ANormal     : out  Vec  from  gp; 
      ABiNormal   : out  Vec  from  gp) 
     ---Purpose: Get average value of Tangent(t) and Normal(t) it is usefull to 
     --          make fast approximation of rational  surfaces.        
  is  redefined; 
   
  
--   =================== To help Particular case   ===============	
   
    IsConstant(me) 
    ---Purpose: Say if the law is Constant.        
    returns  Boolean   
    is redefined;   
     
    IsOnlyBy3dCurve(me) 
     ---Purpose: Return True.        
    returns  Boolean   
    is redefined;   
     
fields  
 
    B :  Vec  from  gp; 
    myAngle  :  Real  from  Standard;  
    myCos    :  Real;
   
end  DraftTrihedron; 


