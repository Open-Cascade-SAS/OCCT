-- Created on: 1995-07-17
-- Created by: Laurent BUCHARD
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



generic class HCurve2dToolGen from BRepBlend (
     CurveGen  as any)

uses 
     Array1OfReal    from TColStd,
     Shape           from GeomAbs,
     CurveType       from GeomAbs,
     Vec2d             from gp,
     Pnt2d             from gp,
     Circ2d            from gp,
     Elips2d           from gp,
     Hypr2d            from gp,
     Parab2d           from gp,
     Lin2d             from gp,
     BezierCurve     from Geom2d,
     BSplineCurve    from Geom2d
     
raises
    
    OutOfRange          from Standard,
    NoSuchObject        from Standard,
    DomainError         from Standard
 
is

    --
    --     Global methods - Apply to the whole curve.
    --     
    
    FirstParameter(myclass; C: CurveGen) returns Real
    	---C++: inline
    ;
    

    LastParameter(myclass; C: CurveGen) returns Real
    	---C++: inline    
    ;

    --
    -- Services to break the curves to the expected continuity
    -- 
    --  If  for example you  need the  curve to  be C2  and the method
    --  Continuity   returns you something lower than   C2 (say C1 for
    --  example).
    --  
    --  First  compute the   number  of intervals  with  the requested
    --  continuity with the method  NbIntervals().   Note that if  the
    --  continuity  is higher than the one   you need NbIntervals will
    --  return 1.
    --  
    --  Then you get the parameters  bounding  the intervals with  the
    --  method  Intervals,   using   an array    of  length  at  least
    --  NbIntervals()+1.
    -- 
    -- If you need  to create a curve  with a restricted span you  can
    -- use the method Trim().

    
    Continuity(myclass; C: CurveGen) returns Shape from GeomAbs
	---Purpose: 
	---C++: inline
    ;
    
    NbIntervals(myclass; C: CurveGen; S : Shape from GeomAbs) returns Integer
	---Purpose: Returns  the number  of  intervals for  continuity
	--          <S>. May be one if Continuity(myclass) >= <S>
	---C++: inline
    ;
    
    Intervals(myclass; C: CurveGen; T : in out Array1OfReal from TColStd; 
    	          S : Shape from GeomAbs)
	---Purpose: Stores in <T> the  parameters bounding the intervals
	--          of continuity <S>.
	--          
	--          The array must provide  enough room to  accomodate
	--          for the parameters. i.e. T.Length() > NbIntervals()
    raises
    	OutOfRange from Standard
    ---C++: inline
    ;
    
    IsClosed(myclass; C: CurveGen) returns Boolean
    ---C++: inline    
    ;
     
    IsPeriodic(myclass; C: CurveGen) returns Boolean
    ---C++: inline
    ;
    
    Period(myclass; C: CurveGen) returns Real
    raises
    	DomainError from Standard -- if the curve is not periodic
    ---C++: inline	
    ;
     
    Value(myclass; C: CurveGen; U : Real) returns Pnt2d from gp
         --- Purpose : Computes the point of parameter U on the curve.
    ---C++: inline
    ;
    
    D0 (myclass; C: CurveGen; U : Real; P : out Pnt2d from gp)
         --- Purpose : Computes the point of parameter U on the curve.
    ---C++: inline
    ;
    
    D1 (myclass; C: CurveGen; U : Real; P : out Pnt2d from gp ; V : out Vec2d from gp)
         --- Purpose : Computes the point of parameter U on the curve with its
         --  first derivative.
     raises 
    	DomainError from Standard
        --- Purpose : Raised if the continuity of the current interval
        --  is not C1.
    ---C++: inline
    ;
    
    D2 (myclass; C: CurveGen; U : Real; P : out Pnt2d from gp; V1, V2 : out Vec2d from gp)
        --- Purpose :
        --  Returns the point P of parameter U, the first and second
        --  derivatives V1 and V2.
     raises 
    	DomainError from Standard
        --- Purpose : Raised if the continuity of the current interval
        --  is not C2.
    ---C++: inline
     ;

    D3 (myclass; C: CurveGen; U : Real; P : out Pnt2d from gp; V1, V2, V3 : out Vec2d from gp)
        --- Purpose :
        --  Returns the point P of parameter U, the first, the second 
        --  and the third derivative.
     raises 
    	DomainError from Standard
        --- Purpose : Raised if the continuity of the current interval
        --  is not C3.
    ---C++: inline
     ;
        
    DN (myclass; C: CurveGen; U : Real; N : Integer)   returns Vec2d from gp
        --- Purpose :
        --  The returned vector gives the value of the derivative for the 
        --  order of derivation N.
     raises  
    	DomainError from Standard,
        --- Purpose : Raised if the continuity of the current interval
        --  is not CN.
        OutOfRange from Standard
        --- Purpose : Raised if N < 1.            
    ---C++: inline
     ;

    Resolution(myclass; C: CurveGen; R3d : Real) returns Real
         ---Purpose :  Returns the parametric  resolution corresponding
         --         to the real space resolution <R3d>.
    ---C++: inline
    ;   
        
    GetType(myclass; C: CurveGen) returns CurveType from GeomAbs
	---Purpose: Returns  the  type of the   curve  in the  current
	--          interval :   Line,   Circle,   Ellipse, Hyperbola,
	--          Parabola, BezierCurve, BSplineCurve, OtherCurve.
    ---C++: inline
    ;

    --
    --     The following methods must  be called when GetType returned
    --     the corresponding type.
    --     

     Line(myclass; C: CurveGen) returns Lin2d from gp
     raises 
    	NoSuchObject from Standard
    ---C++: inline
     ;
     
     Circle(myclass; C: CurveGen) returns Circ2d from gp
     raises 
    	NoSuchObject from Standard
    ---C++: inline
     ;
     
     Ellipse(myclass; C: CurveGen) returns Elips2d from gp
     raises 
    	NoSuchObject from Standard
    ---C++: inline
     ;
     
     Hyperbola(myclass; C: CurveGen) returns  Hypr2d from gp
     raises 
    	NoSuchObject from Standard
    ---C++: inline
     ;
     
     Parabola(myclass; C: CurveGen) returns Parab2d from gp
     raises 
    	NoSuchObject from Standard
    ---C++: inline
     ;
     
     Bezier(myclass; C: CurveGen) returns BezierCurve from Geom2d
     raises 
    	NoSuchObject from Standard
    ---C++: inline
     ;
    
     BSpline(myclass; C: CurveGen) returns BSplineCurve from Geom2d
     raises 
    	NoSuchObject from Standard
    ---C++: inline
     ;

    



    NbSamples(myclass; C: CurveGen; U0,U1: Real from Standard) 
    returns Integer from Standard;

end HCurve2dToolGen;


