-- Created on: 2000-01-28
-- Created by: data exchange team
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class BasicMsgRegistrator from ShapeExtend inherits TShared from MMgt

    ---Purpose: Abstract class that can be used for attaching messages
    --          to the objects (e.g. shapes).
    --          It is used by ShapeHealing algorithms to attach a message
    --          describing encountered case (e.g. removing small edge from
    --          a wire).
    --
    --          The methods of this class are empty and redefined, for instance,
    --          in the classes for Data Exchange processors for attaching
    --          messages to interface file entities or CAS.CADE shapes.

uses

    Shape   from TopoDS,
    Msg     from Message,
    Gravity from Message
     
is

    Create returns mutable BasicMsgRegistrator from ShapeExtend;
    	---Purpose: Empty constructor.

    Send (me: mutable; object : Transient;
    	    	       message: Msg from Message;
    	    	       gravity: Gravity from Message) is virtual;
    	---Purpose: Sends a message to be attached to the object.
	--          Object can be of any type interpreted by redefined MsgRegistrator.

    Send (me: mutable; shape  : Shape from TopoDS;
    	    	       message: Msg from Message;
    	    	       gravity: Gravity from Message) is virtual;
    	---Purpose: Sends a message to be attached to the shape.

    Send (me: mutable; message: Msg from Message;
    	    	       gravity: Gravity from Message) is virtual;
    	---Purpose: Calls Send method with Null Transient.

end BasicMsgRegistrator;
