-- Created on: 1991-05-16
-- Created by: Isabelle GRIGNON
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class IntLinTorus from IntAna 

	---Purpose: Intersection between a line and a torus.

uses Lin          from gp,
     Torus        from gp,
     Pnt          from gp

raises NotDone    from StdFail,
       OutOfRange from Standard


is

    Create
    
    	returns IntLinTorus from IntAna;

    Create(L : Lin from gp; T : Torus from gp)
    
    	---Purpose: Creates the intersection between a line and a torus.

    	returns IntLinTorus from IntAna;


    Perform(me: in out; L : Lin from gp; T : Torus from gp)
    
    	---Purpose: Intersects a line and a torus.

    	is static;


    IsDone(me)
    
	---Purpose: Returns True if the computation was successful.
	--          
	---C++: inline

    	returns Boolean from Standard
	
	is static;


    NbPoints(me)
    
    	---Purpose: Returns the number of intersection points.
	--          
	---C++: inline

    	returns Integer from Standard
	
	raises NotDone     from StdFail
    	--     The exception NotDone is raised if IsDone returns False. 

	is static;


    Value(me; Index : Integer from Standard)
    
    	---Purpose: Returns the intersection point of range Index.
	--          
	---C++: inline
	---C++: return const&

    	returns Pnt from gp

    	raises NotDone    from StdFail,
               OutOfRange from Standard
    	--     The exception NotDone is raised if IsDone returns False. 
    	--     The exception OutOfRange is raised if Index <= 0 or
    	--        Index > NbPoints
	
	is static;


    ParamOnLine(me; Index : Integer from Standard)
    
    	---Purpose: Returns the parameter on the line of the intersection
    	--          point of range Index.
	--          
	---C++: inline

    	returns Real from Standard

    	raises NotDone    from StdFail,
               OutOfRange from Standard
    	--     The exception NotDone is raised if IsDone returns False. 
    	--     The exception OutOfRange is raised if Index <= 0 or
    	--        Index > NbPoints
	
	is static;


    ParamOnTorus(me; Index : Integer from Standard;
                     FI,THETA: out Real from Standard)
    
    	---Purpose: Returns the parameters on the torus of the intersection
    	--          point of range Index.
	--          
	---C++: inline

    	raises NotDone    from StdFail,
               OutOfRange from Standard
    	--     The exception NotDone is raised if IsDone returns False. 
    	--     The exception OutOfRange is raised if Index <= 0 or
    	--        Index > NbPoints
	
	is static;


fields

    done    : Boolean      from Standard;
    nbpt    : Integer      from Standard;
    thePoint: Pnt          from gp [4];
    theParam: Real         from Standard [4];
    theFi   : Real         from Standard [4];
    theTheta: Real         from Standard [4];

end IntLinTorus;
