-- Created on: 1999-11-26
-- Created by: Andrey BETENEV
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0

class ProductCategoryRelationship from StepBasic
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity ProductCategoryRelationship

uses
    HAsciiString from TCollection,
    ProductCategory from StepBasic

is
    Create returns ProductCategoryRelationship from StepBasic;
	---Purpose: Empty constructor

    Init (me: mutable; aName: HAsciiString from TCollection;
                       hasDescription: Boolean;
                       aDescription: HAsciiString from TCollection;
                       aCategory: ProductCategory from StepBasic;
                       aSubCategory: ProductCategory from StepBasic);
	---Purpose: Initialize all fields (own and inherited)

    Name (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Name
    SetName (me: mutable; Name: HAsciiString from TCollection);
	---Purpose: Set field Name

    Description (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Description
    SetDescription (me: mutable; Description: HAsciiString from TCollection);
	---Purpose: Set field Description
    HasDescription (me) returns Boolean;
	---Purpose: Returns True if optional field Description is defined

    Category (me) returns ProductCategory from StepBasic;
	---Purpose: Returns field Category
    SetCategory (me: mutable; Category: ProductCategory from StepBasic);
	---Purpose: Set field Category

    SubCategory (me) returns ProductCategory from StepBasic;
	---Purpose: Returns field SubCategory
    SetSubCategory (me: mutable; SubCategory: ProductCategory from StepBasic);
	---Purpose: Set field SubCategory

fields
    theName: HAsciiString from TCollection;
    theDescription: HAsciiString from TCollection; -- optional
    theCategory: ProductCategory from StepBasic;
    theSubCategory: ProductCategory from StepBasic;
    defDescription: Boolean; -- flag "is Description defined"

end ProductCategoryRelationship;
