-- Created on: 1992-09-28
-- Created by: Remi GILET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MakeMirror

from GC

    ---Purpose: This class implements elementary construction algorithms for a
    -- symmetrical transformation in 3D space about a point,
    -- axis or plane. The result is a Geom_Transformation transformation.
    -- A MakeMirror object provides a framework for:
    -- -   defining the construction of the transformation,
    -- -   implementing the construction algorithm, and
    -- -   consulting the result.

uses Pnt            from gp,
     Ax1            from gp,
     Ax2            from gp,
     Dir            from gp,
     Pln            from gp,
     Lin            from gp,
     Transformation from Geom,
     Real           from Standard
     
is

Create(Point : Pnt from gp) returns MakeMirror;
    ---Puprose: Make a symetry transformation of center <Point>.

Create(Axis : Ax1 from gp) returns MakeMirror;
    ---Puprose: Make a symetry transformation of axis <Axis>.

Create(Line : Lin from gp) returns MakeMirror;
    ---Puprose: Make a symetry transformation of axis <Line>.

Create(Point : Pnt from gp;
       Direc : Dir from gp) returns MakeMirror;
    ---Purpose: Make a symetry transformation af axis defined by 
    --          <Point> and <Direc>.

Create(Plane : Pln from gp) returns MakeMirror;
    ---Purpose: Make a symetry transformation of plane <Plane>.

Create(Plane : Ax2 from gp) returns MakeMirror;
    ---Purpose: Make a symetry transformation of plane <Plane>.

Value(me) returns Transformation from Geom
    is static;
    ---Purpose: Returns the constructed transformation.
    ---C++: return const&
    ---C++: alias "operator const Handle(Geom_Transformation)& () const { return Value(); }"

fields

    TheMirror : Transformation from Geom;

end MakeMirror;

