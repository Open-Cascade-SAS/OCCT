-- Created on: 2001-07-25
-- Created by: Julia DOROVSKIKH
-- Copyright (c) 2001-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class DocumentRetrievalDriver from XmlLDrivers inherits RetrievalDriver from PCDM

uses
    ExtendedString		from TCollection,
    SequenceOfExtendedString	from TColStd,
    Document			from PCDM,
    Document			from CDM,
    Document			from TDocStd,
    Application			from CDM,
    ADriver		        from XmlMDF, 
    ADriverTable		from XmlMDF,
    RRelocationTable		from XmlObjMgt,
    Element			from XmlObjMgt,
    MessageDriver               from CDM

is
    Create returns mutable DocumentRetrievalDriver from XmlLDrivers;
    -- Constructor

    SchemaName		(me)
	returns ExtendedString from TCollection is redefined virtual;
    -- pure virtual method definition

    Make		(me : mutable; PD : Document from PCDM;
				       TD : Document from CDM)
	is redefined virtual;
    -- pure virtual method definition

    CreateDocument	(me : mutable)
	returns Document from CDM is redefined virtual;
    -- pure virtual method definition

    Read(me:mutable; theFileName:    ExtendedString from TCollection;
    	    	     theNewDocument: Document    from CDM;
    	    	     theApplication: Application from CDM) is redefined virtual;
    -- 

    ReadFromDomDocument (me : mutable; theDomElement: Element from XmlObjMgt;
				       theNewDocument: Document from CDM;
				       theApplication: Application from CDM)
	is virtual protected;

    MakeDocument	(me : mutable; thePDoc: Element  from XmlObjMgt;
    	    	    	       theTDoc: Document from CDM)
    	returns Boolean from Standard
	is virtual protected;

    AttributeDrivers	(me : mutable; theMsgDriver: MessageDriver from CDM)
	returns ADriverTable from XmlMDF
	is virtual; 
	
    ReadShapeSection (me:mutable; thePDoc  :  Element from XmlObjMgt; 
    	    	    	    	  theMsgDriver : MessageDriver from CDM) 
        returns ADriver from XmlMDF
        is virtual protected; 
	 
    ShapeSetCleaning(me:mutable; theDriver : ADriver from XmlMDF) 
        is virtual protected;  
	
    PropagateDocumentVersion(me:mutable; theDocVersion : Integer from Standard) 
        is virtual protected; 
	
fields
    myDrivers	: ADriverTable		from XmlMDF      is protected;
    myRelocTable: RRelocationTable	from XmlObjMgt   is protected;
    myFileName  : ExtendedString        from TCollection is protected;

end DocumentRetrievalDriver;
