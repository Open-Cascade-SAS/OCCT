-- Created on: 1999-05-21
-- Created by: Pavel DURANDIN
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ConvertSurfaceToBezierBasis from ShapeUpgrade inherits SplitSurface from ShapeUpgrade

	---Purpose: Converts a plane, bspline surface, surface of revolution, surface 
    	--          of extrusion, offset surface to grid of bezier basis surface (
	--           bezier surface,
	--           surface of revolution based on bezier curve,
	--           offset surface based on any previous type).

uses

    CompositeSurface from ShapeExtend

is

    Create returns mutable ConvertSurfaceToBezierBasis from ShapeUpgrade;
    	---Purpose: Empty constructor.
    
    Build (me: mutable; Segment: Boolean) is redefined;
    	---Purpose: Splits a list of beziers computed by Compute method according
	--          the split values and splitting parameters.
    
    Compute(me: mutable; Segment: Boolean) is redefined;
    	---Purpose: Converts surface into a grid of bezier based surfaces, and
	--          stores this grid.
    
    Segments(me) returns CompositeSurface from ShapeExtend;
    	---Purpose: Returns the grid of bezier based surfaces correspondent to 
        --          original surface.
    
    --Methods for handling surface modes

    SetPlaneMode(me: mutable; mode: Boolean);
    	---Purpose: Sets mode for conversion Geom_Plane to Bezier
	---C++: inline
    
    GetPlaneMode(me) returns Boolean;
    	---Purpose: Returns the Geom_Pline conversion mode.
    	---C++: inline
    
    SetRevolutionMode(me: mutable; mode: Boolean);
    	---Purpose: Sets mode for conversion Geom_SurfaceOfRevolution to Bezier
	---C++: inline
    
    GetRevolutionMode(me) returns Boolean;
    	---Purpose: Returns the Geom_SurfaceOfRevolution conversion mode.
    	---C++: inline
    
    SetExtrusionMode(me: mutable; mode: Boolean);
    	---Purpose: Sets mode for conversion Geom_SurfaceOfLinearExtrusion to Bezier
	---C++: inline
    
    GetExtrusionMode(me) returns Boolean;
    	---Purpose: Returns the Geom_SurfaceOfLinearExtrusion conversion mode.
    	---C++: inline
    
    SetBSplineMode(me: mutable; mode: Boolean);
    	---Purpose: Sets mode for conversion Geom_BSplineSurface to Bezier
	---C++: inline
    
    GetBSplineMode(me) returns Boolean;
    	---Purpose: Returns the Geom_BSplineSurface conversion mode.
    	---C++: inline
    
fields

    mySegments      : CompositeSurface from ShapeExtend;
    myPlaneMode     : Boolean;
    myRevolutionMode: Boolean;
    myExtrusionMode : Boolean;
    myBSplineMode   : Boolean;
    
end ConvertSurfaceToBezierBasis;
