-- Created on: 1999-01-14
-- Created by: Xuan PHAM PHU
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class face from TopOpeBRepTool

uses
    Wire from TopoDS,
    Face from TopoDS
is
    Create returns face from TopOpeBRepTool;
    Init (me : in out; W : Wire from TopoDS; Fref : Face from TopoDS) 
    returns Boolean;
    -- Builds face f for <myW> on <Fref>, 
    -- updates <myfinite> to true if f is finite,
    -- <myFfinite> is finite.
    -- returns false if the compute fails
    W(me) returns Wire from TopoDS;
    ---C++: return const &
    
    IsDone(me)  returns Boolean;    
    
    Finite(me)  returns Boolean;    
    Ffinite(me) returns Face from TopoDS; 
    ---C++: return const &   
    RealF(me)   returns Face from TopoDS;
    -- Raises if !IsDone
    
fields
    myW       : Wire from TopoDS;
    myfinite  : Boolean;
    myFfinite : Face from TopoDS;
    
end face;
