-- Created on: 2001-09-11
-- Created by: Julia DOROVSKIKH
-- Copyright (c) 2001-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class LocationDriver from XmlMXCAFDoc  inherits ADriver from XmlMDF



        ---Purpose: Attribute Driver.

uses    Location         from TopLoc,
        Element          from XmlObjMgt,
        SRelocationTable from XmlObjMgt,
        RRelocationTable from XmlObjMgt,
        Persistent       from XmlObjMgt,
        MessageDriver    from CDM,
        Attribute        from TDF,
        LocationSetPtr   from TopTools

is
    Create (theMessageDriver:MessageDriver from CDM)
        returns mutable LocationDriver from XmlMXCAFDoc;



    NewEmpty (me)  returns mutable Attribute from TDF;




    Paste(me; Source     : Persistent from XmlObjMgt;
              Target     : mutable Attribute from TDF;
              RelocTable : out RRelocationTable from XmlObjMgt)
        returns Boolean from Standard;

    Paste(me; Source     : Attribute from TDF;
              Target     : in out Persistent from XmlObjMgt;
              RelocTable : out SRelocationTable from XmlObjMgt);

    Translate (me; theLoc    : Location from TopLoc;
                        theParent : in out Element from XmlObjMgt;
                        theMap    : in out SRelocationTable from XmlObjMgt);
        ---Purpose: Translate a non storable Location to a storable Location.
        ---Level: Internal

    Translate (me; theParent : Element from XmlObjMgt;
                        theLoc    : in out Location from TopLoc;
                        theMap    : in out RRelocationTable from XmlObjMgt)
    returns Boolean from Standard;
        ---Purpose: Translate a storable Location to a non storable Location.
        ---Level: Internal

    SetSharedLocations(me: mutable;
                       theLocations:  in LocationSetPtr  from TopTools);
    ---C++: inline

fields
    myLocations : LocationSetPtr   from TopTools;
end LocationDriver;
