-- Created on: 1992-09-29
-- Created by: Remi GILET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


private deferred class Root from gce 

    ---Purpose : This class implements the common services for
    --           all classes of gce which report error.

uses 

ErrorType from gce

is

    IsDone(me) returns Boolean
    	is static;
    ---C++: inline
    ---Purpose: Returns true if the construction is successful.
    
    Status(me) returns ErrorType from gce
    	is static;
    ---C++: inline
    ---Purpose:
    -- Returns the status of the construction:
    -- -   gce_Done, if the construction is successful, or
    -- -   another value of the gce_ErrorType enumeration
    --   indicating why the construction failed.

fields

    TheError     : ErrorType from gce is protected;
    ---Purpose: Enumeration to know why the algorithm didn t succeed.

end Root;

