-- Created on: 1997-11-28
-- Created by: Robert COUBLANC
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ExclusionFilter from AIS inherits Filter from SelectMgr

    	---Purpose:  A framework to reject or to accept only objects of
    	-- given types and/or signatures.
    	-- Objects are stored, and the stored objects - along
    	-- with the flag settings - are used to define the filter.
    	-- Objects to be filtered are compared with the stored
    	-- objects added to the filter, and are accepted or
    	-- rejected according to the exclusion flag setting.
    	-- -   Exclusion flag on
    	--   -   the function IsOk answers true for all objects,
    	--    except those of the types and signatures stored
    	--    in the filter framework
    	-- -   Exclusion flag off
    	--   -   the funciton IsOk answers true for all objects
    	--    which have the same type and signature as the stored ones.

uses
    
     EntityOwner from SelectMgr,
     KindOfInteractive from AIS,
     ListOfInteger from TColStd,
     DataMapOfIntegerListOfInteger from TColStd
is
    
    Create(ExclusionFlagOn:Boolean from Standard = Standard_True)
    returns mutable ExclusionFilter from AIS;
    	---Purpose: Constructs an empty exclusion filter object defined by
    	-- the flag setting ExclusionFlagOn.
    	-- By default, the flag is set to true.
    
    Create(TypeToExclude : KindOfInteractive from AIS;
	   ExclusionFlagOn : Boolean from Standard = Standard_True)
    returns  mutable ExclusionFilter from AIS;
    	---Purpose: All the AIS objects of <TypeToExclude>
    	--          Will be rejected by the IsOk Method.
    
    
    Create(TypeToExclude : KindOfInteractive from AIS;
    	   SignatureInType :Integer from Standard ;
	   ExclusionFlagOn : Boolean from Standard = Standard_True)
    returns  mutable ExclusionFilter from AIS;
    	---Purpose: Constructs an exclusion filter object defined by the
    	-- enumeration value TypeToExclude, the signature
    	-- SignatureInType, and the flag setting ExclusionFlagOn.
    	-- By default, the flag is set to true.
    

    IsOk(me; anObj : EntityOwner from SelectMgr)
    returns Boolean from Standard
    is redefined virtual;





	    ---Category: Load Filter...

    Add(me:mutable;TypeToExclude : KindOfInteractive from AIS) 
    returns Boolean from Standard;
   	---Purpose: Adds the type TypeToExclude to the list of types.

    Add(me:mutable;
    	TypeToExclude   : KindOfInteractive from AIS;
        SignatureInType : Integer from Standard) 
    returns Boolean from Standard;
	
    Remove(me:mutable;
    	   TypeToExclude:KindOfInteractive from AIS)
    returns Boolean from Standard;

    Remove(me:mutable;
    	   TypeToExclude:KindOfInteractive from AIS;
           SignatureInType : Integer from Standard) 
    returns Boolean from Standard;

    Clear(me:mutable);

	    ---Category: Information about Filter...



    IsExclusionFlagOn(me) returns Boolean from Standard;
    	---C++: inline

    SetExclusionFlag(me:mutable; Status : Boolean from Standard);
    	---C++: inline


    IsStored(me;aType:KindOfInteractive from AIS) returns Boolean from Standard;
    
    ListOfStoredTypes( me; TheList: in out ListOfInteger from TColStd);
    
    ListOfSignature(me;
    	    	    aType         : KindOfInteractive from AIS;
    	    	    TheStoredList : in out ListOfInteger from TColStd);
		

    IsSignatureIn(me;aType:KindOfInteractive from AIS;aSignature:Integer from Standard)
    returns Boolean from Standard is static private;

fields
    myIsExclusionFlagOn : Boolean from Standard;
    myStoredTypes       : DataMapOfIntegerListOfInteger from TColStd;
end ExclusionFilter;
