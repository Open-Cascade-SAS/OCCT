-- Created on: 1994-05-31
-- Created by: Christian CAILLET
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class SelectVisibleStatus  from IGESSelect  inherits SelectExtract

    ---Purpose : This selection looks at Blank Status of IGES Entities
    --           Direct  selection keeps Visible Entities (Blank = 0),
    --           Reverse selection keeps Blanked Entities (Blank = 1)


uses AsciiString from TCollection, Transient, InterfaceModel

is

    Create returns mutable SelectVisibleStatus;
    ---Purpose : Creates a SelectVisibleStatus

    Sort (me; rank : Integer; ent : Transient; model : InterfaceModel)
    	returns Boolean;
    ---Purpose : Returns True if <ent> is an IGES Entity with Blank Status = 0

    ExtractLabel (me) returns AsciiString from TCollection;
    ---Purpose : Returns the Selection criterium : "IGES Entity, Status Visible"

end SelectVisibleStatus;
