-- Created on: 1995-01-09
-- Created by: Modelistation
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Wedge from BRepPrim inherits GWedge from BRepPrim

	---Purpose: Provides constructors without Builders.

uses
    Ax2 from gp,
    Pnt from gp

raises
    DomainError

is

    Create(Axes : Ax2 from gp; dx, dy, dz : Real)
    returns Wedge from BRepPrim
	---Purpose: Creates a  Wedge  algorithm.   <Axes> is  the axis
	--          system for the primitive.
	--          
	--          XMin, YMin, ZMin are set to 0
	--          XMax, YMax, ZMax are set to dx, dy, dz
	--          Z2Min = ZMin
	--          Z2Max = ZMax
	--          X2Min = XMin
	--          X2Max = XMax
	--          The result is a box
	--          dx,dy,dz should be positive
	raises DomainError;

    Create(Axes : Ax2 from gp; dx, dy, dz, ltx : Real)
    returns Wedge from BRepPrim
	---Purpose: Creates  a Wedge  primitive. <Axes> is   the  axis
	--          system for the primitive.
	--          
	--          XMin, YMin, ZMin are set to 0
	--          XMax, YMax, ZMax are set to dx, dy, dz
	--          Z2Min = ZMin
	--          Z2Max = ZMax
	--          X2Min = ltx
	--          X2Max = ltx
	--          The result is a STEP right angular wedge
	--          dx,dy,dz should be positive
	--          ltx should not be negative
	raises DomainError;

    Create(Axes : Ax2 from gp; xmin, ymin, zmin, z2min, x2min,
                                   xmax, ymax, zmax, z2max, x2max : Real)
    returns Wedge from BRepPrim
	---Purpose: Create  a Wedge primitive.   <Axes>  is  the  axis
	--          system for the primitive.
	--          
	--          all the fields are set to the corresponding value
	--          XYZMax - XYZMin should be positive
	--          ZX2Max - ZX2Min should not be negative 
	raises DomainError;

end Wedge;
