-- Created by: TCL
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


deferred class Tolerance from Prs2d inherits Line from Graphic2d

	---Purpose: Groups all the tolerances
	
uses

	GraphicObject from Graphic2d,
	Drawer        from Graphic2d,
	Length	      from Quantity

is
	
	Initialize( aGO                    : GraphicObject from Graphic2d;
		        aX, aY                 : Real          from Standard;
			    aLength                : Real          from Standard;
                anAngle                : Real          from Standard );
	---Level: Public
	---Purpose: Creates a tolerance with the center in the point (<aX>, <aY>); 
	--          reference point is <aXPosition>, <aYPosition>
	---Category: Constructor

    SetCoord( me: mutable; aX, aY: Real from Standard );
    ---Level: Public
    ---Purpose: Changes the coordinates of this tolerance

    SetSize( me: mutable; aLen: Real from Standard );
    ---Level: Public
    ---Purpose: Defines the size of this one

    Pick( me : mutable; X, Y: ShortReal from Standard;
		  aPrecision: ShortReal from Standard;
		  aDrawer: Drawer from Graphic2d )
	returns Boolean from Standard is protected;
	---Level: Internal
	---Purpose: Returns Standard_True if the Tolerance is picked,
	--	        Standard_False if not.


fields

   myX      : ShortReal from Standard is protected;
   myY      : ShortReal from Standard is protected;
   myLength : ShortReal from Standard is protected;
   myAngle  : ShortReal from Standard is protected;

friends

   class ToleranceFrame from Prs2d
    
end Tolerance from Prs2d;
