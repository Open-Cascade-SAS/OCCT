-- Created on: 1992-08-18
-- Created by: Arnaud BOUZY
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class GenFct from ExprIntrp inherits Generator from ExprIntrp

	---Purpose: Implements an interpreter for defining functions. 
	--          All its functionnalities can be found in class 
	--          GenExp. 

uses NamedFunction from Expr,
    SequenceOfNamedFunction from ExprIntrp,
    AsciiString from TCollection

raises NoSuchObject

is

    Create
    ---Level: Internal 
    returns mutable GenFct is private;

    Create( myclass ) returns GenFct;
        
    Process(me : mutable; str : AsciiString)
    ---Level: Internal 
    is static;

    IsDone(me)
    ---Level: Internal 
    returns Boolean
    is static;
	    
fields

    done : Boolean;
    
end GenFct;
