-- Created on: 1993-12-24
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class S from Law inherits BSpFunc from Law

	---Purpose: Describes an "S" evolution law. 

is

    Create
    returns S from Law;

    	---Purpose: Constructs an empty "S" evolution law.
    Set(me: mutable; Pdeb,Valdeb,Pfin,Valfin: Real from Standard)
    is static;
    	---Purpose:
    	-- Defines this S evolution law by assigning both:
    	-- -   the bounds Pdeb and Pfin of the parameter, and
    	-- -   the values Valdeb and Valfin of the function at these
    	--   two parametric bounds.
    	-- The function is assumed to have the first derivatives
    	-- equal to 0 at the two parameter points Pdeb and Pfin.

    Set(me: mutable; Pdeb,Valdeb,Ddeb,Pfin,Valfin,Dfin: Real from Standard)
    is static;
    	---Purpose: Defines this S evolution law by assigning
    	-- -   the bounds Pdeb and Pfin of the parameter,
    	-- -   the values Valdeb and Valfin of the function at these
    	--   two parametric bounds, and
	-- -   the values Ddeb and Dfin of the first derivative of the
    	--   function at these two parametric bounds.

end S;
