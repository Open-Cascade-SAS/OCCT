-- File:	RWStepAP214_RWAppliedPersonAndOrganizationAssignment.cdl
-- Created:	Fri Mar 12 14:32:39 1999
-- Author:	data exchange team
--		<det@androx.nnov.matra-dtv.fr>
---Copyright:	 Matra Datavision 1999


class RWAppliedPersonAndOrganizationAssignment from RWStepAP214 

	---Purpose: Read & Write Module for AppliedPersonAndOrganizationAssignment

uses
     Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     AppliedPersonAndOrganizationAssignment from StepAP214,
     EntityIterator from Interface

is
    	Create returns RWAppliedPersonAndOrganizationAssignment;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable AppliedPersonAndOrganizationAssignment from StepAP214);

	WriteStep (me; SW : in out StepWriter; ent : AppliedPersonAndOrganizationAssignment from StepAP214);

	Share(me; ent : AppliedPersonAndOrganizationAssignment from StepAP214; iter : in out EntityIterator);



end RWAppliedPersonAndOrganizationAssignment;
