-- Created on: 1995-03-16
-- Created by: Christian CAILLET
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class FuncShape  from XSControl

    ---Purpose : Defines additionnal commands for XSControl to :
    --           - control of initialisation (xinit, xnorm, newmodel)
    --           - analyse of the result of a transfer (recorded in a
    --             TransientProcess for Read, FinderProcess for Write) :
    --             statistics, various lists (roots,complete,abnormal), what
    --             about one specific entity, producing a model with the
    --             abnormal result
    --             
    --           This appendix of XSControl is compiled separately to distinguish
    --           basic features from user callable forms

uses CString, AsciiString from TCollection,
     WorkSession from XSControl, HSequenceOfShape from TopTools

is

    Init (myclass);
    ---Purpose : Defines and loads all functions which work on shapes for XSControl (as ActFunc)

    MoreShapes (myclass; session : WorkSession from XSControl;
    	    	list : in out mutable HSequenceOfShape from TopTools;
                name : CString) returns Integer;
    ---Purpose : Analyses a name as designating Shapes from a Vars or from
    --           XSTEP transfer (last Transfer on Reading). <name> can be :
    --           "*" : all the root shapes produced by last Transfer (Read)
    --                 i.e. considers roots of the TransientProcess
    --           a name : a name of a variable DRAW
    --           
    --           Returns the count of designated Shapes. Their list is put in
    --           <list>. If <list> is null, it is firstly created. Then it is
    --           completed (Append without Clear) by the Shapes found
    --           Returns 0 if no Shape could be found

    FileAndVar (myclass; session : WorkSession from XSControl;
    	    	file, var, def : CString;
                 resfile, resvar : out AsciiString from TCollection)
        returns Boolean;
    ---Purpose : Analyses given file name and variable name, with a default
    --           name for variables. Returns resulting file name and variable
    --           name plus status "file to read"(True) or "already read"(False)
    --           In the latter case, empty resfile means no file available
    --           
    --           If <file> is null or empty or equates ".", considers Session
    --             and returned status is False
    --           Else, returns resfile = file and status is True
    --           If <var> is neither null nor empty, resvar = var
    --           Else, the root part of <resfile> is considered, if defined
    --           Else, <def> is taken


end FuncShape;
