-- Created on: 1994-03-28
-- Created by: Remi LEQUETTE
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class Point from DrawTrSurf inherits Drawable3D from Draw

	---Purpose: A drawable point.

uses
    	Pnt from gp,
    	Pnt2d from gp,
	MarkerShape from Draw,
     	Color from Draw,
     	Display from Draw,
     	Drawable3D from Draw,
	Interpretor from Draw

is

    Create( P : Pnt from gp; 
    	    Shape : MarkerShape from Draw;
	    Col   : Color from Draw) 
    returns mutable Point from DrawTrSurf;
    
    Create( P : Pnt2d from gp; 
    	    Shape : MarkerShape from Draw;
	    Col   : Color from Draw) 
    returns mutable Point from DrawTrSurf;
    
    DrawOn (me; dis : in out Display from Draw);
     
    Is3D(me) returns Boolean
	---Purpose: Is a 3D object. (Default True).
    is redefined;
    
    Point(me) returns Pnt from gp
    is static;
    
    Point(me : mutable; P : Pnt from gp)
    is static;

    Point2d(me) returns Pnt2d from gp
    is static;
    
    Point2d(me : mutable; P : Pnt2d from gp)
    is static;

  Color(me : mutable; aColor : Color from Draw)
     is static;

  Color (me)  returns Color from Draw
     is static;
     
  Shape(me : mutable; S : MarkerShape from Draw)
  is static;
  
  Shape(me) returns MarkerShape from Draw
  is  static;
     
  Copy(me) returns mutable Drawable3D from Draw
	---Purpose: For variable copy.
  is redefined;
  
  Dump(me; S : in out OStream)
	---Purpose: For variable dump.
  is redefined;

  Whatis(me; I : in out Interpretor from Draw)
	---Purpose: For variable whatis command.
  is redefined;

fields

    myPoint : Pnt from gp;
    is3D    : Boolean;
    myShape : MarkerShape from Draw;
    myColor : Color from Draw;

end Point;


