-- Created on: 2013-02-05
-- Created by: Julia GERASIMOVA
-- Copyright (c) 2001-2013 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DiscreteTrihedron from GeomFill
    inherits TrihedronLaw  from  GeomFill 
    
       	---Purpose: Defined Discrete Trihedron Law.        
       	--          The requirement for path curve is only G1.
       	--          The result is C0-continuous surface
       	--          that can be later approximated to C1.

uses
    HCurve from  Adaptor3d, 
    Shape  from  GeomAbs, 
    Pnt    from  gp,
    Vec    from  gp,
    Array1OfReal from TColStd,
    Frenet from GeomFill,
    HSequenceOfAx2 from GeomFill,
    HSequenceOfReal from TColStd

raises
 OutOfRange,  ConstructionError
is  

   Create  
      returns DiscreteTrihedron from GeomFill 
      raises  ConstructionError; 
    
   Copy(me)   
   returns  TrihedronLaw  from  GeomFill          
   is  redefined;
 
   Init(me: mutable)   
   is  static; 

   SetCurve(me : mutable;  C  :  HCurve  from  Adaptor3d) 
   is  redefined;

-- 
-- 
--========== To compute Location and derivatives Location
--              
   D0(me : mutable; 
      Param: Real; 
      Tangent    : out  Vec  from  gp; 
      Normal     : out  Vec  from  gp; 
      BiNormal   : out  Vec  from  gp)
      ---Purpose: compute Trihedron on curve at parameter <Param>         
   returns Boolean  is  redefined;
	
   D1(me : mutable;
      Param: Real;       
      Tangent    : out  Vec  from  gp;  
      DTangent   : out  Vec  from  gp; 
      Normal     : out  Vec  from  gp; 
      DNormal    : out  Vec  from  gp;                 
      BiNormal   : out  Vec  from  gp; 
      DBiNormal  : out  Vec  from  gp)
      ---Purpose: compute Trihedron and  derivative Trihedron  on curve
      --          at parameter <Param>                
      --  Warning : It used only for C1 or C2 aproximation
      --  For the moment it returns null values for DTangent, DNormal
      --  and DBiNormal.
   returns Boolean  
   is  redefined; 
   
   D2(me : mutable;
      Param: Real;       
      Tangent    : out  Vec  from  gp;  
      DTangent   : out  Vec  from  gp; 
      D2Tangent  : out  Vec  from  gp; 
      Normal     : out  Vec  from  gp; 
      DNormal    : out  Vec  from  gp;                 
      D2Normal   : out  Vec  from  gp; 
      BiNormal   : out  Vec  from  gp; 
      DBiNormal  : out  Vec  from  gp; 
      D2BiNormal : out  Vec  from  gp)    
      ---Purpose: compute  Trihedron on curve          
      --          first and seconde  derivatives.
      --  Warning : It used only for C2 aproximation
      --  For the moment it returns null values for DTangent, DNormal
      --  DBiNormal, D2Tangent, D2Normal, D2BiNormal.
   returns Boolean
   is  redefined; 
--
--  =================== Management  of  continuity  ===================
--                 
   NbIntervals(me; S : Shape from GeomAbs) 
	---Purpose: Returns  the number  of  intervals for  continuity
	--          <S>. 
        --          May be one if Continuity(me) >= <S>
   returns Integer  is  redefined;

   Intervals(me; T : in out Array1OfReal from TColStd; 
    	         S : Shape from GeomAbs)
	---Purpose: Stores in <T> the  parameters bounding the intervals
	--          of continuity <S>.
	--          
	--          The array must provide  enough room to  accomodate
	--          for the parameters. i.e. T.Length() > NbIntervals()
    raises
    	OutOfRange from Standard 
    is redefined;  
     
	  
--  ===================  To help   computation of  Tolerance   ===============	 
    GetAverageLaw(me  :  mutable;
      ATangent    : out  Vec  from  gp; 
      ANormal     : out  Vec  from  gp; 
      ABiNormal   : out  Vec  from  gp) 
     ---Purpose: Get average value of Tangent(t) and Normal(t) it is usful to 
     --          make fast approximation of rational  surfaces.        
  is  redefined;

--   =================== To help Particular case   ===============	
   
    IsConstant(me) 
    ---Purpose: Say if the law is Constant.        
    returns  Boolean   
    is redefined;
 
   IsOnlyBy3dCurve(me) 
     ---Purpose: Return True.        
    returns  Boolean   
    is redefined;  
    

fields 

   myPoint      : Pnt  from  gp;
   myTrihedrons : HSequenceOfAx2  from GeomFill;
   myKnots      : HSequenceOfReal from TColStd;
   myFrenet     : Frenet  from GeomFill;
   myUseFrenet  : Boolean from Standard;
   
end DiscreteTrihedron;
