-- Created on: 1997-03-16
-- Created by: SMO
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package TPrsStd 

	---Purpose: The visualization attribute implements the
    	-- Application Interactive Services in the context
    	-- of Open CASCADE Application Framework.


    ---Category: GUID 
    --           04fb4d05-5690-11d1-8940-080009dc3333   TPrsStd_AISViewer
    --           04fb4d00-5690-11d1-8940-080009dc3333	TPrsStd_AISPresentation
   
uses
    Standard,
    TCollection,
    TColStd,
    MMgt,
    Quantity,
    Graphic3d,
    AIS,
    V3d,    
    TDF,
    TDataXtd,
    Geom,
    TopoDS,
    gp
    
    
is


    ---Category: Attributes 
    --           ==========
    
    class AISViewer;
    
    class AISPresentation;  

    ---Category : Drivers to build and/or update AIS objects
    --            ==========================================

    deferred class Driver;
      class PointDriver ;         -- to display Point
      class AxisDriver ;          -- to display Axis
      class PlaneDriver ;         -- to display Plane
      class GeometryDriver;       -- to display Geometry
      class ConstraintDriver;     -- to display Constraint
      class NamedShapeDriver;     -- to display NamedShape
    
    class DriverTable ;               
    
    ---Category: Tools
    --           =====

    class ConstraintTools;

    class DataMapOfGUIDDriver
    instantiates DataMap from TCollection(GUID      from Standard, 
	    	 		       	  Driver from TPrsStd, 
				          GUID      from Standard); 
end TPrsStd;

