-- Created on: 2003-01-22
-- Created by: data exchange team
-- Copyright (c) 2003-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class CurveElementIntervalLinearlyVarying from StepFEA
inherits CurveElementInterval from StepFEA

    ---Purpose: Representation of STEP entity CurveElementIntervalLinearlyVarying

uses
    CurveElementLocation from StepFEA,
    EulerAngles from StepBasic,
    HArray1OfCurveElementSectionDefinition from StepElement

is
    Create returns CurveElementIntervalLinearlyVarying from StepFEA;
	---Purpose: Empty constructor

    Init (me: mutable; aCurveElementInterval_FinishPosition: CurveElementLocation from StepFEA;
                       aCurveElementInterval_EuAngles: EulerAngles from StepBasic;
                       aSections: HArray1OfCurveElementSectionDefinition from StepElement);
	---Purpose: Initialize all fields (own and inherited)

    Sections (me) returns HArray1OfCurveElementSectionDefinition from StepElement;
	---Purpose: Returns field Sections
    SetSections (me: mutable; Sections: HArray1OfCurveElementSectionDefinition from StepElement);
	---Purpose: Set field Sections

fields
    theSections: HArray1OfCurveElementSectionDefinition from StepElement;

end CurveElementIntervalLinearlyVarying;
