-- Created on: 1996-01-30
-- Created by: Christian CAILLET
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package IGESControl

    ---Purpose : This package provide external access and control to use IGES
    --           See also IGESToBRep for reading IGES to Shapes

uses

    TColStd,
    Interface,
    Transfer,
    IFSelect,
    XSControl,
    IGESData,
    TopoDS,
    IGESToBRep,
    ShapeExtend, 
    Message

is

    class Controller;
    class Writer;
    class Reader;
    class ActorWrite;
    class IGESBoundary;
    class AlgoContainer;
    class ToolContainer;

end;
