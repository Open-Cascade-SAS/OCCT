-- Created on: 1992-09-04
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package IntStart

    	---Purpose: This package provides generic algorithms to
    	--          find specific points (points on boundaries
    	--          and points inside a surface) used as starting
    	--          points for marching algorithms.

        ---Level: Internal
        --
        -- All the methods of the classes of this package are Internal.
	--

uses Standard, MMgt, TCollection, StdFail, TopAbs, GeomAbs, gp, IntSurf, math

is

    generic class Segment;
    
    generic class PathPoint;

    generic class SearchOnBoundaries, ThePathPoint, SequenceOfPathPoint, 
                                      TheSegment, SequenceOfSegment;

    deferred class SITopolTool;

    generic class SearchInside;


end IntStart;



