-- File:        CompositeCurveSegment.cdl
-- Created:     Mon Dec  4 12:02:24 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWCompositeCurveSegment from RWStepGeom

	---Purpose : Read & Write Module for CompositeCurveSegment

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     CompositeCurveSegment from StepGeom,
     EntityIterator from Interface

is

	Create returns RWCompositeCurveSegment;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable CompositeCurveSegment from StepGeom);

	WriteStep (me; SW : in out StepWriter; ent : CompositeCurveSegment from StepGeom);

	Share(me; ent : CompositeCurveSegment from StepGeom; iter : in out EntityIterator);

end RWCompositeCurveSegment;
