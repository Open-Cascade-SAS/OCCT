-- Created on: 1997-10-22
-- Created by: Jean-Louis Frenkel
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

---Copy:	 Matra Datavision 1997

deferred class Application from CDM inherits Transient from Standard

uses Document           from CDM,
     MetaData           from CDM,
     Reference          from CDM,
     MessageDriver      from CDM,
     Manager            from Resource,
     ExtendedString     from TCollection
is

    Retrieve(me: mutable; aMetaData: MetaData from CDM; UseStorageConfiguration: Boolean from Standard)
    returns mutable Document from CDM
    is deferred private;


    DocumentVersion(me: mutable; aMetaData: MetaData from CDM)
    returns Integer from Standard
    is deferred private;
    ---Purpose: returns -1 if the metadata has no modification counter.
    
    SetDocumentVersion(me; aDocument: Document from CDM; aMetaData: MetaData from CDM)
    is protected;

    SetReferenceCounter(me:mutable ; aDocument: Document from CDM; aReferenceCounter: Integer from Standard)
    is protected;
    
    Resources(me: mutable)
    returns Manager from Resource
    is deferred;
    ---Purpose: the manager returned by  this virtual  method will be
    --          used to search for Format`.Retrieval  resource items. 
    --          
    
    MessageDriver(me: mutable) returns MessageDriver from CDM
    is virtual;
    ---Purpose: By default returns a NullMessageDriver;

    BeginOfUpdate(me:mutable; aDocument: Document from CDM)
    is virtual;
    ---Purpose: this method is called before the update of a document.
    --         By default, writes in MessageDriver().

    EndOfUpdate(me:mutable; aDocument: Document from CDM; Status: Boolean from Standard; ErrorString: ExtendedString from TCollection)
    is virtual;
    ---Purpose: this method is called affter the update of a document.
    --         By default, writes in MessageDriver().

    Write(me: mutable; aString: ExtString from Standard);
    ---Purpose: writes the string in the application MessagerDriver.

friends     

    class Reference from CDM,
    class MetaData from CDM

end Application from CDM;
