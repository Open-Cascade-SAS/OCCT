-- Created on: 1993-01-09
-- Created by: CKY / Contract Toubro-Larsen ( SIVA )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SelectedComponent from IGESSolid  inherits IGESEntity

        ---Purpose: defines SelectedComponent, Type <182> Form Number <0>
        --          in package IGESSolid
        --          The Selected Component entity provides a means of
        --          selecting one component of a disjoint CSG solid

uses

        BooleanTree     from IGESSolid,
        XYZ             from gp,
        Pnt             from gp

is

        Create returns mutable SelectedComponent;

        -- Specific Methods pertaining to the class

        Init (me        : mutable;
              anEntity  : BooleanTree;
              selectPnt : XYZ);
        ---Purpose : This method is used to set the fields of the class
        --           SelectedComponent
        --       - anEntity  : the Boolean tree entity
        --       - selectPnt : Point in or on the desired component

        Component(me) returns BooleanTree;
        ---Purpose : returns the Boolean tree entity

        SelectPoint(me) returns Pnt;
        ---Purpose : returns the point on/in the selected component

        TransformedSelectPoint(me) returns Pnt;
        ---Purpose : returns the point on/in the selected component
        -- after applying TransformationMatrix

fields

--
-- Class    : IGESSolid_SelectedComponent
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class SelectedComponent.
--
-- Reminder : A SelectedComponent instance is defined by :
--            a pointer to the Boolean Tree entity(Entity) and the X, Y
--            and Z components (X,Y,Z) of a selected point.

        theEntity      : BooleanTree;
            -- the desired boolean tree entity

        theSelectPoint : XYZ;
            -- the X, Y and Z coordinates of the point

end SelectedComponent;
