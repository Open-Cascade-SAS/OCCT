-- Created on: 1993-06-11
-- Created by: Martine LANGLOIS
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package StepToGeom

--- Purpose: Creation des entites geometriques de Geom a partir du schema 
--  StepGeom (Part42, geometric)

uses  gp, Geom, Geom2d, StepGeom, StdFail

is

private deferred class Root;
class MakeCartesianPoint;
class MakeCartesianPoint2d;
class MakeAxisPlacement;
class MakeAxis1Placement;
class MakeAxis2Placement;
class MakeDirection;
class MakeDirection2d;
class MakeVectorWithMagnitude;
class MakeVectorWithMagnitude2d;
class MakeCurve;
class MakeTrimmedCurve;
class MakeTrimmedCurve2d;
class MakeCurve2d;
class MakeConic;
class MakeConic2d;
class MakeBoundedCurve;
class MakeBoundedCurve2d;
class MakeEllipse;
class MakeEllipse2d;
class MakeHyperbola;
class MakeHyperbola2d;
class MakeParabola;
class MakeParabola2d;
class MakeCircle;
class MakeCircle2d;
class MakeBSplineCurve;
class MakeBSplineCurve2d;
class MakeLine;
class MakeLine2d;
class MakePolyline;
class MakePolyline2d;
class MakePlane;
class MakeSurface;
class MakeBoundedSurface;
class MakeElementarySurface;
class MakeSweptSurface;
class MakeConicalSurface;
class MakeCylindricalSurface;
class MakeRectangularTrimmedSurface;
class MakeSphericalSurface;
class MakeSurfaceOfLinearExtrusion;
class MakeSurfaceOfRevolution;
class MakeToroidalSurface;
class MakeBSplineSurface;
class MakeTransformation3d;
class MakeTransformation2d;

-- class CheckSurfaceClosure;

end StepToGeom;
