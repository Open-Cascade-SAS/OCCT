-- Created on: 1993-08-06
-- Created by: Denis PASCAL
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



package GraphDS 

    ---Purpose: This  package  <GraphDS> provides  generic  classes to
    --          describe transient graph data structure.

uses Standard,
     MMgt,
     TCollection,
     TColStd

is
    enumeration EntityRole is 
    	OnlyInput, 
    	OnlyOutput, 
    	InputAndOutput
    end EntityRole;
    
    enumeration RelationRole is 
        OnlyFront, 
    	OnlyBack, 
    	FrontAndBack
    end RelationRole;

    class EntityRoleMap instantiates DataMap from TCollection
                                    (Transient  from Standard,
				     EntityRole from GraphDS,
				     MapTransientHasher from TColStd);

    generic class DirectedGraph,
                  Vertex,
		  Edge,
		  VerticesIterator,
		  EdgesIterator;
		 
    
    generic class RelationGraph,
                  Entity,
		  Relation,
    	    	  EntitiesIterator,
                  IncidentEntitiesIterator,
                  RelationsIterator,
                  IncidentRelationsIterator;		  

end GraphDS;










