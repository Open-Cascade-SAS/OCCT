-- File:	StepToGeom_MakeConicalSurface.cdl
-- Created:	Mon Jun 14 16:05:32 1993
-- Author:	Martine LANGLOIS
---Copyright:	 Matra Datavision 1993

class MakeConicalSurface from StepToGeom

    ---Purpose: This class implements the mapping between class
    --          ConicalSurface from StepGeom which describes a
    --          conical_surface from Prostep and ConicalSurface from Geom 

uses ConicalSurface from Geom,
     ConicalSurface from StepGeom

is 

    Convert ( myclass; SS : ConicalSurface from StepGeom;
                       CS : out ConicalSurface from Geom )
    returns Boolean from Standard;

end MakeConicalSurface;
