-- Created on: 1999-05-11
-- Created by: Sergei ZERTCHANINOV
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class EdgeConnect  from ShapeFix

    ---Purpose : Makes vertices to be shared to connect edges,
    --           updates positions and tolerances for shared vertices.
    --           Accepts edges bounded by two vertices each.

uses 
    DataMapOfShapeShape from TopTools,
    DataMapOfShapeListOfShape from TopTools,
    Edge from TopoDS, Shape from TopoDS

is

    Create returns EdgeConnect from ShapeFix;

    Add (me : in out; aFirst : Edge from TopoDS; aSecond : Edge from TopoDS);
    ---Purpose : Adds information on connectivity between start vertex
    --           of second edge and end vertex of first edge,
    --           taking edges orientation into account

    Add (me : in out; aShape : Shape from TopoDS);
    ---Purpose : Adds connectivity information for the whole shape.
    --           Note: edges in wires must be well ordered
    --           Note: flag Closed should be set for closed wires

    Build (me : in out);
    ---Purpose : Builds shared vertices, updates their positions and tolerances

    Clear (me : in out);
    ---Purpose : Clears internal data structure

fields

    myVertices : DataMapOfShapeShape from TopTools;       -- Map of pairs (vertex, shared)
    myLists    : DataMapOfShapeListOfShape from TopTools; -- Map of pairs (shared, list of vertices/edges)

end EdgeConnect;
