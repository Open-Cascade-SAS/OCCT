-- Created on: 2001-04-24
-- Created by: Atelier IED
-- Copyright (c) 2001-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class LimitsAndFits  from StepShape    inherits TShared

    ---Purpose : Added for Dimensional Tolerances

uses
    HAsciiString from TCollection

is

    Create returns mutable LimitsAndFits;

    Init (me : mutable; form_variance, zone_variance, grade, source :
    	    	        HAsciiString from TCollection);

    FormVariance (me) returns HAsciiString from TCollection;
    SetFormVariance (me : mutable; form_variance : HAsciiString from TCollection);

    ZoneVariance (me) returns HAsciiString from TCollection;
    SetZoneVariance (me : mutable; zone_variance : HAsciiString from TCollection);

    Grade (me) returns HAsciiString from TCollection;
    SetGrade (me : mutable; grade : HAsciiString from TCollection);

    Source (me) returns HAsciiString from TCollection;
    SetSource (me : mutable; source : HAsciiString from TCollection);

fields

    theFormVariance : HAsciiString from TCollection;
    theZoneVariance : HAsciiString from TCollection;
    theGrade  : HAsciiString from TCollection;
    theSource : HAsciiString from TCollection;

end LimitsAndFits;
