-- Created by: Peter KURNEV
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

package BOPTools 

        ---Purpose: 

uses
    gp,  
    Bnd,
    TopAbs, 
    Geom,   
    Geom2d,
    GeomAPI, 
    BRepClass3d,
    TopoDS, 
    TopTools, 
    IntTools,   
    ProjLib,
    --                 
    BOPCol, 
    BOPInt 
is 

    -- 
    -- classes
    -- 
    class ShapeSet; 
    class EdgeSet; 
    class AlgoTools; 
    class Set; 
    class SetMapHasher;  
    class AlgoTools2D; 
    class AlgoTools3D;
    -- 
    imported MapOfSet;
    imported DataMapOfShapeSet;
    --
    -- primitives
    --
    imported ListOfShapeSet from BOPTools;
    imported ListOfEdgeSet from BOPTools;
    imported ConnexityBlock from BOPTools;
    imported ListOfConnexityBlock from BOPTools;
    imported CoupleOfShape from BOPTools;
    imported ListOfCoupleOfShape from BOPTools;
    --
    --  static methods 
    -- 
    MapShapes(S : Shape from TopoDS;
                  M : in out MapOfShape from BOPCol); 
               
    MapShapes(S : Shape from TopoDS;
                  M : in out IndexedMapOfShape from BOPCol); 
              
    MapShapes(S : Shape from TopoDS;
                  T : ShapeEnum from TopAbs;
                  M : in out IndexedMapOfShape from BOPCol);
          

    MapShapesAndAncestors
            (S  : Shape from TopoDS;
             TS : ShapeEnum from TopAbs;
         TA : ShapeEnum from TopAbs;
         M  : in out IndexedDataMapOfShapeListOfShape from BOPCol);
    
end BOPTools;
