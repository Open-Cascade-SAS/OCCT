-- Created on: 1993-03-23
-- Created by: BBL
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ColorCubeColorMap from Aspect inherits ColorMap from Aspect

	---Version: 0.0

	---Purpose: This class defines a ColorCube ColorMap object.
	---Keywords:
	---Warning:
	---References:

uses
	Color		from Quantity,
	ColorMapEntry 	from Aspect

raises
	BadAccess 	from Aspect,
	RangeError from Standard

is
	Create( base_pixel, redmax,   redmult,
			    greenmax, greenmult,
			    bluemax,  bluemult : in Integer from Standard )
	returns mutable ColorCubeColorMap from Aspect
	raises RangeError from Standard ;
	---Level: Public
	---Purpose : Create a ColorCube ColorMap.

	ColorCubeDefinition( me : in ;
			  base_pixel,
			  redmax,   redmult,
			  greenmax, greenmult,
			  bluemax,  bluemult : out Integer from Standard );

	FindColorMapIndex ( me ;
			AColorMapEntryIndex : Integer from Standard )
	returns Integer from Standard
	raises BadAccess from Aspect ;
	---Level: Public
	---Purpose: Returns the index in the ColorMap of the
	--	    ColorMapEntry.Index() equal to <AnEntryIndex>.
	--  Warning: Raises BadAccess if the index is not defined in the
	--	    ColorMap.

	FindEntry ( me ; AColorMapEntryIndex : Integer from Standard )
	returns ColorMapEntry from Aspect
	raises BadAccess from Aspect ;
	---Level: Public
	---Purpose: Returns the ColorMapEntry with ColorMapEntry.Index()
	--	    equal to <AnEntryIndex>.
	--  Warning: Raises BadAccess if the index is not defined in the
	--	    ColorMap.
    	---C++: return const &

	NearestColorMapIndex( me ; aColor : Color from Quantity )
	returns Integer from Standard ;
	---Level: Public
	---Purpose: Returns the index in the ColorMap of the nearest
	--	    matching ColorMapEntry

	NearestEntry( me ; aColor : Color from Quantity )
	returns ColorMapEntry from Aspect ;
	---Level: Public
	---Purpose: Returns the nearest ColorMapEntry that match aColor .
    	---C++: return const &

        AddEntry (me : mutable; aColor : Color from Quantity)
                returns Integer from Standard;
        ---Level: Public
        ---Purpose: Search an identical color entry in the color map <me>
        -- or returns the nearest ColorMapEntry Index.

fields
	mybasepixel 		 : Integer from Standard ;
	mygreenmax , mygreenmult : Integer from Standard ;
	myredmax   , myredmult   : Integer from Standard ;
	mybluemax  , mybluemult  : Integer from Standard ;
		-- ColorCube definition for a ColorCube ColorMap.

end ColorCubeColorMap ;
