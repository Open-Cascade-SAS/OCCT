-- File:	MakeMirror.cdl
-- Created:	Mon Sep 28 11:52:47 1992
-- Author:	Remi GILET
--		<reg@sdsun2>
---Copyright:	 Matra Datavision 1992

class MakeMirror

from GCE2d

    ---Purpose: This class implements elementary construction algorithms for a
    -- symmetrical transformation in 2D space about a point
    -- or axis. The result is a Geom2d_Transformation transformation.
    -- A MakeMirror object provides a framework for:
    -- -   defining the construction of the transformation,
    -- -   implementing the construction algorithm, and
    -- -   consulting the result.

uses Pnt2d          from gp,
     Ax2d           from gp,
     Dir2d          from gp,
     Lin2d          from gp,
     Transformation from Geom2d,
     Real           from Standard
     
is

Create(Point : Pnt2d from gp) returns MakeMirror;
    ---Puprose: Make a symetry transformation of center <Point>.

Create(Axis : Ax2d from gp) returns MakeMirror;
    ---Puprose: Make a symetry transformation of axis <Axis>.

Create(Line : Lin2d from gp) returns MakeMirror;
    ---Puprose: Make a symetry transformation of axis <Line>.

Create(Point : Pnt2d from gp;
       Direc : Dir2d from gp) returns MakeMirror;
    ---Purpose: Make a symetry transformation af axis defined by 
    --          <Point> and <Direc>.

Value(me) returns Transformation from Geom2d
    is static;
    ---C++: return const&
    ---Purpose: Returns the constructed transformation.

Operator(me) returns Transformation from Geom2d
    is static;
    ---C++: return const&
    ---C++: alias "Standard_EXPORT operator Handle_Geom2d_Transformation() const;"

fields

    TheMirror : Transformation from Geom2d;

end MakeMirror;

