-- Created on: 1999-11-26
-- Created by: Andrey BETENEV
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0

class ActionRequestAssignment from StepBasic
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity ActionRequestAssignment

uses
    VersionedActionRequest from StepBasic

is
    Create returns ActionRequestAssignment from StepBasic;
	---Purpose: Empty constructor

    Init (me: mutable; aAssignedActionRequest: VersionedActionRequest from StepBasic);
	---Purpose: Initialize all fields (own and inherited)

    AssignedActionRequest (me) returns VersionedActionRequest from StepBasic;
	---Purpose: Returns field AssignedActionRequest
    SetAssignedActionRequest (me: mutable; AssignedActionRequest: VersionedActionRequest from StepBasic);
	---Purpose: Set field AssignedActionRequest

fields
    theAssignedActionRequest: VersionedActionRequest from StepBasic;

end ActionRequestAssignment;
