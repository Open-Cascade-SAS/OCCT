-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ShapeDefinition from StepRepr inherits SelectType from StepData

	-- <ShapeDefinition> is an EXPRESS Select Type construct translation.
	-- it gathers : ProductDefinitionShape, ShapeAspect, ShapeAspectRelationship

uses

	ProductDefinitionShape,
	ShapeAspect,
	ShapeAspectRelationship
is

	Create returns ShapeDefinition;
	---Purpose : Returns a ShapeDefinition SelectType

	CaseNum (me; ent : Transient) returns Integer;
	---Purpose: Recognizes a ShapeDefinition Kind Entity that is :
	--        1 -> ProductDefinitionShape
	--        2 -> ShapeAspect
	--        3 -> ShapeAspectRelationship
	--        0 else

	ProductDefinitionShape (me) returns any ProductDefinitionShape;
	---Purpose : returns Value as a ProductDefinitionShape (Null if another type)

	ShapeAspect (me) returns any ShapeAspect;
	---Purpose : returns Value as a ShapeAspect (Null if another type)

	ShapeAspectRelationship (me) returns any ShapeAspectRelationship;
	---Purpose : returns Value as a ShapeAspectRelationship (Null if another type)


end ShapeDefinition;

