-- Created on: 1991-07-18
-- Created by: Arnaud BOUZY
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package ExprIntrp 

	---Purpose: Describes an interpreter for GeneralExpressions, 
	--          GeneralFunctions, and GeneralRelations defined in 
	--          package Expr. 

uses Expr, MMgt, TCollection, TColStd

is

    deferred class Generator;
    
    class GenExp;
    
    class GenFct;
    
    class GenRel;
    
    private class Analysis;
    
    class SequenceOfNamedFunction instantiates 
    	Sequence from TCollection(NamedFunction from Expr);

    class SequenceOfNamedExpression instantiates 
    	Sequence from TCollection(NamedExpression from Expr);

    exception SyntaxError inherits Failure from Standard;
    
    private class StackOfGeneralExpression instantiates 
    	Stack from TCollection (GeneralExpression from Expr);
    
    private class StackOfGeneralRelation instantiates 
    	Stack from TCollection (GeneralRelation from Expr);

    private class StackOfGeneralFunction instantiates 
    	Stack from TCollection (GeneralFunction from Expr);
        
    
    private class StackOfNames instantiates 
    	Stack from TCollection (AsciiString from TCollection);

    Parse(gen : Generator; str : AsciiString from TCollection)
    returns Boolean
    is private;
    
end ExprIntrp;

