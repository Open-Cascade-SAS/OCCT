-- Created by: Tanya COOL
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Arrow from Prs2d inherits Line from Graphic2d
  
  ---Purpose: Constructs the primitive arrow

uses

    Drawer	      from Graphic2d,
    GraphicObject     from Graphic2d,
    Length            from Quantity,
    Array1OfShortReal from TShort,
    ExtendedString    from TCollection,
    Ax2d              from gp,
    TypeOfArrow       from Prs2d,
    FStream           from Aspect,
    HArray1OfPnt2d    from TColgp

is
	Create( aGraphicObject: GraphicObject from Graphic2d;
	        Location      : Ax2d from gp;
	        OpenAngle     : Real from Standard = 5.0;
		Length        : Real from Standard = 5.0;
            	theType       : TypeOfArrow from Prs2d = Prs2d_TOA_CLOSED )
	
	returns mutable Arrow from Prs2d;
	
	---Purpose: create an arrow:
   	--          "Location"  gives the location and direction,
   	--          "OpenAngle" gives the opening angle (in radians),
   	--          "Length"    gives the length.

	----------------------------------
	---Category: Draw and Pick
	----------------------------------

	Draw( me : mutable; aDrawer: Drawer from Graphic2d )
     	is static protected;
	---Level: Internal
	---Purpose: Draws the arrow <me>.

    	DrawElement( me : mutable; aDrawer: Drawer from Graphic2d;
                 anIndex: Integer from Standard)
        is redefined protected;
	---Level: Internal
	---Purpose: Draws element <anIndex> of the arrow <me>.

	DrawVertex( me : mutable; aDrawer: Drawer from Graphic2d;
        	                  anIndex: Integer from Standard)
        is redefined protected;
     	---Level: Internal
    	---Purpose: Draws vertex <anIndex> of the arrow <me>.
		
	ArrayOfPnt2d( me ; withTrsf: Boolean from Standard = Standard_False) returns HArray1OfPnt2d from TColgp;
	---Level: Public
	---C++: return const
	
	TypeOfArrow( me ) returns TypeOfArrow from Prs2d;
	---Level: Public
	---Purpose: Returns type of arrow
	--          Type is:
	--             TOA_OPENED,
        --             TOA_CLOSED,
        --             TOA_FILLED


    	Pick (me : mutable; X, Y: ShortReal from Standard;
		    	aPrecision: ShortReal from Standard;
		    	aDrawer: Drawer from Graphic2d)
	returns Boolean from Standard
	is static protected;
	---Level: Internal
	---Purpose: Returns Standard_True if the arrow <me> is picked,
	--	    Standard_False if not.

    	Save( me; aFStream: in out FStream from Aspect ) is virtual;
    
													
fields
 
	myXVert       : Array1OfShortReal from TShort;
	myYVert       : Array1OfShortReal from TShort;
        myTypeOfArrow : TypeOfArrow from Prs2d;
	
end Arrow from Prs2d;
