-- File:        AutoDesignPresentedItem.cdl
-- Created:     Fri Dec  1 11:11:14 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class AutoDesignPresentedItem from StepAP214 

    -- updated for CC1 Rev4 (usage of Select)

inherits PresentedItem from StepVisual

uses

	HArray1OfAutoDesignPresentedItemSelect from StepAP214, 
	AutoDesignPresentedItemSelect from StepAP214
is

	Create returns mutable AutoDesignPresentedItem;
	---Purpose: Returns a AutoDesignPresentedItem

	Init (me : mutable;
	      aItems : mutable HArray1OfAutoDesignPresentedItemSelect from StepAP214) is virtual;

	-- Specific Methods for Field Data Access --

	SetItems(me : mutable; aItems : mutable HArray1OfAutoDesignPresentedItemSelect);
	Items (me) returns mutable HArray1OfAutoDesignPresentedItemSelect;
	ItemsValue (me; num : Integer) returns AutoDesignPresentedItemSelect;
	NbItems (me) returns Integer;

fields

	items : HArray1OfAutoDesignPresentedItemSelect from StepAP214;

end AutoDesignPresentedItem;
