-- Created on: 2002-08-02
-- Created by: Alexander KARTOMIN  (akm)
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- NB:          This originates from BRepLProp being abstracted of BRep.

package LProp3d

    ---Purpose: Handles local properties of curves and surfaces from the 
    --          package Adaptor3d.
    -- SeeAlso: Package LProp.

uses Standard, gp, Adaptor3d, GeomAbs, LProp

is
    
    class CurveTool;
    class SurfaceTool;
    
                                            
    class CLProps from LProp3d 
            instantiates CLProps from LProp(HCurve     from Adaptor3d,
                                            Vec        from gp,
                                            Pnt        from gp,
                                            Dir        from gp,
                                            CurveTool  from LProp3d);

    class SLProps from LProp3d 
            instantiates SLProps from LProp(HSurface    from Adaptor3d,
                                            SurfaceTool from LProp3d);

    
end LProp3d;    
