-- File:	ItemLocation.cdl
-- Created:	Mon Jan 21 14:00:31 1991
-- Author:	Christophe MARION
--		<cma@topsn3>
---Copyright:	 Matra Datavision 1991



private class ItemLocation from TopLoc

	---Purpose: An ItemLocation is an elementary coordinate system
	--          in a Location.
	--          
	--          The  ItemLocation     contains :
	--          
	--          * The elementary Datum.
	--          
	--          * The exponent of the elementary Datum.
	--          
	--          * The transformation associated to the composition.
	--          

uses
    Datum3D   from TopLoc,
    Trsf      from gp,
    TrsfPtr from TopLoc
    
is
    Create(D : Datum3D      from TopLoc; 
    	   P : Integer      from Standard;
           fromTrsf : Boolean from Standard = Standard_False) returns ItemLocation from TopLoc;
	---Purpose: Sets the elementary Datum to <D>
	--          Sets the exponent to <P>

    Create(anOther : ItemLocation from TopLoc) returns ItemLocation from TopLoc;
    
    Assign(me : in out; anOther : ItemLocation from TopLoc) returns ItemLocation from TopLoc;
    ---C++: alias operator=
    ---C++: return &

    Destroy(me : in out);
    ---C++: alias ~

fields
    myDatum  : Datum3D   from TopLoc;
    myPower  : Integer   from Standard;
    myTrsf   : TrsfPtr   from TopLoc;

friends
    class Location from TopLoc
    
end ItemLocation;
