-- File:        ApplicationContextElement.cdl
-- Created:     Mon Dec  4 12:02:23 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWApplicationContextElement from RWStepBasic

	---Purpose : Read & Write Module for ApplicationContextElement

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     ApplicationContextElement from StepBasic,
     EntityIterator from Interface

is

	Create returns RWApplicationContextElement;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable ApplicationContextElement from StepBasic);

	WriteStep (me; SW : in out StepWriter; ent : ApplicationContextElement from StepBasic);

	Share(me; ent : ApplicationContextElement from StepBasic; iter : in out EntityIterator);

end RWApplicationContextElement;
