-- Created on: 1999-03-10
-- Created by: data exchange team
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class OrganizationItem from StepAP214 
inherits ApprovalItem from StepAP214
	

uses

	AppliedOrganizationAssignment from StepAP214,   	
    	Approval from StepBasic
is

    Create returns OrganizationItem;
	---Purpose : Returns a OrganizationItem SelectType

    CaseNum (me; ent : Transient) returns Integer is redefined;
	---Purpose: Recognizes a OrganizationItem Kind Entity that is :
    	
    	--        1 -> AppliedOrganizationAssignment
    	--        2 -> Approval  
    	--        3 -> AssemblyComponentUsageSubstitute
	--        4 -> DocumentFile
    	--        5 -> MaterialDesignation
    	--        6 -> MechanicalDesignGeometricPresentationRepresentation
	--        7 -> PresentationArea
    	--        8 -> Product
	--        9 -> ProductDefinition
    	--        10 -> ProductDefinitionFormation
	--        11 -> ProductDefinitionRelationship
	--        12 -> PropertyDefinition
    	--        13 -> ShapeRepresentation
    	--        14 -> SecurityClassification 
	--        0 else
	
    AppliedOrganizationAssignment (me) returns any AppliedOrganizationAssignment;
	---Purpose : returns Value as a AppliedOrganizationAssignment (Null if another type)
	
    Approval (me) returns any Approval;
    	---Purpose : returns Value as a Approval (Null if another type)
	
	
end OrganizationItem;
