-- Created by: DCB
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


private class TextManager from PlotMgt inherits TextManager from MFT 

uses
  Length           from Quantity,
  PlaneAngle       from Quantity,
  TypeOfText       from Aspect,
  PlotterDriver    from PlotMgt,
  PlotterDriverPtr from PlotMgt

is
  -------------------------
  -- Category: Constructors
  -------------------------
  Create (aDriver : PlotterDriver from PlotMgt)
  returns mutable TextManager from PlotMgt;

  -------------------------
  -- Category: Draw methods
  -------------------------
  BeginString (me: mutable;
               X,Y: Length from Quantity;
               anOrientation: PlaneAngle from Quantity;
               aWidth,aHeight: Length from Quantity;
               aSlant: PlaneAngle from Quantity;
               aPaintType: Integer from Standard) is redefined;
  ---Purpose: Calls when string drawing is started.
  --          with a string aspect <aPaintType> :
  --            0 for filled string
  --            1 for stroke string
  --            2 for outline string
  --          The origine of the string <X>,<Y>,
  --          The orientation of the string <anOrientation>,
  --          The medium size of the char <aWidth,aHeight>,
  --          The Slant of the char <aSlant>,

  BeginChar (me: mutable;
             aCharCode: Integer from Standard;
             X,Y: Length from Quantity)
  returns Boolean from Standard is redefined;
  ---Purpose: Calls when a char drawing is started
  --          and give the current string position for this char.
  --          and give the relative char position from the beginning
  --          of the string.
  --The application can returns FALSE for skipping the char drawing.

  SetCharBoundingBox (me: mutable;
                      X1,Y1,X2,Y2,X3,Y3,X4,Y4: Length from Quantity) 
  returns Boolean from Standard is redefined;
  ---Purpose: Calls to defines the current char bounding-box. 
  -- The application can returns FALSE for ending the char drawing.

  SetCharEncoding (me: mutable;
                   anEncoding: CString from Standard)
  returns Boolean from Standard is redefined;
  ---Purpose: Calls to defines the current char encoding.
  --  Warning: The application can returns FALSE for skipping the char drawing.

  Moveto (me: mutable; X,Y: Length from Quantity) 
  returns Boolean from Standard is redefined;
  ---Purpose: Calls to sets the current string position. 
  -- The application can returns FALSE for ending the char drawing.

  Lineto (me: mutable; X,Y: Length from Quantity) 
  returns Boolean from Standard is redefined;
  ---Purpose: Calls to drawn to the current string position. 
  -- The application can returns FALSE for ending the char drawing.

  Curveto (me: mutable; X1,Y1,X2,Y2,X3,Y3,X4,Y4: Length from Quantity)
  returns Boolean from Standard is redefined;
  ---Purpose: Calls to drawn to the current string position.
  --          The application can drawn the curve defined by
  --          his descriptor P1,P2,P3,P4 or
  --          returns FALSE to let the interpretor compute the curve
  --          vectors.

  ClosePath (me: mutable) is redefined;
  ---Purpose: Calls when a char path drawing is ended 

  EndChar (me: mutable; X,Y: Length from Quantity)
  returns Boolean from Standard is redefined;
  ---Purpose: Calls when a char drawing is ended
  --          and give the relative char ending position from the
  --          beginning of the string.
  --          The application can returns FALSE for skipping the string
  --          drawing.

  EndString (me: mutable ) is redefined;
  ---Purpose: Calls when string drawing is ended (Normally the last call).

  -- Category: Private methods
  -------------------------
  SetTextAttribs (me: mutable;
                  aTextColor: Integer from Standard;
                  aTypeOfText: TypeOfText from Aspect;
                  anUnderlinePosition: Length from Quantity = 0.0)
  is private;
  ---Purpose: Sets the current attribs of the text.

fields
  myDriver           : PlotterDriverPtr from PlotMgt;

friends
  class PlotterDriver from PlotMgt

end TextManager from PlotMgt;
