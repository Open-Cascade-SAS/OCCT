-- Created on: 1991-05-14
-- Created by: Laurent PAINNOT
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class GaussSingleIntegration from math
    	---Purpose:
    	-- This class implements the integration of a function of a single variable
    	-- between the parameter bounds Lower and Upper.
    	--  Warning: Order must be inferior or equal to 61.


uses Function from math,
     OStream from Standard

raises NotDone from StdFail

is
     Create
     returns GaussSingleIntegration;
     
     Create(F: in out Function; Lower, Upper: Real; Order: Integer)
     	---Purpose:
     	-- The Gauss-Legendre integration with N = Order points of integration,
     	-- is done on the function F between the bounds Lower and Upper. 
    
     returns GaussSingleIntegration;
     
     Create(F: in out Function; Lower, Upper: Real; Order: Integer; Tol: Real)
     	---Purpose:
     	-- The Gauss-Legendre integration with N = Order points of integration  and 
     	-- given tolerance = Tol is done on the function F between the bounds  
     	-- Lower and Upper. 
    
     returns GaussSingleIntegration;

     Perform(me: in out; F: in out Function; Lower, Upper: Real; Order: Integer)      
	---Purpose:  perfoms  actual  computation  
     is private;
	
     IsDone(me)
     	---Purpose: returns True if all has been correctly done.
    	---C++: inline

     returns Boolean
     is static;
     
     
     Value(me)
     	---Purpose: returns the value of the integral.
    	---C++: inline

     returns Real
     raises NotDone
     is static;


    Dump(me; o: in out OStream)
    	---Purpose: Prints information on the current state of the object.

    is static;


fields

Val: Real;
Done: Boolean;

end GaussSingleIntegration;
