-- Created on: 1995-06-02
-- Created by: Xavier BENVENISTE
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class SameParameter from Approx

    ---Purpose: Approximation of a  PCurve  on a surface to  make  its
    --          parameter be the same that the parameter of a given 3d
    --          reference curve.

uses     
         HSurface        from   Adaptor3d,
         HCurve          from   Adaptor3d,
         HCurve2d        from   Adaptor2d,
         Surface         from   Geom,
         Curve           from   Geom,
         Curve           from   Geom2d,
    	 BSplineCurve    from   Geom2d  

raises  OutOfRange        from Standard,
        ConstructionError from Standard

is  

    Create (C3D  :  Curve    from  Geom; 
            C2D  :  Curve    from  Geom2d;
	    S    :  Surface  from  Geom; 
            Tol  :  Real)   

    returns  SameParameter    from  Approx 
    ---Purpose: 
    --  Warning: the C3D and C2D must have the same parametric domain.
    --           
    raises ConstructionError; 


    Create (C3D  :  HCurve    from  Adaptor3d; 
            C2D  :  Curve     from  Geom2d;
	    S    :  HSurface  from  Adaptor3d; 
            Tol  :  Real)   

    returns  SameParameter    from  Approx 
    ---Purpose: 
    --Warning: the C3D and C2D must have the same parametric domain.
               
    raises ConstructionError; 
   

    Create (C3D  :  HCurve    from  Adaptor3d; 
            C2D  :  HCurve2d  from  Adaptor2d; 
	    S    :  HSurface  from  Adaptor3d; 
            Tol  :  Real)   

    returns  SameParameter    from  Approx 
   ---Purpose: 
    --  Warning: the C3D and C2D must have the same parametric domain.
    --           
    raises ConstructionError; 
   

    Build (me   : in out;
           Tol  :  Real from Standard)
    ---Purpose: Compute the Pcurve (internal use only).
    is static private;


    IsDone(me) returns Boolean from Standard;
    ---C++: inline
     
    TolReached(me) returns Real from Standard;
    ---C++: inline
     
     
    IsSameParameter(me)  
    ---C++: inline  

    ---Purpose: Tells whether the original data  had already the  same
    --          parameter up to  the tolerance :  in that case nothing
    --          is done.
    
    returns  Boolean  from Standard; 


    Curve2d(me)   
    ---C++: inline

    ---Purpose: Returns the 2D  curve that has  the same parameter  as
    --          the  3D curve once evaluated on  the surface up to the
    --          specified tolerance
    returns  BSplineCurve  from  Geom2d;


fields  

   mySameParameter  :  Boolean       from Standard;
   myDone           :  Boolean       from Standard;
   myTolReached     :  Real          from Standard;
   myCurve2d        :  BSplineCurve  from Geom2d;
   myHCurve2d       :  HCurve2d      from Adaptor2d;
   myC3d            :  HCurve        from Adaptor3d;
   mySurf           :  HSurface      from Adaptor3d;

end  SameParameter; 
