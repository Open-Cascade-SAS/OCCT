-- Created on: 1996-09-04
-- Created by: Christian CAILLET
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class ActorOfFinderProcess  from Transfer  inherits ActorOfProcessForFinder

    ---Purpose : The original class was renamed. Compatibility only
    --         
    --         ModeTrans : a simple way of transmitting a transfer mode from
    --         a user. To be interpreted for each norm

uses Finder, FinderProcess, ProcessForFinder, Binder

is

    Create  returns mutable ActorOfFinderProcess;

    ModeTrans (me : mutable) returns Integer;
    ---Purpose : Returns the Transfer Mode, modifiable
    ---C++ : return &

    Transferring (me : mutable; start : Finder; TP : mutable ProcessForFinder)
        returns mutable Binder  is redefined;
    -- calls the one below

    Transfer (me : mutable; start : Finder; TP : mutable FinderProcess)
        returns mutable Binder  is virtual;
    -- default calls TransferTransient if <start> is a TransientMapper,
    -- i.e. does nothing, to be redefined

    TransferTransient (me : mutable; start : Transient;
    	    	       TP : mutable FinderProcess)
	returns mutable Transient  is virtual;
    -- default does nothing, can be redefined
    -- usefull when a result is Transient, simpler to define than Transfer with
    -- a Finder

fields

    themodetrans : Integer  is protected;

end ActorOfFinderProcess;
