-- Created on: 1994-10-28
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class FaceEdgeInterference from TopOpeBRepDS 
    inherits ShapeShapeInterference from TopOpeBRepDS

uses

    Transition from TopOpeBRepDS,
    Config     from TopOpeBRepDS,
    OStream    from Standard    
    
is

    Create(T : Transition from TopOpeBRepDS;
	   S : Integer from Standard;
	   G : Integer from Standard;
      	   GIsBound : Boolean from Standard;
    	   C : Config from TopOpeBRepDS)
	   
    	---Purpose: Create an interference of EDGE <G> on FACE <S>.

    returns FaceEdgeInterference from TopOpeBRepDS; 
	    
    Dump(me; OS : in out OStream from Standard) returns OStream
    is redefined;
    ---C++: return &
    
end FaceEdgeInterference from TopOpeBRepDS;
