-- Created on: 2002-01-16
-- Created by: Michael PONIKAROV
-- Copyright (c) 2002-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class ExtStringArray from TDataStd inherits Attribute from TDF

	---Purpose: ExtStringArray Attribute. Handles an
    	-- array of UNICODE strings (represented by the
    	-- TCollection_ExtendedString class).

uses GUID                     from Standard,
     ExtendedString           from TCollection,
     HArray1OfExtendedString  from TColStd, 
     Attribute                from TDF,     
     Label                    from TDF, 
     DeltaOnModification      from TDF,     
     RelocationTable          from TDF

is 

    ---Purpose: class methods
    --          =============

    GetID (myclass)   
    ---C++: return const &  
    ---Purpose: Returns the GUID for the attribute.  
    returns GUID from Standard;

    Set (myclass; label : Label from TDF; lower, upper : Integer from Standard; 
    	    	  isDelta : Boolean from Standard = Standard_False)
    ---Purpose: Finds, or creates, an ExtStringArray attribute with <lower> 
    --          and <upper> bounds.  The ExtStringArray  attribute is returned. 
    --          If <isDelta> == False, DefaultDeltaOnModification is used.     
    -- 	        If attribute is already set, all input parameters are refused 
    --          and the found attribute is returned.
    returns ExtStringArray from TDataStd;

    
    ---Category: ExtStringArray methods
    --          ===============

    Init(me : mutable; lower, upper : Integer from Standard);
    ---Purpose: Initializes the inner array with bounds from <lower> to <upper>

    SetValue (me : mutable; Index : Integer from Standard; Value : ExtendedString from TCollection);
    ---Purpose: Sets  the   <Index>th  element  of   the  array to <Value>

    Value (me; Index : Integer from Standard)
    ---Purpose: Returns the value of  the  <Index>th element of the array
    --
    ---C++: return const &
    ---C++: alias operator ()
    returns ExtendedString from TCollection;

    Lower (me) returns Integer from Standard;
    ---Purpose:  Return the lower bound.

    Upper (me) returns Integer from Standard;
    ---Purpose: Return the upper bound
    
    Length (me) returns Integer from Standard;
    ---Purpose: Return the number of elements of <me>.
   
    ChangeArray(me : mutable; newArray : HArray1OfExtendedString from TColStd; 
    	    	    	      isCheckItems : Boolean = Standard_True); 	    
    ---Purpose: Sets the inner array <myValue> of the ExtStringArray attribute to <newArray>. 
    -- If value of <newArray> differs from <myValue>, Backup performed and myValue 
    -- refers to new instance of HArray1OfExtendedString that holds <newArray> values
    -- If <isCheckItems> equal True each item of <newArray> will be checked with each 
    -- item of <myValue> for coincidence (to avoid backup). 
    
    Array(me) returns HArray1OfExtendedString from TColStd;
    ---Purpose: Return the inner array of the ExtStringArray attribute    
    ---C++: inline 
    ---C++: return const     
    
    GetDelta(me) returns Boolean from Standard;  
    ---C++: inline  
    
    SetDelta(me : mutable; isDelta : Boolean from Standard);     
    ---C++: inline  
    ---Purpose: for  internal  use  only!   
     
    RemoveArray(me  : mutable) is private;      
    ---C++: inline 
         
    ---Category: methodes of TDF_Attribute
    --           =========================

    Create returns mutable ExtStringArray from TDataStd; 
    
    ID (me)
    	---C++: return const & 
    returns GUID from Standard;

    Restore (me: mutable; With : Attribute from TDF);

    NewEmpty (me)
    returns mutable Attribute from TDF;

    Paste (me; Into : mutable Attribute from TDF;
	       RT   : mutable RelocationTable from TDF);    

    Dump(me; anOS : in out OStream from Standard)
    	returns OStream from Standard
    	is redefined;
	---C++: return &

    ---Category: methods to be added for using in DeltaOn Modification  
    --           =====================================================
    DeltaOnModification(me; anOldAttribute : Attribute from TDF)
    	returns DeltaOnModification from TDF
    	---Purpose : Makes a DeltaOnModification between <me> and
    	--         <anOldAttribute>.  
    	is redefined virtual;  
	
fields

    myValue : HArray1OfExtendedString from TColStd;
    myIsDelta : Boolean from Standard;   
     
friends   
    class DeltaOnModificationOfExtStringArray from TDataStd     
    
end ExtStringArray;
