-- Created on: 1992-09-24
-- Created by: Denis PASCAL
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


generic class DFSIterator from GraphTools 
	                 (Graph     as any;
                          Vertex    as any;
			  VHasher   as any;
                          VIterator as any)

    ---Purpose: This generic  class implement  the Depth  First Search
    --          algorithm from  a  Vertex with an iterator  to reached
    --          adjacent vertices of a  given  one.  The  interface of
    --          this algorithm is made as an iterator.

--generic class DFSIterator from GraphTools
--            (Graph     as any;
--    	       Vertex    as any;
--    	       VHasher   as MapHasher from TCollection (Vertex);
--	       VIterator as VertexIterator (Graph,Vertex))

raises NoMoreObject from Standard,
       NoSuchObject from Standard

    class DFSMap   instantiates IndexedMap from TCollection (Vertex,VHasher); 
    
is

    Create
    returns DFSIterator;
	---Purpose: Create an empty iterator.

    Perform (me : in out; G : Graph; V : Vertex);
	---Purpose: Initializes the research from <V> member vertex of
	--          <G>.
        ---Level: Public

    More (me) returns Boolean from Standard;
	---Purpose: Returns True if there are other vertices.
        ---Level: Public

    Next(me : in out) 
    	---Purpose: Set the iterator to the next vertex.
        ---Level: Public
    raises NoMoreObject from Standard;

    Value (me) returns any Vertex 
	---Purpose: returns the vertex  value for the current position
	--          of the iterator.
	---C++: return const &
        ---Level: Public
    raises NoSuchObject from Standard;


fields

    myVisited      : DFSMap from GraphTools;
    myCurrentIndex : Integer from Standard;

end DFSIterator;
    
    








