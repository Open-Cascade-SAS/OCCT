-- Created on: 1993-08-30
-- Created by: Modelistation
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class OrientedShapeMapHasher from TopTools 

uses
    Shape from TopoDS

is

    HashCode(myclass; S : Shape from TopoDS; Upper : Integer) returns Integer;
	---Purpose: Returns a HasCode value  for  the  Key <K>  in the
	--          range 0..Upper.
	--
	---C++: inline
	
    IsEqual(myclass; S1, S2 : Shape from TopoDS) returns Boolean;
	---Purpose: Returns True when the two keys are equal. Two same
	--          keys must have the same hashcode,  the contrary is
	--          not necessary.
	--          
	---C++: inline
	

end OrientedShapeMapHasher;
