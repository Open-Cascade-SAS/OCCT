-- File:        ConicalSurface.cdl
-- Created:     Mon Dec  4 12:02:24 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWConicalSurface from RWStepGeom

	---Purpose : Read & Write Module for ConicalSurface

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     ConicalSurface from StepGeom,
     EntityIterator from Interface

is

	Create returns RWConicalSurface;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable ConicalSurface from StepGeom);

	WriteStep (me; SW : in out StepWriter; ent : ConicalSurface from StepGeom);

	Share(me; ent : ConicalSurface from StepGeom; iter : in out EntityIterator);

end RWConicalSurface;
