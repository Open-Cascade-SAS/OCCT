-- File:	IGESSolid_ToolPlaneSurface.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolPlaneSurface  from IGESSolid

    ---Purpose : Tool to work on a PlaneSurface. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses PlaneSurface from IGESSolid,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolPlaneSurface;
    ---Purpose : Returns a ToolPlaneSurface, ready to work


    ReadOwnParams (me; ent : mutable PlaneSurface;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : PlaneSurface;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : PlaneSurface;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a PlaneSurface <ent>, from
    --           its specific (own) parameters

    DirChecker (me; ent : PlaneSurface) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : PlaneSurface;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : PlaneSurface; entto : mutable PlaneSurface;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : PlaneSurface;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolPlaneSurface;
