-- Created on: 1992-07-20
-- Created by: Arnaud BOUZY
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class Generator from ExprIntrp inherits TShared from MMgt

	---Purpose: Implements general services for interpretation of 
	--          expressions.

uses NamedExpression from Expr,
    NamedFunction from Expr,
    SequenceOfNamedFunction from ExprIntrp,
    SequenceOfNamedExpression from ExprIntrp,
    AsciiString from TCollection

is

    Initialize;
    
    Use(me : mutable; func : NamedFunction)
    ---Level: Internal 
    is static;

    Use(me : mutable; named : NamedExpression)
    ---Level: Internal 
    is static;
        
    GetNamed(me)
    returns SequenceOfNamedExpression
    ---C++: return const &
    ---Level: Internal 
    is static;
    
    GetFunctions(me)
    returns SequenceOfNamedFunction
    ---C++: return const &
    ---Level: Internal 
    is static;

    GetNamed(me; name : AsciiString)
    ---Purpose: Returns NamedExpression with name <name> already 
    --          interpreted if it exists. Returns a null handle if 
    --          not. 
    ---Level: Advanced
    returns any NamedExpression
    is static;
    
    GetFunction(me; name : AsciiString)
    ---Purpose: Returns NamedFunction with name <name> already 
    --          interpreted if it exists. Returns a null handle if 
    --          not.
    ---Level: Advanced 
    returns any NamedFunction
    is static;
    
fields

    myFunctions : SequenceOfNamedFunction;
    myNamed : SequenceOfNamedExpression;
    
end Generator;
