-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package TShort 

                             
uses TCollection

is


--                  Instantiations de TCollection                         --
--                  *****************************                         --
------------------------------------------------------------------------

--          
-- Instantiations Array1 -- *************************************************************
--       
    class Array1OfShortReal instantiates Array1 from TCollection (ShortReal);

--          
-- Instantiations HArray1 -- **************************************************************
--       
    class HArray1OfShortReal instantiates 
    	HArray1 from TCollection (ShortReal, Array1OfShortReal from TShort);

--          
-- Instantiations Array2 -- ***************************************************************************
--       
    class Array2OfShortReal instantiates 
	Array2 from TCollection (ShortReal);

--          
-- Instantiations HArray2
-- ****************************************************************************
--       
    class HArray2OfShortReal instantiates 
    	HArray2 from TCollection ( ShortReal,
	    	    	    	   Array2OfShortReal from TShort);
--                    
--       Instantiations Sequence      *****************************************************
--       
    class SequenceOfShortReal instantiates 
	Sequence from TCollection (ShortReal); 

--                    
--       Instantiations HSequence      ***********************************************
--       
class HSequenceOfShortReal instantiates 
	HSequence from TCollection (ShortReal,
    	    	    	    	    SequenceOfShortReal from TShort);
end TShort;

