-- Created on: 2000-09-08
-- Created by: data exchange team
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Volume from XCAFDoc inherits Attribute from TDF

	---Purpose: attribute to store volume

uses
     Attribute       from TDF,
     Label           from TDF,
     GUID            from Standard,
     Real            from Standard,
     RelocationTable from TDF
    
is
    Create returns Volume from XCAFDoc;
    
    ---Purpose: class methods
    --          =============

    GetID (myclass) 
    	---C++: return const &  
    returns GUID from Standard;

    ID (me)
    	---C++: return const & 
    returns GUID from Standard;

    Set (me: mutable; vol: Real from Standard);
    	---Purpose: Sets a value of volume

    Set (myclass ; label : Label from TDF; vol: Real from Standard)
    returns Volume from XCAFDoc;
        ---Purpose: Find, or create, an Volume attribute and set its value

    Get (me)
    returns Real from Standard;
    
    Get (myclass ; label : Label from TDF; vol: in out Real from Standard)
    returns Boolean from Standard;
        ---Purpose: Returns volume as argument
	--          returns false if no such attribute at the <label>

    Restore (me: mutable; With : Attribute from TDF);

    NewEmpty(me)
    returns Attribute from TDF;

    Paste (me; Into : Attribute from TDF;
	       RT   : RelocationTable from TDF);    

    Dump(me; anOS : in out OStream from Standard)
    returns OStream from Standard
    is redefined;
    ---C++: return &

fields

    myValue     : Real     from Standard;

end Volume from XCAFDoc;
