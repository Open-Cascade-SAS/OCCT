-- File:	PCDM_Reader.cdl
-- Created:	Thu Dec 18 09:16:27 1997
-- Author:	Jean-Louis Frenkel
--		<rmi@frilox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1997

deferred class Reader from PCDM inherits Transient from Standard


uses
    Document from CDM, 
    ExtendedString from TCollection,  
    Application from CDM, 
    ReaderStatus from PCDM

raises  DriverError from PCDM


is

    CreateDocument(me: mutable) returns Document from CDM
    is deferred;
    ---Purpose: this method is called by the framework before the read method.
    
    Read(me: mutable; aFileName: ExtendedString from TCollection; 
                      aNewDocument: mutable Document from CDM;
		      anApplication: Application from CDM)
    raises DriverError from PCDM
    is deferred;
    ---Purpose: retrieves the content of the file into a new Document.  
    
    GetStatus(me) returns ReaderStatus from PCDM; 
    ---C++: inline
fields 

    myReaderStatus : ReaderStatus from  PCDM is protected;
    
end Reader from PCDM;

