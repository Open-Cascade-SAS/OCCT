-- Created on: 1993-06-15
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PaveSet from TopOpeBRepBuild 
    inherits LoopSet from TopOpeBRepBuild

---Purpose: 
-- class providing an exploration of a set of vertices to build edges.
-- It is similar to LoopSet from TopOpeBRepBuild where Loop is Pave.

uses 
    
    Shape from TopoDS,
    Edge from TopoDS,
    Loop from TopOpeBRepBuild,
    Pave from TopOpeBRepBuild,
    ListOfPave from TopOpeBRepBuild,
    ListIteratorOfListOfPave from TopOpeBRepBuild
    
is

    Create(E : Shape from TopoDS) returns PaveSet from TopOpeBRepBuild;
    ---Purpose: Create a Pave set on edge <E>. It contains <E> vertices. 

    RemovePV(me:in out; B : Boolean); -- particular case B = T/F : try/don't try
    -- to remove Pave in Prepare() (T by default)
		
    Append(me : in out; PV : Pave from TopOpeBRepBuild) is static;
    ---Purpose: Add <PV> in the Pave set.
    
    -- === start signature LoopSet
    InitLoop(me : in out) is redefined;
    MoreLoop(me) returns Boolean is redefined;
    NextLoop(me : in out) is redefined;
    Loop(me) returns Loop from TopOpeBRepBuild is redefined;
    ---C++: return const &
    -- === end signature LoopSet

    Edge(me) returns Edge from TopoDS is static;
    ---C++: return const &

    HasEqualParameters(me : in out) returns Boolean is static;
    EqualParameters(me) returns Real is static;
    ClosedVertices(me : in out) returns Boolean is static;

    Prepare(me : in out) is static private;
    SortPave(myclass; Lin:ListOfPave; Lout:out ListOfPave);
    
fields

    myEdge       : Edge from TopoDS;
    myVertices   : ListOfPave from TopOpeBRepBuild;
    myVerticesIt : ListIteratorOfListOfPave from TopOpeBRepBuild;

    myHasEqualParameters : Boolean from Standard;
    myEqualParameters    : Real from Standard;
    myClosed             : Boolean from Standard;
    myPrepareDone        : Boolean from Standard;
    myRemovePV : Boolean;
    
end PaveSet from TopOpeBRepBuild;
