-- Created on: 1996-09-04
-- Created by: Christian CAILLET
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ActorOfTransientProcess  from Transfer  inherits ActorOfProcessForTransient from Transfer

    ---Purpose : The original class was renamed. Compatibility only

uses Transient, TransientProcess, ProcessForTransient, Binder

is

    Create  returns mutable ActorOfTransientProcess;

    Transferring (me : mutable; start : Transient; TP : mutable ProcessForTransient)
        returns mutable Binder  is redefined;
    -- calls the one below

    Transfer (me : mutable; start : Transient; TP : mutable TransientProcess)
        returns mutable Binder  is virtual;
    -- default calls TransferTransient i.e. does nothing, to be redefined

    TransferTransient (me : mutable; start : Transient;
    	    	       TP : mutable TransientProcess)
	returns mutable Transient  is virtual;
    -- default does nothing, can be redefined
    -- usefull when a result is Transient, simpler to define than Transfer with
    -- a Binder

end ActorOfTransientProcess;
