-- Created on: 1995-12-19
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Loop from TopOpeBRepBuild inherits TShared from MMgt

---Purpose: 
-- a Loop is an existing shape (Shell,Wire) or a set
-- of shapes (Faces,Edges) which are connex.
-- a set of connex shape is represented by a BlockIterator

uses

    Shape from TopoDS,
    BlockIterator from TopOpeBRepBuild,
    ShapeEnum from TopAbs

is

    Create(S : Shape from TopoDS) returns mutable Loop;
    Create(BI : BlockIterator) returns mutable Loop;
	
    IsShape(me) returns Boolean from Standard is virtual;

    Shape(me) returns Shape from TopoDS is virtual;
    ---C++: return const &
    -- only when IsShape() is true
    
    BlockIterator(me) returns BlockIterator is static;
    ---C++: return const &
    -- only when IsShape() is false

    Dump(me) is virtual;	

fields

    myIsShape       : Boolean from Standard is protected;
    myShape         : Shape from TopoDS     is protected;
    myBlockIterator : BlockIterator         is protected;

end Loop from TopOpeBRepBuild;
