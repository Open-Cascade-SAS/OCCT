-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class CurveStyleFont from StepVisual 

inherits TShared from MMgt

uses

	HAsciiString from TCollection, 
	HArray1OfCurveStyleFontPattern from StepVisual, 
	CurveStyleFontPattern from StepVisual
is

	Create returns mutable CurveStyleFont;
	---Purpose: Returns a CurveStyleFont

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aPatternList : mutable HArray1OfCurveStyleFontPattern from StepVisual) is virtual;

	-- Specific Methods for Field Data Access --

	SetName(me : mutable; aName : mutable HAsciiString);
	Name (me) returns mutable HAsciiString;
	SetPatternList(me : mutable; aPatternList : mutable HArray1OfCurveStyleFontPattern);
	PatternList (me) returns mutable HArray1OfCurveStyleFontPattern;
	PatternListValue (me; num : Integer) returns mutable CurveStyleFontPattern;
	NbPatternList (me) returns Integer;

fields

	name : HAsciiString from TCollection;
	patternList : HArray1OfCurveStyleFontPattern from StepVisual;

end CurveStyleFont;
