-- Created on: 1993-03-10
-- Created by: JCV
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class  SphericalSurface from Geom inherits ElementarySurface from Geom

        --- Purpose :  Describes a sphere.
    	-- A sphere is defined by its radius, and is positioned in
    	-- space by a coordinate system (a gp_Ax3 object), the
    	-- origin of which is the center of the sphere.
    	-- This coordinate system is the "local coordinate
    	-- system" of the sphere. The following apply:
    	-- - Rotation around its "main Axis", in the trigonometric
    	--   sense given by the "X Direction" and the "Y
    	--   Direction", defines the u parametric direction.
    	-- - Its "X Axis" gives the origin for the u parameter.
    	-- - The "reference meridian" of the sphere is a
    	--   half-circle, of radius equal to the radius of the
    	--   sphere. It is located in the plane defined by the
    	--   origin, "X Direction" and "main Direction", centered
    	--   on the origin, and positioned on the positive side of the "X Axis".
    	-- - Rotation around the "Y Axis" gives the v parameter
    	--   on the reference meridian.
    	-- - The "X Axis" gives the origin of the v parameter on
    	--   the reference meridian.
    	-- - The v parametric direction is oriented by the "main
    	--   Direction", i.e. when v increases, the Z coordinate
    	--   increases. (This implies that the "Y Direction"
    	--   orients the reference meridian only when the local
    	--   coordinate system is indirect.)
    	-- - The u isoparametric curve is a half-circle obtained
    	--   by rotating the reference meridian of the sphere
    	--   through an angle u around the "main Axis", in the
    	--   trigonometric sense defined by the "X Direction"
    	--   and the "Y Direction".
    	--   The parametric equation of the sphere is:
    	-- P(u,v) = O + R*cos(v)*(cos(u)*XDir + sin(u)*YDir)+R*sin(v)*ZDir
    	-- where:
    	-- - O, XDir, YDir and ZDir are respectively the
    	--   origin, the "X Direction", the "Y Direction" and the "Z
    	--   Direction" of its local coordinate system, and
    	-- - R is the radius of the sphere.
    	--   The parametric range of the two parameters is:
    	-- - [ 0, 2.*Pi ] for u, and
    	-- - [ - Pi/2., + Pi/2. ] for v.

uses Ax3      from gp, 
     Pnt      from gp, 
     Sphere   from gp,
     Trsf     from gp,
     Vec      from gp, 
     Curve    from Geom,
     Geometry from Geom

raises ConstructionError from Standard,
       RangeError        from Standard

is

  Create (A3 : Ax3; Radius : Real)   returns mutable SphericalSurface
        --- Purpose :
        --  A3 is the local coordinate system of the surface.
        --  At the creation the parametrization of the surface is defined
        --  such as the normal Vector (N = D1U ^ D1V) is directed away from
        --  the center of the sphere.
        --  The direction of increasing parametric value V is defined by the
        --  rotation around the "YDirection" of A2 in the trigonometric sense
        --  and the orientation of increasing parametric value U is defined 
        --  by the rotation around the main direction of A2 in the
        --  trigonometric sense.
        --  Warnings :
        --  It is not forbidden to create a spherical surface with 
        --  Radius = 0.0
     raises ConstructionError;
        --- Purpose : Raised if Radius < 0.0.


  Create (S : Sphere)   returns mutable SphericalSurface;
        --- Purpose :
        --  Creates a SphericalSurface from a non persistent Sphere from 
        --  package gp.


  SetRadius (me : mutable; R : Real)
     raises ConstructionError;
        --- Purpose : Assigns the value R to the radius of this sphere.
    	-- Exceptions Standard_ConstructionError if R is less than 0.0.


  SetSphere (me : mutable; S : Sphere);
    	--- Purpose : Converts the gp_Sphere S into this sphere.
      

  Sphere (me)  returns Sphere;
        --- Purpose : Returns a non persistent sphere with the same geometric
        --  properties as <me>.


  UReversedParameter(me; U : Real) returns Real;
  	---Purpose: Computes the u parameter on the modified
    	-- surface, when reversing its u  parametric
    	-- direction, for any point of u parameter U on this sphere.
    	-- In the case of a sphere, these functions returns 2.PI - U.
        

  VReversedParameter(me; V : Real) returns Real;
  	---Purpose: Computes the v parameter on the modified
    	-- surface, when reversing its v parametric
    	-- direction, for any point of v parameter V on this sphere.
    	-- In the case of a sphere, these functions returns   -U.


  Area (me)   returns Real;
        --- Purpose : Computes the aera of the spherical surface.


  Bounds (me; U1, U2, V1, V2 : out Real);
        --- Purpose : Returns the parametric bounds U1, U2, V1 and V2 of this sphere.
    	-- For a sphere: U1 = 0, U2 = 2*PI, V1 = -PI/2, V2 = PI/2.


  Coefficients (me; A1, A2, A3, B1, B2, B3, C1, C2, C3, D : out Real);
       	--- Purpose : Returns the coefficients of the implicit equation of the 
       	--  quadric in the absolute cartesian coordinates system :
       	--  These coefficients are normalized.
       	--  A1.X**2 + A2.Y**2 + A3.Z**2 + 2.(B1.X.Y + B2.X.Z + B3.Y.Z) +
       	--  2.(C1.X + C2.Y + C3.Z) + D = 0.0


  Radius (me)  returns Real;

       	---Purpose: Computes the coefficients of the implicit equation of
       	-- this quadric in the absolute Cartesian coordinate system:
       	-- A1.X**2 + A2.Y**2 + A3.Z**2 + 2.(B1.X.Y + B2.X.Z + B3.Y.Z) +
       	-- 2.(C1.X + C2.Y + C3.Z) + D = 0.0
    	-- An implicit normalization is applied (i.e. A1 = A2 = 1.
    	-- in the local coordinate system of this sphere).
        
  Volume (me)  returns Real;
        --- Purpose : Computes the volume of the spherical surface.

  
  IsUClosed (me)  returns Boolean;
        --- Purpose : Returns True.


  IsVClosed (me)  returns Boolean;
        --- Purpose : Returns False.


  IsUPeriodic (me)  returns Boolean;
        --- Purpose : Returns True.


  IsVPeriodic (me) returns Boolean;
        --- Purpose : Returns False.


  UIso (me; U : Real)   returns mutable Curve;
        --- Purpose : Computes the U isoparametric curve.
        --  The U isoparametric curves of the surface are defined by the 
        --  section of the spherical surface with plane obtained by rotation
        --  of the plane (Location, XAxis, ZAxis) around ZAxis. This plane
        --  defines the origin of parametrization u.
        --  For a SphericalSurface the UIso curve is a Circle.
        -- Warnings : The radius of this circle can be zero.


  VIso (me; V : Real)  returns mutable Curve;
        --- Purpose : Computes the V isoparametric curve.
        --  The V isoparametric curves of the surface  are defined by 
        --  the section of the spherical surface with plane parallel to the
        --  plane (Location, XAxis, YAxis). This plane defines the origin of
        --  parametrization V.
        --  Be careful if  V is close to PI/2 or 3*PI/2 the radius of the 
        --  circle becomes tiny. It is not forbidden in this toolkit to 
        --  create circle with radius = 0.0
        --  For a SphericalSurface the VIso curve is a Circle.
        --  Warnings : The radius of this circle can be zero.


  D0 (me; U, V : Real; P : out Pnt);
        --- Purpose :
        --  Computes the  point P (U, V) on the surface.
        --  P (U, V) = Loc + Radius * Sin (V) * Zdir +
        --             Radius * Cos (V) * (cos (U) * XDir + sin (U) * YDir)
        --  where Loc is the origin of the placement plane (XAxis, YAxis)
        --  XDir is the direction of the XAxis and YDir the direction of
        --  the YAxis and ZDir the direction of the ZAxis.


  D1 (me; U, V : Real; P : out Pnt; D1U, D1V : out Vec);
        --- Purpose :
        --  Computes the current point and the first derivatives in the
        --  directions U and V.


  D2 (me; U, V : Real; P : out Pnt; D1U, D1V, D2U, D2V, D2UV : out Vec);
        --- Purpose :
        --  Computes the current point, the first and the second derivatives
        --  in the directions U and V.


  D3 (me; U, V : Real;  P : out Pnt; 
      D1U, D1V, D2U, D2V, D2UV, D3U, D3V, D3UUV, D3UVV : out Vec);
        --- Purpose :
        --  Computes the current point, the first,the second and the third 
        --  derivatives in the directions U and V.


  DN (me; U, V : Real; Nu, Nv : Integer)   returns Vec
        --- Purpose :
        --  Computes the derivative of order Nu in the direction u 
        --  and Nv in the direction v.
     raises RangeError;
        --- Purpose : Raised if Nu + Nv < 1 or Nu < 0 or Nv < 0.


  Transform (me : mutable; T : Trsf) ;
    	---Purpose: Applies the transformation T to this sphere.
  Copy (me)  returns mutable like me;
    	---Purpose: Creates a new object which is a copy of this sphere.
fields 

  radius : Real;


end;
