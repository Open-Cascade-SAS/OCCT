-- Created on: 1998-05-07
-- Created by: Andre LIEUTIER
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class LineConstraint from Plate
---Purpose: constraint a point to belong to a straight line
--          
--          

uses 
 XY from gp, 
 Lin  from  gp,
 LinearScalarConstraint from Plate

is
    Create(point2d : XY ; lin  :  Lin  from  gp; 
           iu : Integer = 0; iv : Integer = 0) returns LineConstraint;
-- constraint the iu th  derivative in u and iv  th derivative in v at
-- the point2d parametre to belong to the lin  line.

    -- Accessors :
    LSC(me) returns  LinearScalarConstraint ;
    ---C++: inline 
    ---C++: return const &


fields
    myLSC : LinearScalarConstraint;
    
end;

