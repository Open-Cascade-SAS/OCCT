-- Created on: 1992-09-28
-- Created by: Didier PIFFAULT
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class InterferencePolygon2d from Intf

inherits Interference from Intf

	---Purpose: Computes the  interference between two  polygons or
	--          the    self intersection of    a  polygon  in  two
	--          dimensions.

uses    Pnt2d             from gp,
    	SectionPoint      from Intf,
    	SeqOfSectionPoint from Intf,
    	TangentZone       from Intf,
    	SeqOfTangentZone  from Intf,
        Polygon2d         from Intf

raises  OutOfRange from Standard

is

-- Interface :

    Create          returns InterferencePolygon2d from Intf;
    ---Purpose: Constructs an empty interference of Polygon.


    Create         (Obje1, Obje2 : in Polygon2d) 
    	            returns InterferencePolygon2d from Intf;
    ---Purpose: Constructs and computes an interference between two Polygons.


    Create         (Obje       : in Polygon2d) 
    	            returns InterferencePolygon2d from Intf;
    ---Purpose: Constructs and computes the auto interference of a Polygon.


    Perform        (me         : in out;
    	    	    Obje1, Obje2 : in Polygon2d);
    ---Purpose: Computes an interference between two Polygons.


    Perform        (me         : in out;
    	    	    Obje       : in Polygon2d);
    ---Purpose: Computes the self interference of a Polygon.


    Pnt2dValue     (me;
    	    	    Index      : in Integer)
		    returns Pnt2d from gp
    	    	    raises OutOfRange from Standard
    	    	    is static;
    ---Purpose: Gives the  geometrical 2d point   of the  intersection
    --          point at address <Index> in the interference.


-- Implementation :

    Interference   (me : in out; Obje1, Obje2 : in Polygon2d)
    	    	    is private;

    Interference   (me : in out; Obje : in Polygon2d)
    	    	    is private;

    Clean          (me   : in out) is private;

    Intersect      (me         : in out;
                    iO, iT     : Integer from Standard;
                    BegO, EndO : in Pnt2d from gp;
                    BegT, EndT : in Pnt2d from gp)
    	    	    is private;
    ---Purpose: Computes the intersection between two segments 
    --          <BegO><EndO> et <BegT><EndT>.

fields

    oClos, tClos         : Boolean from Standard;
    nbso                 : Integer from Standard;

end InterferencePolygon2d;
