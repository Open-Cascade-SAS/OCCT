-- Created on: 1991-10-10
-- Created by: Jean Claude VAUTHIER
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class ParabolaToBSplineCurve   from Convert   inherits ConicToBSplineCurve

        --- Purpose :
        --  This algorithm converts a parabola into a non rational B-spline
        --  curve.
        --  The parabola is a Parab2d from package gp with the parametrization
        --  P (U) = Loc + F * (U*U * Xdir + 2 * U * Ydir) where Loc is the 
        --  apex of the parabola, Xdir is the normalized direction of the 
        --  symmetry axis of the parabola, Ydir is the normalized direction of
        --  the directrix and F is the focal length.
        --- KeyWords :
        --  Convert, Parabola, BSplineCurve, 2D .

uses Parab2d from gp

is


  Create (Prb : Parab2d; U1, U2 : Real)   returns ParabolaToBSplineCurve;
        --- Purpose : 
        --  The parabola Prb is limited between the parametric values U1, U2
        --  and the equivalent B-spline curve as the same orientation as the
        --  parabola Prb.


end ParabolaToBSplineCurve;
