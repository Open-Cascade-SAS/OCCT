-- Created on: 1992-08-26
-- Created by: Remi GILET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MakeHypr2d from gce inherits Root from gce

    ---Purpose :This class implements the following algorithms used to 
    --          create a 2d Hyperbola from gp.
    --          * Create a 2d Hyperbola from its center and two points:
    --            one on its axis of symmetry giving the major radius, the 
    --            other giving the value of the small radius.
    --          * Create a 2d Hyperbola from its major axis and its major
    --            radius and its minor radius.
    --            
    --
    --                         ^YAxis                
    --                         |                   
    --                  FirstConjugateBranch     
    --                         |        
    --        Other            |                Main
    --   --------------------- C ------------------------------>XAxis
    --        Branch           |                Branch
    --                         |
    --                         |         
    --                   SecondConjugateBranch
    --                         |         
    --
    --  An axis placement (one axis) is associated with the hyperbola.
    --  This axis is the "XAxis" or major axis of the hyperbola. It is
    --  the symmetry axis of the main branch of hyperbola. 
    --  The "YAxis" is normal to this axis and pass throught its location 
    --  point. It is the minor axis.
    --  
    --  The major radius is the distance between the Location point
    --  of the hyperbola C and the vertex of the Main Branch (or the
    --  Other branch). The minor radius is the distance between the
    --  Location point of the hyperbola C and the vertex of the First 
    --  (or Second) Conjugate branch.
    --  The major radius can be lower than the minor radius.

uses Pnt2d   from gp,
     Ax2d    from gp,
     Ax22d   from gp,
     Hypr2d  from gp,
     Boolean from Standard

raises NotDone from StdFail

is

Create(S1,S2  : Pnt2d from gp;
       Center : Pnt2d from gp) returns MakeHypr2d;
    ---Purpose: Constructs a hyperbola
    --   centered on the point Center, where:
    --   -   the major axis of the hyperbola is defined by Center and point S1,
    --   -   the major radius is the distance between Center and S1, and
    --   -   the minor radius is the distance between point S2 and the major axis.

Create (MajorAxis   : Ax2d    from gp      ; 
    	MajorRadius : Real    from Standard; 
    	MinorRadius : Real    from Standard;
    	Sense       : Boolean from Standard)  returns MakeHypr2d;
    --- Purpose : Constructs a hyperbola with major and minor radii MajorRadius and
    --   MinorRadius, where:
    --   -   the center of the hyperbola is the origin of the axis MajorAxis, and
    --   -   the major axis is defined by MajorAxis if Sense
    -- is true, or the opposite axis to MajorAxis if Sense is false; or
    -- -   centered on the origin of the coordinate system
    --   A, with major and minor radii MajorRadius and
    --   MinorRadius, where its major axis is the "X Axis"
    --   of A (A is the local coordinate system of the hyperbola).
 
Create (A           : Ax22d   from gp      ; 
    	MajorRadius : Real    from Standard; 
    	MinorRadius : Real    from Standard)  returns MakeHypr2d;
    --- Purpose :Creates a Hypr2d centered on the origin of the coordinate system
    --  A, with major and minor radii MajorRadius and
    --  MinorRadius, where its major axis is the "X Axis"
    --  of A (A is the local coordinate system of the hyperbola).


Value(me) returns Hypr2d from gp
    raises NotDone
    is static;
    ---C++: return const&
    ---Purpose: Returns the constructed hyperbola.
    -- Exceptions StdFail_NotDone if no hyperbola is constructed.
    
Operator(me) returns Hypr2d from gp
    is static;
    ---C++: return const&
    ---C++ : alias "Standard_EXPORT operator gp_Hypr2d() const;"

fields

    TheHypr2d : Hypr2d from gp;
    --The solution from gp.
    
end MakeHypr2d;




