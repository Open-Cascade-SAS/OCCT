-- File:	BRepExtrema_ExtPF.cdl
-- Created:	Wed Feb  9 08:33:21 1994
-- Author:	Laurent PAINNOT
--		<lpa@phylox>
---Copyright:	 Matra Datavision 1994

class ExtPF from BRepExtrema

uses
    Integer           from Standard,
    Real              from Standard,
    Boolean           from Standard,
    Face              from TopoDS,
    Vertex            from TopoDS,
    ExtPS             from Extrema,
    SequenceOfReal    from TColStd,
    SequenceOfPOnSurf from Extrema,
    Pnt               from gp,
    Surface           from BRepAdaptor
     
raises 
    NotDone      from StdFail,
    OutOfRange   from Standard,
    TypeMismatch from Standard

is
    Create returns ExtPF from BRepExtrema;

    Create(V : Vertex from TopoDS;
           E : Face   from TopoDS)
    	---Purpose: It calculates all the distances.
    returns ExtPF from BRepExtrema;

    Initialize(me: in out; E : Face from TopoDS)
    	---Purpose: 
    is static;
    
    Perform(me: in out; V : Vertex from TopoDS;
     	    	    	E : Face   from TopoDS)
    	---Purpose: An exception is raised if the fields have not been
    	--          initialized.
    	--          Be careful: this method uses the Face only for 
    	--          classify not for the fields.
    raises TypeMismatch from Standard
    is static;
    
    IsDone(me) returns Boolean from Standard
    	---Purpose: True if the distances are found.
    is static;
    
    NbExt(me) returns Integer from Standard
    	---Purpose: Returns the number of extremum distances.
    raises NotDone from StdFail
    is static;

    
    SquareDistance(me; N : Integer from Standard) returns Real from Standard
    	---Purpose: Returns the value of the <N>th extremum square distance.
    raises NotDone    from StdFail,
    	   OutOfRange from Standard
    is static;
    
    Parameter(me; N : Integer from Standard; U, V: out Real) 
    	---Purpose: Returns the parameters on the  Face  of the  <N>th
    	--          extremum distance.
    raises NotDone    from StdFail,
    	   OutOfRange from Standard
    is static;
    
    
    Point(me; N : Integer from Standard) returns Pnt from gp
    	---Purpose: Returns the Point of the <N>th extremum distance.
    raises NotDone    from StdFail, 
    	   OutOfRange from Standard
    is static;
    
    
fields
    myExtrem  : ExtPS             from Extrema;
    mynbext   : Integer           from Standard;
    mySqDist  : SequenceOfReal    from TColStd;
    myPoints  : SequenceOfPOnSurf from Extrema;
    mySurf    : Surface           from BRepAdaptor;

end ExtPF;
