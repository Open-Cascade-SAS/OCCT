-- File:        MarkerSelect.cdl
-- Created:     Fri Dec  1 11:11:11 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993



class MarkerSelect from StepVisual inherits SelectType from StepData

	-- <MarkerSelect> is an EXPRESS Select Type construct translation.
	-- it gathers : enum MarkerType

uses Transient, SelectMember from StepData, MarkerMember from StepVisual

is

	Create returns MarkerSelect;
	---Purpose : Returns a MarkerSelect SelectType

	CaseNum (me; ent : Transient) returns Integer;
	---Purpose: Recognizes a MarkerSelect Kind Entity that is :
	--        0 else

    NewMember (me) returns SelectMember from StepData  is redefined;
    ---Purpose : Returns a new MarkerMember

    CaseMem (me; sm : SelectMember from StepData) returns Integer is redefined;
    ---Purpose : Returns 1 for a SelectMember enum, named MARKER_TYPE

    MarkerMember (me) returns MarkerMember  from StepVisual;
    ---Purpose : Gives access to the MarkerMember in order to get/set its value

end MarkerSelect;
