-- Created on: 2002-12-12
-- Created by: data exchange team
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class Volume3dElementRepresentation from StepFEA
inherits ElementRepresentation from StepFEA

    ---Purpose: Representation of STEP entity Volume3dElementRepresentation

uses
    HAsciiString from TCollection,
    HArray1OfRepresentationItem from StepRepr,
    RepresentationContext from StepRepr,
    HArray1OfNodeRepresentation from StepFEA,
    FeaModel3d from StepFEA,
    Volume3dElementDescriptor from StepElement,
    ElementMaterial from StepElement

is
    Create returns Volume3dElementRepresentation from StepFEA;
	---Purpose: Empty constructor

    Init (me: mutable; aRepresentation_Name: HAsciiString from TCollection;
                       aRepresentation_Items: HArray1OfRepresentationItem from StepRepr;
                       aRepresentation_ContextOfItems: RepresentationContext from StepRepr;
                       aElementRepresentation_NodeList: HArray1OfNodeRepresentation from StepFEA;
                       aModelRef: FeaModel3d from StepFEA;
                       aElementDescriptor: Volume3dElementDescriptor from StepElement;
                       aMaterial: ElementMaterial from StepElement);
	---Purpose: Initialize all fields (own and inherited)

    ModelRef (me) returns FeaModel3d from StepFEA;
	---Purpose: Returns field ModelRef
    SetModelRef (me: mutable; ModelRef: FeaModel3d from StepFEA);
	---Purpose: Set field ModelRef

    ElementDescriptor (me) returns Volume3dElementDescriptor from StepElement;
	---Purpose: Returns field ElementDescriptor
    SetElementDescriptor (me: mutable; ElementDescriptor: Volume3dElementDescriptor from StepElement);
	---Purpose: Set field ElementDescriptor

    Material (me) returns ElementMaterial from StepElement;
	---Purpose: Returns field Material
    SetMaterial (me: mutable; Material: ElementMaterial from StepElement);
	---Purpose: Set field Material

fields
    theModelRef: FeaModel3d from StepFEA;
    theElementDescriptor: Volume3dElementDescriptor from StepElement;
    theMaterial: ElementMaterial from StepElement;

end Volume3dElementRepresentation;
