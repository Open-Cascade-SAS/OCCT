-- Created on: 1994-05-19
-- Created by: Yves FRICAUD
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package Bisector 

    --- Purpose : This package provides the bisecting line between two
    --            geometric elements.

uses 
     MMgt,
     Standard,
     TCollection,
     TColStd,	
     TColgp,
     Geom2d,
     GeomAbs,
     gp,
     math,
     IntCurve,	
     GccInt,
     StdFail,
     IntRes2d
is

    deferred class Curve;
    
   	     class BisecAna;
    	     --- Purpose: This class provides the bisecting line between two
    	     --           geometric elements.The elements are Circles,Lines or
    	     --           Points. 

    	     class BisecPC;
	     ---Purpose: This class provides the bisecting line between a point
	     --          a Curve.
    
    	     class BisecCC;	
	     ---Purpose: This class provides the bisecting line between two
	     --          Curves. 

    class Bisec;
	---Purpose: This class provides the bisecting line between two
	--          geometris  elelements.  The   bisecting   line  is
	--          trimmed by a point, 
    
    class Inter;
    
    class PointOnBis;
    
    class PolyBis;
    
    private class FunctionH;
    
    private class FunctionInter;
    
    IsConvex (Cu : Curve from Geom2d; Sign : Real) 
    returns Boolean from Standard;
    
end Bisector;
