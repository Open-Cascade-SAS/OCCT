-- Created on: 2008-07-30
-- Created by: Vladislav ROMASHKO
-- Copyright (c) 2008-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Selector from Voxel

    ---Purpose: Detects voxels in the viewer 3d under the mouse cursor.

uses

    View from V3d,
    BoolDS from Voxel,
    ColorDS from Voxel,
    ROctBoolDS from Voxel

is

    Create
    ---Purpose: An empty constructor.
    returns Selector from Voxel;
    
    Create(view : View from V3d)
    ---Purpose: A constructor of the selector,
    --          which initializes the classes
    --          by a view, where the user selects the voxels.
    returns Selector from Voxel;
    
    Init(me : in out;
    	 view : View from V3d);
    ---Purpose: Initializes the selector by a view, 
    --          where the user selects the voxels.

    SetVoxels(me : in out;
    	      voxels : BoolDS from Voxel);
    ---Purpose: Defines the voxels (1bit).

    SetVoxels(me : in out;
    	      voxels : ColorDS from Voxel);
    ---Purpose: Defines the voxels (4bit).

    SetVoxels(me : in out;
    	      voxels : ROctBoolDS from Voxel);
    ---Purpose: Defines the voxels (1bit recursive splitting).

    Detect(me : in out;
    	   winx : Integer from Standard;
	   winy : Integer from Standard;
	   ix : out Integer from Standard;
	   iy : out Integer from Standard;
	   iz : out Integer from Standard)
    ---Purpose: Detects a voxel under the mouse cursor.
    returns Boolean from Standard;

fields

    myView : View from V3d;
    myVoxels : Address from Standard;
    myIsBool : Integer from Standard; -- 0 - ColorDS, 1 - BoolDS, 2 - ROctBoolDS
    
end Selector;
