-- Created on: 1999-03-09
-- Created by: data exchange team
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DateItem from StepAP214 inherits ApprovalItem from StepAP214


uses
    	ApprovalPersonOrganization from StepBasic,
	AppliedPersonAndOrganizationAssignment from StepAP214,
    	AppliedOrganizationAssignment from StepAP214,
    	Effectivity from StepBasic

is
    Create returns DateItem;
	---Purpose : Returns a DateItem SelectType
	
	CaseNum (me; ent : Transient) returns Integer is redefined;
	---Purpose: Recognizes a DateItem Kind Entity that is :
	--        1 -> ApprovalPersonOrganization
	--        2 -> AppliedDateAndPersonAssignment
    	--        3 -> AppliedOrganizationAssignment
    	--        4 -> AssemblyComponentUsageSubstitute
	--        5 -> DocumentFile
	--        6 -> Effectivity
    	--        7 -> MaterialDesignation
    	--        8 -> MechanicalDesignGeometricPresentationRepresentation
	--        9 -> PresentationArea
    	--        10 -> Product
	--        11 -> ProductDefinition
    	--        12 -> ProductDefinitionFormation
	--        13 -> ProductDefinitionRelationship
    	--    	  14 -> PropertyDefinition
    	--        15 -> ShapeRepresentation
	--        0 else

	ApprovalPersonOrganization (me) returns any ApprovalPersonOrganization ;
	---Purpose : returns Value as a ApprovalPersonOrganization (Null if another type)

	AppliedPersonAndOrganizationAssignment (me) returns any AppliedPersonAndOrganizationAssignment ; 
	---Purpose : returns Value as a AppliedDateAndPersonAssignment (Null if another type)

    	AppliedOrganizationAssignment (me) returns any AppliedOrganizationAssignment ;
    	---Purpose : returns Value as a AppliedOrganizationAssignment (Null if another type)

	Effectivity (me) returns any Effectivity ;
	---Purpose : returns Value as a Effectivity (Null if another type)
	

end DateItem;
