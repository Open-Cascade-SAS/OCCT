-- Created on: 1997-04-17
-- Created by: Christophe MARION
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class VertexList from HLRBRep

uses
	Orientation                    from TopAbs,
        Intersection                   from HLRAlgo,
        Interference                   from HLRAlgo,
	ListIteratorOfInterferenceList from HLRAlgo,
	EdgeInterferenceTool           from HLRBRep 
is

    Create(T : EdgeInterferenceTool from HLRBRep;
           I : ListIteratorOfInterferenceList from HLRAlgo)
    returns VertexList from HLRBRep;

    IsPeriodic(me) returns Boolean from Standard
        ---Purpose: Returns True when the curve is periodic.
    is static;
    
    More(me) returns Boolean from Standard
        ---Purpose: Returns True when there are more vertices.
    is static;
    
    Next(me : in out)
        ---Purpose: Proceeds to the next vertex.
    is static;
    
    Current(me) returns Intersection from HLRAlgo
        ---Purpose: Returns the current vertex
        --          
	---C++: return const &
    is static;
    
    IsBoundary(me) returns Boolean from Standard
        ---Purpose: Returns True  if the current  vertex  is is on the
        --          boundary of the edge.
    is static;
    
    IsInterference(me) returns Boolean from Standard
        ---Purpose: Returns  True   if   the current    vertex  is  an
        --          interference. 
    is static;
    
    Orientation(me) returns Orientation from TopAbs
        ---Purpose: Returns the  orientation of the  current vertex if
        --          it is on the boundary of the edge.
    is static;
    
    Transition(me) returns Orientation from TopAbs
        ---Purpose: Returns  the transition  of the  current vertex if
        --          it is an interference.
    is static;
    
    BoundaryTransition(me) returns Orientation from TopAbs
        ---Purpose: Returns  the  transition  of  the  current  vertex
        --          relative to the boundary if it is an interference.
    is static;
    
fields
	
    myIterator   : ListIteratorOfInterferenceList from HLRAlgo;
    myTool       : EdgeInterferenceTool           from HLRBRep;
    fromEdge     : Boolean                        from Standard;
    fromInterf   : Boolean                        from Standard;

end VertexList;
