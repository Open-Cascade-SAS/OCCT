-- File:	BOPTools_PaveBlock.cdl
-- Created:	Thu Feb 15 11:21:52 2001
-- Author:	Peter KURNEV
--		<pkv@irinox>
---Copyright:	 Matra Datavision 2001


class PaveBlock from BOPTools 

	---Purpose:  
    	--  Class for storing info about a couple  
        --- of neighbouring paves on an edge  

uses
    Pave from BOPTools,  
    PointBetween from BOPTools,
    Range        from IntTools, 
    ShrunkRange  from IntTools, 
    Curve        from IntTools



is 
    Create 
    	returns PaveBlock from BOPTools;  
    	---Purpose: 
    	--- Empty constructor 
    	---
    Create (anEdge:  Integer from Standard; 
    	    aPave1:  Pave from BOPTools; 
    	    aPave2:  Pave from BOPTools); 
    	---Purpose:  
    	--- Constructor 
    	--- Index  - DS-index of the edge    	 
    	--- aPave1 - one pave              
    	--- aPave2 - other pave               
    	---
    SetEdge (me:out;   
    	     anEdge:Integer from Standard); 
    	---Purpose:  
    	--- Modifier  
    	--- Sets DS-index for the edge that is between aPave1 and aPave2 
    	---
    SetOriginalEdge  (me:out;   
    	    	      anEdge:Integer from Standard);  
    	---Purpose:  
    	--- Modifier  
    	--- Sets DS-index for the edge from which this pave block comes from 
    	---
    SetPave1(me:out;  
    	     aPave: Pave from BOPTools);	     
    	---Purpose:  
    	--- Modifier  
    	---
    SetPave2(me:out;  
    	     aPave: Pave from BOPTools);	     
    	---Purpose:  
    	--- Modifier  
    	---
    SetShrunkRange  (me:out;   
    	    	     aSR:ShrunkRange from IntTools);  
    	---Purpose:  
    	--- Modifier  
    	--- Sets the Shrunk Range for the pave block 
    	---
    SetPointBetween (me:out; 
    	    	     aP: PointBetween from BOPTools);  
    	---Purpose:  
    	--- Modifier  
    	--- Sets the point between the paves for the pave block  
    	---

    ---  Case  of  Face/Face Pave  Block 
    ---		    	     
    SetCurve        (me:out; 
    	    	     aC:Curve from IntTools);  
    	---Purpose:  
    	--- Modifier  
    	--- Sets the intersection curve to which the pave block belongs to  
    	---
    SetFace1        (me:out; 
    	    	     nF1:Integer from Standard); 
    	---Purpose:  
    	--- Modifier  
    	--- Sets the DS-index of the first face  
    	---
    SetFace2        (me:out; 
    	    	     nF2:Integer from Standard);  
    	---Purpose:  
    	--- Modifier  
    	--- Sets the DS-index of the second face  
    	---
    Edge    (me) 
    	returns Integer from Standard; 
    	---Purpose:  
    	--- Selector  
    	---
    OriginalEdge(me) 
    	returns Integer from Standard; 
    	---Purpose:  
    	--- Selector  
    	---
    Pave1(me) 
    	returns Pave from BOPTools; 
    	---C++:  return const &	 
    	---Purpose:  
    	--- Selector  
    	---
    Pave2(me) 
    	returns Pave from BOPTools; 
    	---C++:  return const &	
    	---Purpose:  
    	--- Selector  
    	---
    IsValid(me) 
	returns Boolean from Standard;	    	     
    	---Purpose:  
    	--- Returns  TRUE if both paves have vertex index !=0            
    	---
    IsEqual(me;  
    	    Other:PaveBlock from BOPTools)    
        returns Boolean from Standard;	
    	---Purpose:  
    	--- Returns  TRUE if <Other> is  equal to me 
    	---
    Parameters   (me; 
                  aT1:out Real from Standard;   
                  aT2:out Real from Standard);    
    	---Purpose:  
    	--- Returns values for paves' parameters      
    	---
    Range  (me) 
    	returns Range from IntTools; 
    	---C++:  return const &	
    	---Purpose:  
    	--- Returns parmetric range for paves' parameters      
    	---
    ShrunkRange(me) 
    	returns ShrunkRange from IntTools; 
    	---C++:  return const &  
    	---Purpose:  
    	--- Selector      
    	---
    PointBetween  (me) 
    	returns  PointBetween from BOPTools; 
    	---C++:  return const & 	 
    	---Purpose:  
    	--- Selector      
    	---
    Curve(me) 
    	returns Curve from IntTools; 
    	---C++:  return const & 
    	---Purpose:  
    	--- Selector      
    	---
    Face1(me) 
    	returns Integer from Standard; 
    	---Purpose:  
    	--- Selector      
    	---
    Face2(me) 
    	returns Integer from Standard; 
    	---Purpose:  
    	--- Selector      
    	---
    IsInBlock(me; 
    	   aPaveX:  Pave from BOPTools) 
    	returns Boolean  from Standard;  
    
fields   

    myEdge         :  Integer from Standard;
    myOriginalEdge :  Integer from Standard;
    myPave1        :  Pave from BOPTools; 
    myPave2        :  Pave from BOPTools; 
    myRange        :  Range from IntTools;     
    myShrunkRange  :  ShrunkRange from IntTools; 
    myCurve        :  Curve from IntTools; 
    myFace1        :  Integer from Standard; 
    myFace2        :  Integer from Standard; 
    myPointBetween :  PointBetween from BOPTools;  
     
end PaveBlock;
