-- Created on: 1992-10-21
-- Created by: Christian CAILLET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



deferred class SingleParentEntity  from IGESData  inherits IGESEntity

    ---Purpose : a SingleParentEntity is a kind of IGESEntity which can refer
    --           to a (Single) Parent, from Associativities list of an Entity
    --           a effective SingleParent definition entity must inherit it

uses Integer

raises OutOfRange

is

    SingleParent (me) returns IGESEntity  is deferred;
    ---Purpose : Returns the parent designated by the Entity, if only one !

    NbChildren (me) returns Integer  is deferred;
    ---Purpose : Returns the count of Entities designated as children

    Child (me; num : Integer) returns IGESEntity
    ---Purpose : Returns a Child given its rank
    	raises OutOfRange  is deferred;
    --           Error if <num> is below one or over <NbChildren>

end SingleParentEntity;
