-- Created on: 1993-04-23
-- Created by: Laurent BUCHARD
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package ApproxInt

uses 
     Standard,TCollection,math,gp,TColStd,TColgp,
     IntImp,IntSurf,
     AppParCurves,StdFail,Approx,MMgt
     
is

    deferred class SvSurfaces;     
    generic class PrmPrmSvSurfaces,TheInt2S;
    generic class ImpPrmSvSurfaces,TheZerImpFunc;
    generic class MultiLine;
    generic class MultiLineTool;
    generic class Approx,ThePrmPrmSvSurfaces,
                         TheImpPrmSvSurfaces,
                         TheMultiLine,
                         TheMultiLineTool,
			 TheComputeLine,
                         TheComputeLineBezier;

end ApproxInt;
