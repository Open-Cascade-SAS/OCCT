-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class OrientedClosedShell from StepShape 

inherits ClosedShell from StepShape 

uses

	Boolean from Standard, 
	HArray1OfFace from StepShape, 
	Face from StepShape, 
	HAsciiString from TCollection
is

	Create returns OrientedClosedShell;
	---Purpose: Returns a OrientedClosedShell


	Init (me : mutable;
	      aName : HAsciiString from TCollection;
	      aCfsFaces : HArray1OfFace from StepShape) is redefined;

	Init (me : mutable;
	      aName : HAsciiString from TCollection;
	      aClosedShellElement : ClosedShell from StepShape;
	      aOrientation : Boolean from Standard) is virtual;

	-- Specific Methods for Field Data Access --

	SetClosedShellElement(me : mutable; aClosedShellElement : ClosedShell);
	ClosedShellElement (me) returns ClosedShell;
	SetOrientation(me : mutable; aOrientation : Boolean);
	Orientation (me) returns Boolean;
	SetCfsFaces(me : mutable; aCfsFaces : HArray1OfFace) is redefined;
	CfsFaces (me) returns HArray1OfFace is redefined;
	CfsFacesValue (me; num : Integer) returns Face is redefined;
	NbCfsFaces (me) returns Integer is redefined;

fields

	closedShellElement : ClosedShell from StepShape;
	orientation : Boolean from Standard;

 -- 
 -- NB : field <cfs_faces> inherited from classe <connected_face_set> is redeclared.
 --      it shall appears in a physical file as a *.
 --

end OrientedClosedShell;
