-- Created on: 1993-03-23
-- Created by: BBL,JLF
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


deferred class AlienImage from AlienImage inherits TShared from MMgt

	---Purpose: This class defines an Alien image.
	-- Alien Image is X11 .xwd image or SGI .rgb image for example

uses
	File  		from OSD,
	Image 		from Image

raises
	TypeMismatch 	from Standard

is
	Initialize ;

	Read ( me : in out mutable ; afile : in out File from OSD )
	  returns Boolean from Standard is deferred;
	---Level: Public
	---Purpose: Reads content of a  AlienImage object from a file .
	--         Returns True if file is a XWD file .

	Write( me : in immutable ; afile : in out File from OSD )
	  returns Boolean from Standard is deferred ;
	---Level: Public
	---Purpose: Writes content of a  AlienImage object to a file .

	ToImage  ( me : in immutable ) 
	  returns mutable Image from Image 
          raises TypeMismatch from Standard is deferred ;
	---Level: Public
	---Purpose : Converts a AlienImage object to a Image object.

	FromImage( me : in out mutable ; anImage : in Image from Image )
          raises TypeMismatch from Standard is deferred ;
	---Level: Public
	---Purpose : Converts a Image object to a AlienImage object.

end AlienImage;
 
