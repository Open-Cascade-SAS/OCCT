-- Created on: 1993-02-05
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package Contap

	---Purpose: 

uses Standard,StdFail,MMgt, GeomAbs, TopAbs, TCollection, gp, TColgp,
     math, IntSurf, IntStart, IntWalk,
     Geom2d, TColStd, Geom, Adaptor3d,  Adaptor2d

is

    deferred generic class ArcTool;        -- template class
    
    deferred generic class SurfaceTool;    -- template class
    
    deferred generic class TopolTool;      -- template class
    
    generic class Point;

    generic class Line;

    generic class SurfFunction;
    
    generic class ArcFunction;
    
    generic class SurfProps;

    generic class ContourGen, ThePoint,TheSequenceOfPoint,TheHSequenceOfPoint,
                              TheLine, TheSequenceOfLine,
			      TheSurfProps, TheSurfFunction, TheArcFunction,
                              TheSearch, TheIWalking, TheSearchInside;
    	    	    	      ---TheLineConstructor;

    class ContAna;		   

    enumeration TFunction is
    	ContourStd,
	ContourPrs,
	DraftStd,
	DraftPrs
    end TFunction;	

    enumeration IType is  -- a replacer dans IntSurf et fusionner avec IntPatch
    -- type of the line of contour

    	Lin,       -- pour conflit avec deferred class Line
    	Circle,
        Walking,
    	Restriction
    end IType;
	
    generic class HContToolGen;
    
    generic class HCurve2dToolGen;
    
    class HCurve2dTool instantiates 
    	HCurve2dToolGen from Contap ( 
	    HCurve2d from Adaptor2d);

    class HContTool instantiates 
        HContToolGen from Contap (
    	 HVertex       from Adaptor3d,
	 HCurve2d      from Adaptor2d,
	 HSurface      from Adaptor3d,
    	 HCurve2dTool  from Contap,
	 HSurfaceTool  from Adaptor3d);
	 
    class Contour instantiates ContourGen from Contap
    	(HVertex       from Adaptor3d,
	 HCurve2d      from Adaptor2d,
	 HSurface      from Adaptor3d,
	 HCurve2dTool  from Contap,
	 HSurfaceTool  from Adaptor3d,
	 HContTool     from Contap,
	 TopolTool     from Adaptor3d);


end Contap;
