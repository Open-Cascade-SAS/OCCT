-- File:        CameraModel.cdl
-- Created:     Mon Dec  4 12:02:24 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWCameraModel from RWStepVisual

	---Purpose : Read & Write Module for CameraModel

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     CameraModel from StepVisual

is

	Create returns RWCameraModel;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable CameraModel from StepVisual);

	WriteStep (me; SW : in out StepWriter; ent : CameraModel from StepVisual);

end RWCameraModel;
