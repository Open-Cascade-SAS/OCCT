-- File:      HLRAppli.cdl
-- Created:   05.12.12 15:50:05
-- Created by: Julia GERASIMOVA
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package HLRAppli

        ---Purpose : This package represents applications
        --           of Hidden Lines Removal algorithm

uses
    TopoDS,
    HLRAlgo

is
    class ReflectLines;
    
end HLRAppli;
