-- Created on: 1997-03-26
-- Created by: Christian CAILLET
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class PresentationLayerUsage  from StepVisual    inherits TShared

    ---Purpose : Added from StepVisual Rev2 to Rev4

uses
     PresentationLayerAssignment from StepVisual,
     PresentationRepresentation from StepVisual

is

    Create returns PresentationLayerUsage;

    Init (me : mutable;
    	  aAssignment : PresentationLayerAssignment from StepVisual;
	  aPresentation : PresentationRepresentation from StepVisual);

    SetAssignment (me : mutable; aAssignment : PresentationLayerAssignment from StepVisual);
    Assignment (me) returns PresentationLayerAssignment from StepVisual;

    SetPresentation (me : mutable; aPresentation : PresentationRepresentation from StepVisual);
    Presentation (me) returns PresentationRepresentation from StepVisual;

fields

    theAssignment : PresentationLayerAssignment from StepVisual;
    thePresentation : PresentationRepresentation from StepVisual;

end PresentationLayerUsage;
