-- Created on: 1992-09-22
-- Created by: Christian CAILLET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package IFGraph

    	---Purpose : Provides tools to operate on an InterfaceModel and its
    	--           Entities as on a Graph. These Tools are based on classes
    	--           Graph and GraphContent  from Interface

uses Interface, GraphTools, TColStd, Standard

is

--  (sub-classes of GraphContent from Interface)
    	class AllShared;
	class AllConnected;
    	class Cumulate;
    	class Compare;
	class ExternalSources;

    	class Articulations;

    class SubPartsIterator;  -- result as several subsets
    	class ConnectedComponants;
    	class StrongComponants;
	class Cycles;
	class SCRoots;

--    class SortedStrongsFrom  instantiates  SortedStrgCmptsFromIterator from GraphTools
--    	(Graph from Interface,Transient,
--    	 MapTransientHasher from TColStd,GraphContent from Interface);

--    class SortedStrongs instantiates SortedStrgCmptsIterator from GraphTools
--    	(Graph from Interface,Transient,
--    	 GraphContent from Interface,SortedStrongsFrom from IFGraph);

--    class SortedStrongs instantiates SortedStrgCmptsIterator
--    	(Graph,Transient,GraphContent,GraphContent);

end IFGraph;
