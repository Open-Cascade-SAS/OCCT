-- Created on: 2000-04-18
-- Created by: Andrey BETENEV
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0

class DimensionalLocationWithPath from StepShape
inherits DimensionalLocation from StepShape

    ---Purpose: Representation of STEP entity DimensionalLocationWithPath

uses
    HAsciiString from TCollection,
    ShapeAspect from StepRepr

is
    Create returns DimensionalLocationWithPath from StepShape;
	---Purpose: Empty constructor

    Init (me: mutable; aShapeAspectRelationship_Name: HAsciiString from TCollection;
                       hasShapeAspectRelationship_Description: Boolean;
                       aShapeAspectRelationship_Description: HAsciiString from TCollection;
                       aShapeAspectRelationship_RelatingShapeAspect: ShapeAspect from StepRepr;
                       aShapeAspectRelationship_RelatedShapeAspect: ShapeAspect from StepRepr;
                       aPath: ShapeAspect from StepRepr);
	---Purpose: Initialize all fields (own and inherited)

    Path (me) returns ShapeAspect from StepRepr;
	---Purpose: Returns field Path
    SetPath (me: mutable; Path: ShapeAspect from StepRepr);
	---Purpose: Set field Path

fields
    thePath: ShapeAspect from StepRepr;

end DimensionalLocationWithPath;
