-- Created on: 1994-09-02
-- Created by: Yves FRICAUD
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class CurAndInf from LProp 

	---Purpose: Stores the parameters of a curve 2d or 3d corresponding
	--          to the curvature's extremas and the Inflection's Points.

uses
    CIType            from LProp,
    SequenceOfReal    from TColStd,
    SequenceOfCIType  from LProp
    
raises 
    OutOfRange from Standard 
    
is
    Create;
    
    AddInflection (me : in out; Param : Real) 
    is static;
    
    AddExtCur (me : in out; Param : Real; IsMin : Boolean)
    is static;
    
    Clear (me : in out) 
    is static;
    
    IsEmpty (me) returns Boolean
    is static;
    
    NbPoints (me) returns Integer
	---Purpose: Returns the number of points.
	--          The Points are stored to increasing parameter.
    is static;
    
    Parameter (me; N : Integer) returns Real
	---Purpose: Returns the parameter of the Nth point.
    raises
    	OutOfRange from Standard
	---Purpose: raises if N not in the range [1,NbPoints()]    
    is static;
    
    Type (me; N : Integer) returns CIType 
    	---Purpose: Returns 
    	--          - MinCur if the Nth parameter corresponds to
    	--          a minimum of the radius of curvature.
    	--          - MaxCur if the Nth parameter corresponds to
    	--          a maximum of the radius of curvature.    
    	--          - Inflection if the parameter corresponds to
    	--          a point of inflection.
    raises
    	OutOfRange from Standard
	---Purpose: raises if N not in the range [1,NbPoints()] 
    is static;	    
    
fields
    theParams : SequenceOfReal    from TColStd;
    theTypes  : SequenceOfCIType  from LProp;

end CurAndInf;


