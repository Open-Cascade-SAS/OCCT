-- Created on: 1995-06-14
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class FaceEdgeFiller from TopOpeBRep

uses

    Shape                      from TopoDS,
    FaceEdgeIntersector              from TopOpeBRep,
    HDataStructure                   from TopOpeBRepDS,
    DataStructure                               from TopOpeBRepDS,
    Interference                     from TopOpeBRepDS,
    ListOfInterference               from TopOpeBRepDS,    
    ListIteratorOfListOfInterference from TopOpeBRepDS,
    Point                            from TopOpeBRepDS
    
is 

    Create returns FaceEdgeFiller from TopOpeBRep;
    
    Insert(me : in out;
    	   F,E : Shape from TopoDS;
    	   FEINT : in out FaceEdgeIntersector from TopOpeBRep;
	   HDS : HDataStructure from TopOpeBRepDS)
    is static;

    -- -------
    -- private
    -- -------

    ScanInterfList(me; 
    	IT : in out ListIteratorOfListOfInterference from TopOpeBRepDS;
	DSP : Point from TopOpeBRepDS;
	BDS : DataStructure from TopOpeBRepDS)
    ---Purpose: 
    -- Search, among a list of interferences accessed by the iterator
    -- <IT>, a geometry <G> whose 3D point is identical to the 3D point
    -- of the TheDSPoint <DSP>.
    -- returns True if such an interference has been found, False else.
    -- if True, iterator It points (by the Value() method) on the first 
    -- interference accessing an identical 3D point.
	
    returns Boolean from Standard
    is static private;

    GetGeometry(me ; 
         IT : in out ListIteratorOfListOfInterference from TopOpeBRepDS;
	 EI : FaceEdgeIntersector from TopOpeBRep;
	 G  : in out Integer from Standard;
    	 DS : DataStructure from TopOpeBRepDS)
    ---Purpose:
    -- Search for an interference in list <IT> which 3D geometry 
    -- equals 3D geometry of the current intersection of <EI>.
    -- The search is performed by ScanInterfList.
    -- if found, set <G> to the geometry of the interference found.
    -- returns found.
	
    returns Boolean from Standard
    is static private;

    MakeGeometry(me ; EI : in out FaceEdgeIntersector from TopOpeBRep;
    	    	      DS  : in out DataStructure from TopOpeBRepDS)
    returns Integer from Standard
    is static private;

    GetGeometry(me ; L   : ListOfInterference from TopOpeBRepDS;
		     DSP : Point from TopOpeBRepDS;
		     G   : in out Integer from Standard;
    	    	     DS  : in out DataStructure from TopOpeBRepDS)
    ---Purpose:
    -- Get the geometry of a DS point <DSP>.
    -- First, search it with ScanInterfList (previous method).
    -- if found, set <G> to the geometry of the interference found.
    -- else, add the point <DSP> in the <DS> and set <G> to the 
    -- value of the new geometry such created.
    -- 
    -- returns the value of ScanInterfList().
	
    returns Boolean from Standard
    is static private;


    StoreInterference(me; 
    	    	      I   : Interference from TopOpeBRepDS;
    	    	      LI  : in out ListOfInterference from TopOpeBRepDS;
		      BDS : in out DataStructure from TopOpeBRepDS)
    ---Purpose: 
    -- Add interference <I> to list <LI>.
    -- Add <I> to the interference list of <I> geometry (via <BDS>).
    is static private;
        
end FaceEdgeFiller from TopOpeBRep;
