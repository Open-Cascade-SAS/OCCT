-- File:	TFunction_DriverTable.cdl
-- Created:	Fri Jun 11 17:25:03 1999
-- Author:	Vladislav ROMASHKO
--		<vro@flox.nnov.matra-dtv.fr>
---Copyright:	 Matra Datavision 1999

class DriverTable from TFunction inherits TShared from MMgt
    	---Purpose: A container for instances of drivers.
    	-- You create a new instance of TFunction_Driver
    	-- and use the method AddDriver to load it into the driver table.
uses 
 
    DataMapOfGUIDDriver from TFunction, 
    Driver              from TFunction, 
    GUID                from Standard, 
    OStream             from Standard,
    DataMapOfGUIDDriver from TFunction,
    HArray1OfDataMapOfGUIDDriver from TFunction
    
is 

    Get (myclass)
    ---Purpose: Returns the driver table. If a driver does not exist, creates it.
    returns mutable DriverTable from TFunction;

    Create returns mutable DriverTable from TFunction; 
    ---Purpose: Default constructor

    AddDriver(me : mutable; guid   : GUID    from Standard;
    	    	    	    driver : Driver  from TFunction;
    	    	    	    thread : Integer from Standard = 0)
    ---Purpose: Returns true if the driver has been added successfully to the driver table.
    returns Boolean from Standard;

    HasDriver (me; guid   : GUID    from Standard;
    	    	   thread : Integer from Standard = 0)
    ---Purpose: Returns true if the driver exists in the driver table.
    returns Boolean from Standard;

    FindDriver(me; guid   :     GUID   from Standard; 
	 	   driver : out Driver from TFunction;
    	    	   thread :     Integer from Standard = 0)  
    ---Purpose: Returns true if the driver was found.
    returns Boolean from Standard;

    Dump(me; anOS : in out OStream from Standard) 
    ---C++: alias operator << 
    ---C++: return &
    returns OStream from Standard;

    RemoveDriver (me : mutable; guid   : GUID    from Standard;
    	    	    	    	thread : Integer from Standard = 0)
    ---Purpose: Removes a driver with the given GUID.
    --     Returns true if the driver has been removed successfully.
    returns Boolean from Standard;

    Clear (me : mutable);
    ---Purpose: Removes all drivers. Returns true if the driver has been removed successfully.

fields

    myDrivers       : DataMapOfGUIDDriver          from TFunction;
    myThreadDrivers : HArray1OfDataMapOfGUIDDriver from TFunction;

end DriverTable;   
