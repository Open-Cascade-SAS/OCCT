-- Created on: 1994-09-21
-- Created by: Christian CAILLET
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package APIHeaderSection

    ---Purpose : This package gives the means to access to the Header of a
    --           Step Model

uses  Standard, TCollection, Interface, IFSelect, StepData, HeaderSection

is

    class MakeHeader;  -- which provide basic access services to Step Header

    class EditHeader;  -- to edit a Step Header

end APIHeaderSection;
