-- File:        FaceBound.cdl
-- Created:     Fri Dec  1 11:11:20 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class FaceBound from StepShape 

inherits TopologicalRepresentationItem from StepShape 

uses

	Loop from StepShape, 
	Boolean from Standard, 
	HAsciiString from TCollection
is

	Create returns mutable FaceBound;
	---Purpose: Returns a FaceBound


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aBound : mutable Loop from StepShape;
	      aOrientation : Boolean from Standard) is virtual;

	-- Specific Methods for Field Data Access --

	SetBound(me : mutable; aBound : mutable Loop);
	Bound (me) returns mutable Loop;
	SetOrientation(me : mutable; aOrientation : Boolean);
	Orientation (me) returns Boolean;

fields

	bound : Loop from StepShape;
	orientation : Boolean from Standard;

end FaceBound;
