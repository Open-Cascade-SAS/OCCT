-- Created on: 1993-01-09
-- Created by: CKY / Contract Toubro-Larsen ( TCD )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DrawingUnits from IGESGraph  inherits IGESEntity

        ---Purpose: defines IGESDrawingUnits, Type <406> Form <17>
        --          in package IGESGraph
        --
        --          Specifies the drawing space units as outlined
        --          in the Drawing entity

uses

        HAsciiString from TCollection

is

        Create returns DrawingUnits;

        -- Specific Methods pertaining to the class

        Init (me      : mutable;
              nbProps : Integer;
              aFlag   : Integer;
              aUnit   : HAsciiString from TCollection);
        ---Purpose : This method is used to set the fields of the class
        --           DrawingUnits
        --      - nbProps : Number of property values (NP = 2)
        --      - aFlag   : DrawingUnits Flag
        --      - aUnit   : DrawingUnits Name

        NbPropertyValues  (me) returns Integer;
        ---Purpose : returns the number of property values in <me>

        Flag (me) returns Integer;
        ---Purpose : returns the drawing space units of <me>

        Unit (me) returns HAsciiString from TCollection;
        ---Purpose : returns the name of the drawing space units of <me>

    	    --  additionnal information, deducted from Flag

    	UnitValue (me) returns Real;
	---Purpose : Computes the value of the unit, in meters, according Flag
	--           (same values as for GlobalSection from IGESData)

fields

--
-- Class    : IGESGraph_DrawingUnits
--
-- Purpose  : Declaration of the variables specific to a Drawing Unit.
--
-- Reminder : A Drawing Unit is defined by :
--                  - Number of property values (NP = 2)
--                  - Units Flag
--                  - Units Name
--

        theNbPropertyValues : Integer;

        theFlag             : Integer;

        theUnit             : HAsciiString from TCollection;

end DrawingUnits;
