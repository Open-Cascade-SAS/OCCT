-- File:	StepRepr_QuantifiedAssemblyComponentUsage.cdl
-- Created:	Mon Jul  3 20:13:37 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class QuantifiedAssemblyComponentUsage from StepRepr
inherits AssemblyComponentUsage from StepRepr

    ---Purpose: Representation of STEP entity QuantifiedAssemblyComponentUsage

uses
    HAsciiString from TCollection,
    ProductDefinition from StepBasic,
    MeasureWithUnit from StepBasic

is
    Create returns QuantifiedAssemblyComponentUsage from StepRepr;
	---Purpose: Empty constructor

    Init (me: mutable; aProductDefinitionRelationship_Id: HAsciiString from TCollection;
                       aProductDefinitionRelationship_Name: HAsciiString from TCollection;
                       hasProductDefinitionRelationship_Description: Boolean;
                       aProductDefinitionRelationship_Description: HAsciiString from TCollection;
                       aProductDefinitionRelationship_RelatingProductDefinition: ProductDefinition from StepBasic;
                       aProductDefinitionRelationship_RelatedProductDefinition: ProductDefinition from StepBasic;
                       hasAssemblyComponentUsage_ReferenceDesignator: Boolean;
                       aAssemblyComponentUsage_ReferenceDesignator: HAsciiString from TCollection;
                       aQuantity: MeasureWithUnit from StepBasic);
	---Purpose: Initialize all fields (own and inherited)

    Quantity (me) returns MeasureWithUnit from StepBasic;
	---Purpose: Returns field Quantity
    SetQuantity (me: mutable; Quantity: MeasureWithUnit from StepBasic);
	---Purpose: Set field Quantity

fields
    theQuantity: MeasureWithUnit from StepBasic;

end QuantifiedAssemblyComponentUsage;
