-- Created on: 1992-11-25
-- Created by: Jean Pierre TIRAULT
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class Array2Descriptor from TCollection

uses 
    Integer from Standard,
    Address from Standard

is
    Initialize (aLowerRow: Integer; aUpperRow: Integer; 
    	    	aLowerCol: Integer; aUpperCol: Integer;
    	    	anAddress: Address);

    UpperRow (me) returns Integer;
    ---Level: Advanced
    
    LowerRow (me) returns Integer;
    ---Level: Advanced

    UpperCol (me) returns Integer;
    ---Level: Advanced
    
    LowerCol (me) returns Integer;
    ---Level: Advanced

    Address(me) returns Address;
    ---Level: Advanced

fields
    myAddress     : Address;
    myLowerRow    : Integer;
    myLowerCol    : Integer;
    myUpperRow    : Integer;
    myUpperCol    : Integer;

    
end;    
