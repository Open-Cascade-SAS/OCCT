-- Created on: 1991-05-14
-- Created by: Annick PANCHER
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Revised:     Mireille MERCIEN


deferred generic class Compare from TCollection ( Item as any )

	---Purpose: Defines a comparison operator which can be used by
	-- any ordered structure.   The  way to compare items
	-- has  to be described  in  subclasses, which inherit
	-- from instantiations of Compare.

is

    IsLower (me; Left, Right: Item)
	---Level: Public
	---Purpose: returns True if <Left> is lower than <Right>.
    returns Boolean
    is virtual;
    
    IsGreater (me; Left, Right: Item)
	---Level: Public
	---Purpose: returns True if <Left> is greater than <Right>.
    returns Boolean
    is virtual;

    IsEqual(me; Left, Right: Item)
	---Level: Public
	---Purpose: returns True when <Right> and <Left> are equal.
    returns Boolean
    is virtual;
	
end;


