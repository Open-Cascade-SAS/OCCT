-- Created on: 1993-12-23
-- Created by: Gilles DEBARBOUILLE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


generic class FuzzyInstance from Dynamic (Dictionary as Transient)

inherits

    FuzzyClass from Dynamic

	---Purpose: This class  describes the  facilities available to
	--          manipulate fuzzy  objects. It  is a  generic class
	--          because the creation of a FuzzyInstance requests a
	--          specific dictionary of definitions.

uses

    CString from Standard,
    Integer from Standard,
    Real    from Standard,
    Boolean from Standard,
    OStream from Standard,
    FuzzyDefinition from Dynamic,
    Parameter       from Dynamic,
    AsciiString     from TCollection

is

    Create(atype : CString from Standard) returns mutable FuzzyInstance from Dynamic;
    --- Purpose: Creates  a   FuzzyInstance    object  of   the   type
    --  <atype>. If  <atype>  is not defined  in the   dictionary, the
    --  object created will have no definition.

    Create(afuzzyinstance : FuzzyInstance from Dynamic) returns mutable FuzzyInstance from Dynamic;
    --- Purpose: Creates a  FuzzyInstance with as definition the fuzzy
    --           instance <afuzzyinstance>.

    Type(me) returns AsciiString from TCollection is redefined;
    ---Purpose: Returns the type of object read in the definition.
    
    Definition(me) returns FuzzyClass from Dynamic is static;
    ---Purpose: Returns   a    reference to  the   definition   of the
    --          FuzzyInstance.
    
    Parameter(me : mutable ; aparameter : CString from Standard; avalue : Boolean from Standard) is redefined;
    ---Purpose: Adds to the  instance <me> the parameter  <aparameter>
    --          with the boolean value <avalue>.
    
    Parameter(me : mutable ; aparameter : CString from Standard; avalue : Integer from Standard) is redefined;
    ---Purpose: Adds  to the instance <me>  the parameter <aparameter>
    --          with the integer value <avalue>.
    
    Parameter(me : mutable ; aparameter : CString from Standard ; avalue : Real from Standard) is redefined;
    ---Purpose: Adds  to the  instance  <me>  the parameter <aparameter>
    --          with the real value <avalue>.
    
    Parameter(me : mutable ; aparameter : CString from Standard; astring : CString from Standard) is redefined;
    ---Purpose: Adds  to the  instance  <me>  the parameter <aparameter>
    --          with the string <astring>.
    
    Parameter(me : mutable ; aparameter : CString from Standard ; anobject : any Transient) is redefined;
    ---Purpose: Adds  to the  instance  <me>  the parameter <aparameter>
    --          with the object value <anobject>.
    
    Value(me ; aparameter : CString from Standard ; avalue : out Boolean from Standard)  
    returns Boolean from Standard is redefined;   
    ---Purpose: Returns True, if   there is a parameter   <aparameter>
    --          previously  stored in the  instance <me>  and there is
    --          the corresponding boolean value in the output argument
    --          <avalue>, False otherwise.
     
    Value(me ; aparameter : CString from Standard ; avalue : out Integer from Standard)  
    returns Boolean from Standard is redefined;    
    ---Purpose: Returns True,  if  there  is a  parameter <aparameter>
    --          previously stored  in the instance   <me> and there is
    --          the corresponding integer value in the output argument
    --          <avalue>, False otherwise.
    
    Value(me ; aparameter : CString from Standard ; avalue : out Real from Standard)  
    returns Boolean from Standard is redefined;   
    ---Purpose: Returns  True,  if there is  a  parameter <aparameter>
    --          previously  stored in the instance  <me>  and there is
    --          the corresponding real  value  in the output  argument
    --          <avalue>, False otherwise.
    
    Value(me ; aparameter : CString from Standard ; avalue : out AsciiString from TCollection)  
    returns Boolean from Standard is redefined; 
    ---Purpose: Returns True,  if  there is  a parameter  <aparameter>
    --          previously  stored in the instance   <me> and there is
    --          the   corresponding string   in  the  output  argument
    --          <avalue>, False otherwise.
    
    Value(me ; aparameter : CString from Standard ; avalue : out any Transient)  
    returns Boolean from Standard is redefined;   
    ---Purpose: Returns  True,  if  there is  a   parameter <aparameter>
    --          previously stored  in the instance <me> and   there is
    --          the corresponding object value  in  the output argument
    --          <avalue>, False otherwise.
    
    Dump(me ; astream : in out OStream from Standard) is redefined;
    ---Purpose: Useful for debugging.
    
fields

    thedefinition : FuzzyClass from Dynamic;

end FuzzyInstance;
