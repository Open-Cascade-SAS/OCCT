-- Created on: 1993-04-07
-- Created by: Laurent BUCHARD
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class IntersectionPoint from IntCurveSurface

    ---Purpose: Definition of an interserction point between a 
    --          curve and a surface. 

    ---Level: Public

   
uses
    Pnt                   from gp,
    TransitionOnCurve     from IntCurveSurface

is 

    Create
    	---Purpose: Empty Constructor.
    	returns IntersectionPoint from IntCurveSurface;
	
    Create(P     : Pnt        from gp; 
    	   USurf : Real       from Standard;
	   VSurf : Real       from Standard;
	   UCurv : Real       from Standard;
	   TrCurv: TransitionOnCurve   from IntCurveSurface)
	---Purpose: Create an IntersectionPoint.
	returns IntersectionPoint from IntCurveSurface;
	
    SetValues(me: in out;
             P     : Pnt        from gp; 
      	     USurf : Real       from Standard;
	     VSurf : Real       from Standard;
	     UCurv : Real       from Standard;
	     TrCurv: TransitionOnCurve   from IntCurveSurface)
	 ---Purpose: Set the fields of the current IntersectionPoint.
	 is static;
	 
    Values(me;
    	  P     : out Pnt        from gp; 
    	  USurf : out Real       from Standard;
	  VSurf : out Real       from Standard;
	  UCurv : out Real       from Standard;
	  TrCurv: out TransitionOnCurve   from IntCurveSurface)
	 ---Purpose: Get the fields of the current IntersectionPoint.
	 is static;
	 
    Pnt(me)
    	 ---Purpose: returns the geometric point.
         ---C++: return const & 
         ---C++: inline
         returns Pnt from gp
         is static;

    U(me)
    	 ---Purpose: returns the U parameter on the surface.
         ---C++: inline
         returns Real from Standard
         is static;

    V(me)
    	 ---Purpose: returns the V parameter on the surface.
         ---C++: inline
         returns Real from Standard
         is static;

    W(me)
    	 ---Purpose: returns the parameter on the curve.
         ---C++: inline
         returns Real from Standard
         is static;

    Transition(me)
    	 ---Purpose: returns the Transition of the point.
         ---C++: inline
         returns TransitionOnCurve from IntCurveSurface
         is static;


    Dump(me) 
    	 ---Purpose: Dump all the fields.
    	 is static;

fields

    myP       : Pnt      from gp;
    myUSurf   : Real     from Standard;
    myVSurf   : Real     from Standard;
    myUCurv   : Real     from Standard;
    myTrOnCurv: TransitionOnCurve   from IntCurveSurface;
 
end IntersectionPoint;

