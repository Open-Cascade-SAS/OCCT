-- Created on: 1995-01-27
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package GeomInt

	---Purpose: Provides intersections on between two surfaces of Geom.
	--          The result are curves from Geom.


uses StdFail,
     TCollection,
     TColStd,
     TopAbs,
     
     gp,
     Geom,
     Geom2d,
     TColGeom,
     TColGeom2d,     
     Adaptor3d,
     GeomAdaptor,

     IntSurf,
     IntPatch,
     ApproxInt,
     Bnd

is

    class IntSS;
    imported VectorOfReal;

    class LineConstructor;

    class LineTool;

    class WLApprox instantiates Approx from ApproxInt
    	(HSurface     from Adaptor3d,
	 HSurfaceTool from Adaptor3d,
	 Quadric      from IntSurf,
	 QuadricTool  from IntSurf,
	 WLine        from IntPatch);
	 
    private class ParameterAndOrientation;

    imported SequenceOfParameterAndOrientation;

    AdjustPeriodic(thePar    : Real from Standard;
            	   theParMin : Real from Standard;
            	   theParMax : Real from Standard;
            	   thePeriod : Real from Standard;
            	   theNewPar : out Real from Standard;
            	   theOffset : out Real from Standard;
            	   theEps    : Real from Standard = 0.0)
    returns Boolean from Standard;        
    ---Purpose:  Adjusts the parameter <thePar> to the range [theParMin,  theParMax]

end GeomInt;
