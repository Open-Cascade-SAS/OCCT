-- Created on: 1995-04-20
-- Created by: Christian CAILLET
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Activator  from StepSelect  inherits Activator  from IFSelect

    ---Purpose : Performs Actions specific to StepSelect, i.e. creation of
    --           Step Selections and Counters, plus dumping specific to Step

uses CString, SessionPilot, ReturnStatus

is

    Create returns mutable Activator from StepSelect;


    Do   (me : mutable; number : Integer; pilot : mutable SessionPilot)
    	returns ReturnStatus;
    ---Purpose : Executes a Command Line for StepSelect

    Help (me; number : Integer) returns CString;
    ---Purpose : Sends a short help message for StepSelect commands

end Activator;
