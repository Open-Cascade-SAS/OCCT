-- Created on: 1993-01-09
-- Created by: CKY / Contract Toubro-Larsen ( TCD )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DefinitionLevel from IGESGraph  inherits LevelListEntity

        ---Purpose: defines IGESDefinitionLevel, Type <406> Form <1>
        --          in package IGESGraph
        --
        --          Indicates the no. of levels on which an entity is
        --          defined

uses

        IGESEntity       from IGESData,
        HArray1OfInteger from TColStd

raises OutOfRange

is

        Create returns mutable DefinitionLevel;

        -- Specific Methods pertaining to the class

        Init (me              : mutable;
              allLevelNumbers : HArray1OfInteger);
        ---Purpose : This method is used to set the fields of the class
        --           DefinitionLevel
        --       - allLevelNumbers : Values of Level Numbers

        NbPropertyValues (me) returns Integer;
        ---Purpose : returns the number of property values in <me>

        NbLevelNumbers (me) returns Integer;
        ---Purpose : Must return the count of levels (== NbPropertyValues)

        LevelNumber (me; LevelIndex : Integer) returns Integer
        raises OutOfRange;
        ---Purpose : returns the Level Number of <me> indicated by <LevelIndex>
        -- raises an exception if LevelIndex is <= 0 or
        -- LevelIndex > NbPropertyValues

fields

--
-- Class    : IGESGraph_DefinitionLevel
--
-- Purpose  : Declaration of the variables specific to a Definition Level.
--
-- Reminder : A Definition Level is defined by :
--              - Level Numbers

        theLevelNumbers : HArray1OfInteger;

end DefinitionLevel;
