--
-- File:	Aspect_LineStyle.cdl
-- Created:	Mardi 7 Septembre 1993
-- Author:	GG
-- Updated:	JLF (Reason LineStyle MUST be given in METER ) 2 Mars 94
--
---Copyright:	MatraDatavision 1991-1993
--

class LineStyle from Aspect

	---Version:

	---Purpose: This class allows the definition of a Line Style.
	--	    The Style can be Predefined or defined by the user

	---Keywords: LineStyle 

	---Warning:
	---References:

uses
	TypeOfLine from Aspect,
	Array1OfLength from TColQuantity,
	HArray1OfLength from TColQuantity

raises
	LineStyleDefinitionError from Aspect

is
	Create
		returns LineStyle from Aspect
	---Level: Public
	---Purpose: Creates a line style with the default value of
	--	    LineStyle type : SOLID
	--
	raises LineStyleDefinitionError from Aspect;
	-- if the maximum number of line style is exceeded

	Create ( Type	: TypeOfLine from Aspect )
		returns LineStyle from Aspect ;
	---Level: Public
	---Purpose: Creates the line style <Type>.

	Create ( Style : Array1OfLength from TColQuantity ) 
		returns LineStyle from Aspect
	---Level: Public
	---Purpose: Creates a line style from METER Float style descriptor .
	--	    Style Descriptor is :
	--	    Each Odd float described the Drawn part of the style .
	--	    Each Even float described the Hidden part of the style .
	--	    (e.g) [0.010,0.002,0.005,0.004] 
	--		  Draw 10 MM ,Move 2 MM,Draw 5 MM ..
	raises LineStyleDefinitionError from Aspect;
	-- if the METER float values are <= 0. 

	---------------------------------------------------
	-- Category: Methods to modify the class definition
	---------------------------------------------------

	Assign ( me	: in out ;
		 Other	: LineStyle from Aspect )
		returns LineStyle from Aspect is static;
	---Level: Public
	---Purpose: Updates the line style <me> from the definition of the
	--	    line style <Other>.
	---Category: Methods to modify the class definition
	---C++: alias operator =
	---C++: return &

	SetValues ( me		: in out ;
		    Type	: TypeOfLine from Aspect )  is static;
	---Level: Public
	---Purpose: Updates the line style <me> from the definition of the
	--	    line style <Type>.
	---Category: Methods to modify the class definition

	SetValues ( me		: in out ;
		    Style : Array1OfLength from TColQuantity )
	---Level: Public
	---Purpose: Updates a line style with the new Float descriptor
	raises LineStyleDefinitionError from Aspect is static;
	-- if the METER float values are <= 0. 
	---Category: Methods to modify the class definition

	----------------------------
	-- Category: Inquire methods
	----------------------------

	Style ( me )
		returns TypeOfLine from Aspect is static;
	---Level: Public
	---Purpose: Returns the type of the line style <me> 
	---Category: Inquire methods

	Length ( me )
		returns Integer from Standard  is static;
	---Level: Public
	---Purpose: Returns the components length of the line style
	---Category: Inquire methods

	Values ( me ) 
		returns Array1OfLength from TColQuantity  is static;
	---Level: Public
	---Purpose: Returns the components of a line style 
	---Category: Inquire methods
	---C++: return const &

    	IsEqual(me; Other : LineStyle from Aspect) returns Boolean;
	    ---C++: alias operator==

    	IsNotEqual(me; Other : LineStyle from Aspect) returns Boolean;
	    ---C++: alias operator!=

	----------------------------
	-- Category: Private methods
	----------------------------

	PredefinedStyle ( me : in out  ;
		          Type : TypeOfLine from Aspect )  
	---Level: Internal
	---Purpose: Set MyLineDescriptor with the predefined style values
	--	    according of type
	---Category: Private methods
	returns HArray1OfLength from TColQuantity is static private;

--

fields

--
-- Class	:	Aspect_LineStyle
--
-- Purpose	:	Declaration of variables specific to line styles
--

	MyLineType		: TypeOfLine from Aspect;
	MyLineDescriptor	: HArray1OfLength from TColQuantity;

end LineStyle;
