-- Created on: 1996-01-09
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Generator from LocOpe

	---Purpose: 

uses GeneratedShape      from LocOpe,

     Shape               from TopoDS,
     Face                from TopoDS,
     Edge                from TopoDS,
     
     ListOfShape         from TopTools,
     DataMapOfShapeListOfShape from TopTools
--     DataMapOfShapeShape from TopTools
     
     
     
raises NotDone      from StdFail,
       NullObject   from Standard,
       NoSuchObject from Standard

is

    Create
	---Purpose: Empty constructor.
    	returns Generator from LocOpe;
    	---C++: inline


    Create(S: Shape from TopoDS)
	---Purpose: Creates the algorithm on the shape <S>.
	---C++: inline
    	returns Generator from LocOpe;


    Init(me: in out; S: Shape from TopoDS)
	---Purpose: Initializes the algorithm on the shape <S>.
	---C++: inline
    	is static;


    Perform(me: in out; G: GeneratedShape from LocOpe)
			
	raises NullObject from Standard		
    	is static;


    IsDone(me)
    
	---C++: inline
    	returns Boolean from Standard
	is static;



    ResultingShape(me)
	---Purpose: Returns the new shape
    	returns Shape from TopoDS
	---C++: return const&
	---C++: inline
	raises NotDone from StdFail
	is static;
	

    Shape(me)
	---Purpose: Returns the initial shape
    	returns Shape from TopoDS
	---C++: return const&
	---C++: inline
	is static;


    DescendantFace(me: in out; F: Face from TopoDS)
    	---Purpose: Returns  the  descendant  face  of <F>.    <F> may
    	--          belong to the original shape or to the "generated"
    	--          shape.  The returned    face may be   a null shape
    	--          (when <F> disappears). 
	---C++: return const&
    	returns ListOfShape from TopTools


	raises NotDone from StdFail,
	--- The exception is raised when IsDone returns <Standard_False>.
	       NoSuchObject from Standard
	--- The exception is  raised when <F> does  not  belong to the
	--  original  shape or to the "generated" one.
	is static;


fields

    myShape     : Shape                 from TopoDS;
    myGen       : GeneratedShape        from LocOpe;
    myDone      : Boolean               from Standard;
    myRes       : Shape                 from TopoDS;
    myModShapes : DataMapOfShapeListOfShape from TopTools;

end Generator;













