-- Created on: 1995-10-20
-- Created by: Yves FRICAUD
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Interval from BRepOffset 

	---Purpose: 

uses
    Type from BRepOffset
    
is

    Create;
    
    Create (U1,U2 : Real from Standard;
    	    Type  : Type from BRepOffset)
    returns Interval from BRepOffset;
    
    First (me : in out; U : Real from Standard)
    	---C++: inline
    is static;
    
    Last  (me : in out; U : Real from Standard)
        ---C++: inline
    is static;    
    
    Type  (me : in out; T : Type from BRepOffset)
       ---C++: inline
    is static;
    
    First (me) returns Real from Standard
       ---C++: inline
    is static;    
    
    Last  (me) returns Real from Standard
       ---C++: inline
    is static;
    
    Type  (me) returns Type from BRepOffset
       ---C++: inline
    is static;    
    

fields

    f,l  : Real from Standard;
    type : Type from BRepOffset;
    
end Interval;
