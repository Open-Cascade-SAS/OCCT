-- Created on: 1996-02-15
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class FindEdges from LocOpe

	---Purpose: 

uses Shape                      from TopoDS,
     Edge                      from TopoDS,
     ListOfShape               from TopTools,
     ListIteratorOfListOfShape from TopTools
     

raises ConstructionError from Standard,
       NoSuchObject      from Standard,
       NoMoreObject      from Standard

is

    Create
    	returns FindEdges from LocOpe;
	---C++: inline



    Create(FFrom,FTo: Shape from TopoDS)
    
	---C++: inline
    	returns FindEdges from LocOpe
	raises ConstructionError from Standard;
	
	
    Set(me: in out; FFrom, FTo: Shape from TopoDS)
    
	raises ConstructionError from Standard
    	is static;


    InitIterator(me: in out)
    
	---C++: inline
    	is static;


    More(me)
    
    	returns Boolean from Standard
	---C++: inline
	is static;


    EdgeFrom(me)
    
    	returns Edge from TopoDS
	---C++: return const&
	---C++: inline
	raises NoSuchObject from Standard
	is static;


    EdgeTo(me)
    
    	returns Edge from TopoDS
	---C++: return const&
	---C++: inline
	raises NoSuchObject from Standard
	is static;


    Next(me: in out)
    
	---C++: inline
    	raises NoMoreObject from Standard
	is static;


fields

    myFFrom  : Shape                     from TopoDS;
    myFTo    : Shape                     from TopoDS;
    myLFrom  : ListOfShape               from TopTools;
    myLTo    : ListOfShape               from TopTools;
    myItFrom : ListIteratorOfListOfShape from TopTools;
    myItTo   : ListIteratorOfListOfShape from TopTools;

end FindEdges;
