-- Created on: 1995-01-06
-- Created by: Christophe MARION
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class FaceIsoLiner from HLRTopoBRep

uses
    Integer from Standard,
    Real    from Standard,
    Pnt     from gp,
    Line    from Geom2d,
    Face    from TopoDS,
    Edge    from TopoDS,
    Vertex  from TopoDS,
    Data    from HLRTopoBRep

is
    Perform( myclass;
             FI     :        Integer from Standard;
             F      :        Face    from TopoDS;
    	     DS     : in out Data    from HLRTopoBRep;
	     nbIsos :        Integer from Standard);

    MakeVertex( myclass;
                E   :        Edge from TopoDS;
                P   :        Pnt  from gp;
                Par :        Real from Standard;
                Tol :        Real from Standard;
    	        DS  : in out Data from HLRTopoBRep)
    returns Vertex from TopoDS; 

    MakeIsoLine( myclass;
             F   :        Face   from TopoDS;
	     Iso :        Line   from Geom2d;	
             V1  : in out Vertex from TopoDS;
             V2  : in out Vertex from TopoDS;
             U1  :        Real   from Standard;
             U2  :        Real   from Standard;
             Tol :        Real   from Standard;
             DS  : in out Data   from HLRTopoBRep);

end FaceIsoLiner;
