-- File:        Vertex.cdl
-- Created:     Mon Dec  4 12:02:33 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWVertex from RWStepShape

	---Purpose : Read & Write Module for Vertex

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     Vertex from StepShape

is

	Create returns RWVertex;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable Vertex from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : Vertex from StepShape);

end RWVertex;
