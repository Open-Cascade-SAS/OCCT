-- Created on: 1997-05-27
-- Created by: Sergey SOKOLOV
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DoubleJacobiPolynomial from PLib 

	---Purpose: 

uses Array1OfReal,HArray1OfReal from TColStd, 
     JacobiPolynomial from PLib

is  
    Create returns DoubleJacobiPolynomial; 
    
    Create ( JacPolU, JacPolV : JacobiPolynomial from  PLib)  
      returns DoubleJacobiPolynomial;

    MaxErrorU ( me; Dimension, DegreeU, DegreeV, dJacCoeff : Integer; 
    	    	JacCoeff : Array1OfReal from TColStd ) returns Real;
     
    MaxErrorV ( me; Dimension, DegreeU, DegreeV, dJacCoeff : Integer; 
    	    	JacCoeff : Array1OfReal from TColStd ) returns Real;
    
    MaxError ( me; Dimension, MinDegreeU, MaxDegreeU,  
    	       MinDegreeV, MaxDegreeV, dJacCoeff : Integer; 
    	       JacCoeff : Array1OfReal from TColStd; Error : Real ) returns Real;

    ReduceDegree ( me; Dimension, MinDegreeU, MaxDegreeU,  
    	       	   MinDegreeV, MaxDegreeV, dJacCoeff : Integer; 
    	       	   JacCoeff : Array1OfReal from TColStd; EpmsCut : Real; 
    	    	   MaxError : in out Real;  NewDegreeU, NewDegreeV : in out Integer);

    AverageError ( me; Dimension, DegreeU, DegreeV, dJacCoeff : Integer; 
    	    	   JacCoeff : Array1OfReal from TColStd ) returns Real;

    WDoubleJacobiToCoefficients ( me; Dimension, DegreeU, DegreeV : Integer; 
    	    	                  JacCoeff : Array1OfReal from TColStd; 
    	    	    	    	  Coefficients : out Array1OfReal from TColStd ); 
				   
    U (me) 
--- Purpose: returns myJacPolU;
    ---C++: inline
    returns JacobiPolynomial from PLib;

    V (me) 
--- Purpose: returns myJacPolV;
    ---C++: inline
    returns JacobiPolynomial from PLib;

    TabMaxU (me) 
--- Purpose: returns myTabMaxU;
    ---C++: inline
    returns HArray1OfReal from TColStd;

    TabMaxV (me) 
--- Purpose: returns myTabMaxV;
    ---C++: inline
    returns HArray1OfReal from TColStd;

fields
 
    myJacPolU     : JacobiPolynomial from PLib;
    myJacPolV     : JacobiPolynomial from PLib; 
    myTabMaxU     : HArray1OfReal from TColStd;
    myTabMaxV     : HArray1OfReal from TColStd;
    
end DoubleJacobiPolynomial;
