-- Created on: 1998-09-03
-- Created by: Julia GERASIMOVA
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

private class FaceAndOrder from BRepFill

	---Purpose: A structure containing Face and Order of constraint

uses
    Face from TopoDS, 
    Shape from GeomAbs
is
    Create returns FaceAndOrder from BRepFill;
    
    Create( aFace   : Face from TopoDS; 
    	    anOrder : Shape from GeomAbs )
    returns FaceAndOrder from BRepFill;

    --Face(me : in out) returns Face from TopoDS;
    -- ---C++: return &
    --Order(me : in out) returns Integer from Standard;
    -- ---C++: return &

fields

    myFace  : Face from TopoDS;
    myOrder : Shape from GeomAbs;

friends
    class Filling from BRepFill

end FaceAndOrder;
