-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class RevolvedAreaSolid from StepShape 

inherits SweptAreaSolid from StepShape 

uses

	Axis1Placement from StepGeom, 
	Real from Standard, 
	HAsciiString from TCollection, 
	CurveBoundedSurface from StepGeom
is

	Create returns mutable RevolvedAreaSolid;
	---Purpose: Returns a RevolvedAreaSolid


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aSweptArea : mutable CurveBoundedSurface from StepGeom) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aSweptArea : mutable CurveBoundedSurface from StepGeom;
	      aAxis : mutable Axis1Placement from StepGeom;
	      aAngle : Real from Standard) is virtual;

	-- Specific Methods for Field Data Access --

	SetAxis(me : mutable; aAxis : mutable Axis1Placement);
	Axis (me) returns mutable Axis1Placement;
	SetAngle(me : mutable; aAngle : Real);
	Angle (me) returns Real;

fields

	axis : Axis1Placement from StepGeom;
	angle : Real from Standard;

end RevolvedAreaSolid;
