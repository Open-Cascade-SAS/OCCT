-- Created on: 1996-01-23
-- Created by: Laurent PAINNOT
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class   GenExtCS from Extrema 

    	---Purpose: It calculates all the extremum distances
    	--          between acurve and a surface.
    	--          These distances can be minimum or maximum.

uses  POnSurf       from Extrema,
      POnCurv       from Extrema,
      Pnt           from gp,
      HArray1OfPnt  from TColgp,
      HArray2OfPnt  from TColgp,
      FuncExtCS     from Extrema,
      Surface       from Adaptor3d,
      SurfacePtr    from Adaptor3d,
      Curve         from Adaptor3d,
      CurvePtr      from Adaptor3d

raises  NotDone      from StdFail,
    	OutOfRange   from Standard,
	TypeMismatch from Standard
	

is

    Create returns GenExtCS;
    
    Create (C: Curve from Adaptor3d; S: Surface from Adaptor3d; 
    	    NbT: Integer; NbU,NbV: Integer; Tol1,Tol2: Real)
    	returns GenExtCS;
      	---Purpose: It calculates all the distances.
        --          The function F(u,v)=distance(S1(u1,v1),S2(u2,v2)) has an 
        --          extremum when gradient(F)=0. The algorithm searchs
        --          all the zeros inside the definition ranges of the 
        --          surfaces.
      	--          NbU and NbV are used to locate the close points on the
      	--          surface and NbT on the curve to find the zeros. 

    Create (C: Curve from Adaptor3d; S: Surface from Adaptor3d; 
    	    NbT,NbU,NbV: Integer; 
    	    tmin, tsup: Real; 
    	    Umin, Usup, Vmin, Vsup: Real; 
    	    Tol1,Tol2: Real)
    	returns GenExtCS;
      	---Purpose: It calculates all the distances.
        --          The function F(u,v)=distance(P,S(u,v)) has an 
        --          extremum when gradient(F)=0. The algorithm searchs
        --          all the zeros inside the definition ranges of the 
        --          surface.
      	--          NbT,NbU and NbV are used to locate the close points
      	--          to find the zeros. 
    
    Initialize(me: in out; S: Surface from Adaptor3d; 
    	       NbU, NbV: Integer; Tol2: Real)
    	---Pupose: sets the fields of the algorithm.
    is static;


    Initialize(me: in out; S: Surface from Adaptor3d; NbU, NbV: Integer; 
    	       Umin, Usup, Vmin, Vsup: Real; Tol2: Real)
    	---Pupose: sets the fields of the algorithm.
    is static;
    

    Perform(me: in out; C: Curve from Adaptor3d; 
    	    NbT: Integer; Tol1: Real)
        ---Purpose: the algorithm is done with S
        --          An exception is raised if the fields have not
        --          been initialized.  
    raises TypeMismatch from Standard
    is static;

    Perform(me: in out; C: Curve from Adaptor3d; NbT: Integer;
            tmin, tsup: Real; Tol1: Real)
        ---Purpose: the algorithm is done with C
        --          An exception is raised if the fields have not
        --          been initialized.  
    raises TypeMismatch from Standard
    is static;


    IsDone (me) returns Boolean
    	---Purpose: Returns True if the distances are found.
    	is static;
    
    NbExt (me) returns Integer
    	---Purpose: Returns the number of extremum distances.
    	raises  NotDone from StdFail
	    	-- if IsDone(me)=False.
    	is static;

    SquareDistance(me; N: Integer) returns Real
    	---Purpose: Returns the value of the Nth resulting square distance.
    	raises  NotDone from StdFail,
    	    	-- if IsDone(me)=False.
    	        OutOfRange
		-- if N < 1 or N > NbPoints(me).
    	is static;

    PointOnCurve (me; N: Integer) returns POnCurv
    	---Purpose: Returns the point of the Nth resulting distance.
    	---C++: return const&
    	raises  NotDone from StdFail,
    	    	-- if IsDone(me)=False.
    	        OutOfRange
		-- if N < 1 or N > NbPoints(me).
    	is static;

    PointOnSurface (me; N: Integer) returns POnSurf
    	---Purpose: Returns the point of the Nth resulting distance.
    	---C++: return const&
    	raises  NotDone from StdFail,
    	    	-- if IsDone(me)=False.
    	        OutOfRange
		-- if N < 1 or N > NbPoints(me).
    	is static;

    BidonCurve(me) returns CurvePtr from Adaptor3d
    is static private;

    BidonSurface(me) returns SurfacePtr from Adaptor3d
    is static private;

fields
    myDone     : Boolean;
    myInit     : Boolean;
    mytmin     : Real;
    mytsup     : Real;
    myumin     : Real;
    myusup     : Real;
    myvmin     : Real;
    myvsup     : Real;
    mytsample  : Integer;
    myusample  : Integer;
    myvsample  : Integer;
    mytol1     : Real;
    mytol2     : Real;
    myF        : FuncExtCS from Extrema;
    myS        : SurfacePtr from Adaptor3d;
    mySurfPnts : HArray2OfPnt from TColgp;

end GenExtCS;
