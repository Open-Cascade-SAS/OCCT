-- Created on: 1993-05-07
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class VPointInterIterator from TopOpeBRep

    -- ==========================
    -- Restriction Point iterator
    -- ==========================

uses

    LineInter from TopOpeBRep,
    PLineInter from TopOpeBRep,
    VPointInter from TopOpeBRep

is

    Create returns VPointInterIterator from TopOpeBRep;
    Create(LI : LineInter from TopOpeBRep)  
    returns VPointInterIterator from TopOpeBRep;

    Init(me:in out; LI : LineInter from TopOpeBRep;
    	    	    checkkeep : Boolean from Standard = Standard_False) is static;
    Init(me:in out) is static;
    More(me) returns Boolean is static;
    Next(me:in out) is static;
 
    CurrentVP(me:in out) returns VPointInter from TopOpeBRep is static;
    ---C++: return const &

    CurrentVPIndex(me) returns Integer is static;

    ChangeCurrentVP(me:in out) returns VPointInter from TopOpeBRep is static;
    ---C++: return &

    PLineInterDummy(me) returns PLineInter from TopOpeBRep;
    
fields

    myLineInter : PLineInter from TopOpeBRep;
    myVPointIndex : Integer;    
    myVPointNb : Integer;
    mycheckkeep : Boolean from Standard;

end VPointInterIterator from TopOpeBRep;
