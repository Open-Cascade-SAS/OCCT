-- Created on: 1993-01-09
-- Created by: CKY / Contract Toubro-Larsen ( TCD )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class IntercharacterSpacing from IGESGraph  inherits IGESEntity

        ---Purpose: defines IGESIntercharacterSpacing, Type <406> Form <18>
        --          in package IGESGraph
        --
        --          Specifies the gap between letters when fixed-pitch
        --          spacing is used

uses  Integer, Real  -- no one specific type


is

        Create returns mutable IntercharacterSpacing;

        -- Specific Methods pertaining to the class

        Init (me       : mutable;
              nbProps  : Integer;
              anISpace : Real);
        ---Purpose : This method is used to set the fields of the class
        --           IntercharacterSpacing
        --       - nbProps  : Number of property values (NP = 1)
        --       - anISpace : Intercharacter spacing percentage

        NbPropertyValues (me) returns Integer;
        ---Purpose : returns the number of property values in <me>

        ISpace (me) returns Real;
        ---Purpose : returns the Intercharacter Space of <me> in percentage
        -- of the text height (Range = 0..100)

fields

--
-- Class    : IGESGraph_IntercharacterSpacing
--
-- Purpose  : Declaration of the variables specific to a
--            Intercharacter Spacing property.
--
-- Reminder : An Intercharacter spacing property is defined by :
--                  - Number of property values (NP=1)
--                  - ISpace
--

        theNbPropertyValues : Integer;

        theISpace           : Real;

end IntercharacterSpacing;
