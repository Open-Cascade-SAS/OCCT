-- File:	StepBasic_ExternallyDefinedItem.cdl
-- Created:	Wed May 10 15:09:07 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class ExternallyDefinedItem from StepBasic
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity ExternallyDefinedItem

uses
    SourceItem from StepBasic,
    ExternalSource from StepBasic

is
    Create returns ExternallyDefinedItem from StepBasic;
	---Purpose: Empty constructor

    Init (me: mutable; aItemId: SourceItem from StepBasic;
                       aSource: ExternalSource from StepBasic);
	---Purpose: Initialize all fields (own and inherited)

    ItemId (me) returns SourceItem from StepBasic;
	---Purpose: Returns field ItemId
    SetItemId (me: mutable; ItemId: SourceItem from StepBasic);
	---Purpose: Set field ItemId

    Source (me) returns ExternalSource from StepBasic;
	---Purpose: Returns field Source
    SetSource (me: mutable; Source: ExternalSource from StepBasic);
	---Purpose: Set field Source

fields
    theItemId: SourceItem from StepBasic;
    theSource: ExternalSource from StepBasic;

end ExternallyDefinedItem;
