-- Created on: 1994-02-21
-- Created by: Laurent PAINNOT
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class MCurvesToBSpCurve from Approx



uses MultiBSpCurve        from AppParCurves,
     MultiCurve           from AppParCurves,
     SequenceOfMultiCurve from AppParCurves

is


    Create returns MCurvesToBSpCurve;
    
    Reset(me: in out) 
    	--- Clear the internal Sequence Of MultiCurve
    is static;
    
    Append(me: in out; MC: MultiCurve from AppParCurves)
    is static;


    Perform(me: in out)
    is static;
    
    Perform(me: in out; TheSeq: SequenceOfMultiCurve from AppParCurves)
    is static;
    
    
    Value(me)
    	---Purpose: return the composite MultiCurves as a MultiBSpCurve.
    	---C++: return const&

    returns MultiBSpCurve
    is static;


    ChangeValue(me: in out)
    	---Purpose: return the composite MultiCurves as a MultiBSpCurve.
    	---C++: return const&

    returns MultiBSpCurve
    is static;


fields


mySpline: MultiBSpCurve           from AppParCurves;
myDone  : Boolean                 from Standard;
myCurves: SequenceOfMultiCurve    from AppParCurves; 

end MCurvesToBSpCurve;
