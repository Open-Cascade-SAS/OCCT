-- Created on: 1991-10-04
-- Created by: Remi GILET
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class BCirc from GccInt 

inherits Bisec from GccInt 

     	---Purpose: Describes a circle as a bisecting curve between two 2D
    	-- geometric objects (such as circles or points).

uses Circ2d from gp,
     IType  from GccInt

is

Create(Circ : Circ2d) returns mutable BCirc;
    	---Purpose: Constructs a bisecting curve whose geometry is the 2D circle Circ.
    
Circle(me) returns Circ2d from gp
    is redefined;
    	---Purpose: Returns a 2D circle which is the geometry of this bisecting curve.    

    ArcType(me) returns IType from GccInt
    is static;
    	---Purpose: Returns GccInt_Cir, which is the type of any GccInt_BCirc bisecting curve.

fields

    cir : Circ2d from gp;
    ---Purpose: The bisecting line.

end BCirc;    


