-- Created on: 1995-06-08
-- Created by: Robert COUBLANC
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class BasicTool from SelectBasics 

	---Purpose: give Tools for sorting Selection results
    --          (example : sensitive entities matching)

uses
    Pnt2d from gp,
    Array1OfPnt2d from TColgp
is

    MatchSegments(myclass;
    	    	  P1,P2 : Pnt2d from gp;
    	    	  P3,P4 : Pnt2d from gp)
    returns Boolean;
    ---Purpose: returns True if The Segment {P1P2} is
    --          intersected by the segment {P3P4}

    MatchSegment(myclass;
		 pBegin,pEnd : Pnt2d from gp;
		 X,Y,aTol    : Real;
	         DMin        : in out Real) returns Boolean;
    ---Level: Internal
    ---Purpose: return True if Segment(pBegin, pEnd) is Selected 
 
    AutoInter(myclass; aPolyg2d: Array1OfPnt2d from TColgp)
    returns Boolean;
      
    MatchPolyg2d (myclass;
    	    	  tabpoint: Array1OfPnt2d from TColgp;
    	    	  X,Y,aTol: Real;
	          DMin    : in out Real;
    	    	  Rank    : in out Integer) returns Boolean;
    ---Level: Internal 
    ---Purpose: package method used to find if a point 
    --          is close enough to a polygon of 2D points
    --          to be Used by Primitives like curves or faces...
    --          Rank gives the index of the touched
    --          segment

    


end BasicTool;
