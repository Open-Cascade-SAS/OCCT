-- Created on: 1993-07-12
-- Created by: Martine LANGLOIS
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MakePolyline from GeomToStep inherits Root from GeomToStep

    ---Purpose: This class implements the mapping between an Array1 of points
    --          from gp and a Polyline from StepGeom.
  
uses Array1OfPnt from TColgp,
     Array1OfPnt2d from TColgp,
     Polyline from StepGeom
     
raises NotDone from StdFail
     
is 

Create ( P : Array1OfPnt from TColgp ) returns MakePolyline;

Create ( P : Array1OfPnt2d from TColgp ) returns MakePolyline;

Value (me) returns Polyline from StepGeom
    raises NotDone
    is static;
    ---C++: return const&

fields

    thePolyline : Polyline from StepGeom;
    	-- The solution from StepGeom
    	
end MakePolyline;


