-- Created on: 2000-04-18
-- Created by: Andrey BETENEV
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0

class DimensionalCharacteristic from StepShape
inherits SelectType from StepData

    ---Purpose: Representation of STEP SELECT type DimensionalCharacteristic

uses
    DimensionalLocation from StepShape,
    DimensionalSize from StepShape

is
    Create returns DimensionalCharacteristic from StepShape;
	---Purpose: Empty constructor

    CaseNum (me; ent: Transient) returns Integer;
	---Purpose: Recognizes a kind of DimensionalCharacteristic select type
	--          1 -> DimensionalLocation from StepShape
	--          2 -> DimensionalSize from StepShape
	--          0 else

    DimensionalLocation (me) returns DimensionalLocation from StepShape;
	---Purpose: Returns Value as DimensionalLocation (or Null if another type)

    DimensionalSize (me) returns DimensionalSize from StepShape;
	---Purpose: Returns Value as DimensionalSize (or Null if another type)

end DimensionalCharacteristic;
