-- File:	StepShape_SeamEdge.cdl
-- Created:	Fri Jan  4 17:42:44 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class SeamEdge from StepShape
inherits OrientedEdge from StepShape

    ---Purpose: Representation of STEP entity SeamEdge

uses
    HAsciiString from TCollection,
    Vertex from StepShape,
    Edge from StepShape,
    Pcurve from StepGeom

is
    Create returns SeamEdge from StepShape;
	---Purpose: Empty constructor

    
		       
    Init (me: mutable; aRepresentationItem_Name: HAsciiString from TCollection;	       
                       aOrientedEdge_EdgeElement: Edge from StepShape;
                       aOrientedEdge_Orientation: Boolean;
                       aPcurveReference: Pcurve from StepGeom);
	---Purpose: Initialize all fields (own and inherited)

    PcurveReference (me) returns Pcurve from StepGeom;
	---Purpose: Returns field PcurveReference
    SetPcurveReference (me: mutable; PcurveReference: Pcurve from StepGeom);
	---Purpose: Set field PcurveReference

fields
    thePcurveReference: Pcurve from StepGeom;

end SeamEdge;
