-- File:	GeomLib_CheckBSplineCurve.cdl
-- Created:	Wed May 28 16:31:08 1997
-- Author:	Xavier BENVENISTE
--		<xab@zozox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1997



class Check2dBSplineCurve from GeomLib

	---Purpose: this class is used to  construct the BSpline curve
	--          from an Approximation ( ApproxAFunction from AdvApprox).
    	

uses
    Pnt2d           from gp,
    BSplineCurve    from Geom2d

raises

    NotDone    from StdFail,
    OutOfRange from Standard
    
is

    Create( Curve : BSplineCurve from Geom2d ;
    	    Tolerance        : Real from Standard ;
            AngularTolerance : Real from Standard) 
    returns Check2dBSplineCurve from GeomLib;
    
    IsDone(me) returns Boolean from Standard
	---C++: inline
    is static;
    
    NeedTangentFix(me; FirstFlag : in out Boolean from Standard ;
    	         SecondFlag : in out Boolean from Standard) ;
    FixTangent  (me : in out ; FirstFlag : Boolean from Standard ;
              		       LastFlag  : Boolean from Standard)  ;	 
	
    FixedTangent  (me : in out ; FirstFlag : Boolean from Standard ;
              		       LastFlag  : Boolean from Standard) 
    ---Purpose:  modifies the curve
    -- by fixing the first or the last tangencies 
    -- 
    returns BSplineCurve from Geom2d
    raises
    	OutOfRange from Standard,
    	---Purpose: if Index3D not in the Range [1,Nb3dSpaces]
	NotDone    from StdFail
	---Purpose: if the Approx is not Done
    is static;
 

fields

    myCurve            : BSplineCurve from Geom2d ;
    myDone             : Boolean from Standard ;
    myFixFirstTangent  : Boolean from Standard ;
    myFixLastTangent   : Boolean from Standard ;
    myAngularTolerance : Real from Standard ;
    myTolerance        : Real from Standard ;
    myFirstPole        : Pnt2d from gp ;
    	-- the second pole that controls first tangency
    myLastPole         : Pnt2d from gp ;
    	-- the before last pole that controls last tangency

end Check2dBSplineCurve;
