-- Created on: 1992-10-14
-- Created by: Christophe MARION
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package HLRBRep 
    ---Purpose: Hidden Lines Removal
    --          algorithms on the BRep DataStructure.
    --          
    --          The class PolyAlgo  is used to remove Hidden lines
    --          on Shapes with Triangulations.

uses
    Standard,
    StdFail,
    MMgt,
    gp,
    Geom,
    Geom2d,
    TCollection,
    TColgp,
    TColStd,
    GeomAbs,
    LProp,
    IntRes2d,
    IntCurve,
    IntCurveSurface,
    TopAbs,
    TopoDS,
    TopExp,
    TopTools,
    HLRAlgo,
    Adaptor3d,
    BRep,
    BRepAdaptor,
    BRepTopAdaptor,
    HLRTopoBRep

is
    class CurveTool;
    class BCurveTool;
    class Curve;
    class SurfaceTool;
    class BSurfaceTool;
    class Surface;

    class CLPropsATool;
    class CLProps       instantiates CLProps          from LProp (
    	Address      from Standard, -- as Curve from HLRBRep
	Vec2d        from gp,
	Pnt2d        from gp,
	Dir2d        from gp,
	CLPropsATool from HLRBRep);

    class SLPropsATool;
    class SLProps       instantiates SLProps          from LProp (
    	Address      from Standard, -- as Surface from HLRBRep
	SLPropsATool from HLRBRep);

    class CInter        instantiates IntCurveCurveGen from IntCurve ( 
    	Address   from Standard,
    	CurveTool from HLRBRep);

    class LineTool;

    class InterCSurf    instantiates Inter            from IntCurveSurface (
    	Lin         from gp,
	LineTool    from HLRBRep,
    	Address     from Standard,
        SurfaceTool from HLRBRep);

    class EdgeFaceTool;

    class Intersector;
    
    class EdgeData;
	
    class FaceData;
    
    class FaceIterator;
	
    imported Array1OfEData;

    imported Array1OfFData;

    class Data;

    class ShapeToHLR;

    class HLRToShape;

    class ShapeBounds;

    imported SeqOfShapeBounds;

    class EdgeInterferenceTool;

    class VertexList;

    class EdgeIList;
    
    class AreaLimit;
    
    class EdgeBuilder;

    class Hider;
    
    class InternalAlgo;
    
    class Algo;

    class PolyAlgo;

    class BiPoint;
    class BiPnt2D;
    
    imported ListOfBPoint;
    
    imported ListIteratorOfListOfBPoint;

    imported ListOfBPnt2D;

    imported ListIteratorOfListOfBPnt2D;

    class PolyHLRToShape;

    MakeEdge(ec    : Curve from HLRBRep;
             U1,U2 : Real  from Standard)
    returns Edge from TopoDS;
    
    MakeEdge3d(ec    : Curve from HLRBRep;
               U1,U2 : Real  from Standard)
    returns Edge from TopoDS;
    
    PolyHLRAngleAndDeflection(InAngl           :     Real from Standard;
                              OutAngl, OutDefl : out Real from Standard);
    
end HLRBRep;
