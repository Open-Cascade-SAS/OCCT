-- Created on: 2002-08-02
-- Created by: Alexander KARTOMIN  (akm)
-- Copyright (c) 2002-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- NB:          This originates from BRepLProp being abstracted of BRep.

class CurveTool from LProp3d

uses Vec   from gp,
     Pnt   from gp,
     Dir   from gp,
     HCurve from Adaptor3d

is

    Value(myclass; C : HCurve from Adaptor3d; U : Real; P : out Pnt);
    ---Purpose: Computes the point <P> of parameter <U> on the HCurve <C>.
        
    D1   (myclass; C : HCurve from Adaptor3d; 
          U : Real; P : out Pnt; V1 : out Vec);
    ---Purpose: Computes the point <P> and first derivative <V1> of 
    --          parameter <U> on the HCurve <C>.

    D2   (myclass; C : HCurve from Adaptor3d; 
          U : Real; P : out Pnt; V1, V2 : out Vec);
    ---Purpose: Computes the point <P>, the first derivative <V1> and second
    --          derivative <V2> of parameter <U> on the HCurve <C>.
    
    D3   (myclass; C : HCurve from Adaptor3d; 
          U : Real; P : out Pnt; V1, V2, V3 : out Vec);
    ---Purpose: Computes the point <P>, the first derivative <V1>, the 
    --          second derivative <V2> and third derivative <V3> of 
    --          parameter <U> on the HCurve <C>.

     Continuity(myclass; C : HCurve from Adaptor3d) returns Integer;
     ---Purpose: returns the order of continuity of the HCurve <C>.
     --          returns 1 : first derivative only is computable
     --          returns 2 : first and second derivative only are computable.
     --          returns 3 : first, second and third are computable.

     FirstParameter(myclass; C : HCurve from Adaptor3d) returns Real;
     ---Purpose: returns the first parameter bound of the HCurve.
     --          
     
     LastParameter(myclass; C : HCurve from Adaptor3d) returns Real;
     ---Purpose: returns the last parameter bound of the HCurve.
     --          FirstParameter must be less than LastParamenter.

end CurveTool;


