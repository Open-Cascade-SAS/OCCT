-- Created on: 1998-06-03
-- Created by: data exchange team
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Geom from ShapeAnalysis 

    ---Purpose: Analyzing tool aimed to work on primitive geometrical objects

uses
    HArray2OfReal from TColStd,
    Trsf from gp,
    Pln from gp,
    Array1OfPnt from TColgp

raises
   OutOfRange from Standard
    
is
    NearestPlane (myclass; Pnts: Array1OfPnt from TColgp;
    	    	     	   aPln: out Pln from gp;
    	    	    	   Dmax: out Real)
    returns Boolean;
    	---Purpose : Builds a plane out of a set of points in array
	--           Returns in <dmax> the maximal distance between the produced
	--           plane and given points

    PositionTrsf (myclass; coefs: HArray2OfReal from TColStd;
                    	   trsf: out Trsf from gp;
    	    	           unit, prec : Real)
    returns Boolean
    	---Purpose: Builds transfromation object out of matrix.
	--          Matrix must be 3 x 4.
    	--          Unit is used as multiplier.
    raises OutOfRange from Standard;
    	--          If numer of rows is greater than 3 or number of columns is
    	--          greater than 4

end Geom;
