-- File:	BRepBuilderAPI_MakeSolid.cdl
-- Created:	Wed Jul 21 16:06:45 1993
-- Author:	Remi LEQUETTE
--		<rle@nonox>
---Copyright:	 Matra Datavision 1993


class MakeSolid from BRepBuilderAPI  inherits MakeShape from BRepBuilderAPI

	---Purpose: Describes functions to build a solid from shells.
    	-- A solid is made of one shell, or a series of shells, which
    	-- do not intersect each other. One of these shells
    	-- constitutes the outside skin of the solid. It may be closed
    	-- (a finite solid) or open (an infinite solid). Other shells
    	-- form hollows (cavities) in these previous ones. Each
    	-- must bound a closed volume.
    	-- A MakeSolid object provides a framework for:
    	-- -   defining and implementing the construction of a solid, and
    	-- -   consulting the result.

uses
    Solid     from TopoDS,
    CompSolid from TopoDS,
    Shell     from TopoDS,
    Shape     from TopoDS,
    MakeSolid from BRepLib

raises
    NotDone from StdFail
    
is

    Create
	---Purpose: Initializes the construction of a solid. An empty solid is
    	-- considered to cover the whole space. The Add function
    	-- is used to define shells to bound it.
    returns MakeSolid from BRepBuilderAPI;

    ----------------------------------------------
    -- From Compsolid
    ----------------------------------------------

    Create(S : CompSolid from TopoDS)
	---Purpose: Make a solid from a CompSolid.
	---Level: Public
    returns MakeSolid from BRepBuilderAPI;

    --  this  algorithm  removes  all  inner  faces  amd  make  solid  from  compsolid

    ----------------------------------------------
    -- From shells
    ----------------------------------------------

    Create(S : Shell from TopoDS)
	---Purpose: Make a solid from a shell.
	---Level: Public
    returns MakeSolid from BRepBuilderAPI;

    
    Create(S1,S2 : Shell from TopoDS)
	---Purpose: Make a solid from two shells.
	---Level: Public
    returns MakeSolid from BRepBuilderAPI;
    
    Create(S1,S2,S3 : Shell from TopoDS)
	---Purpose: Make a solid from three shells.
	---Level: Public
    returns MakeSolid from BRepBuilderAPI;
    
    	---Purpose: Constructs a solid
    	-- -   covering the whole space, or
    	-- -   from shell S, or
    	-- -   from two shells S1 and S2, or
    	-- -   from three shells S1, S2 and S3, or
    	-- Warning
    	-- No check is done to verify the conditions of coherence
    	-- of the resulting solid. In particular, S1, S2 (and S3) must
    	-- not intersect each other.
    	-- Besides, after all shells have been added using the Add
    	-- function, one of these shells should constitute the outside
    	-- skin of the solid; it may be closed (a finite solid) or open
    	-- (an infinite solid). Other shells form hollows (cavities) in
    	-- these previous ones. Each must bound a closed volume.
        
    ----------------------------------------------
    -- From solid and shells
    ----------------------------------------------

    Create(So : Solid from TopoDS)
	---Purpose: Make a solid from a solid. Usefull for adding later.
	---Level: Public
    returns MakeSolid from BRepBuilderAPI;
    
    Create(So : Solid from TopoDS; S : Shell from TopoDS)
	---Purpose: Add a shell to a solid.
	---Level: Public
    returns MakeSolid from BRepBuilderAPI;
    
    	---Purpose:
    	-- Constructs a solid:
    	-- -   from the solid So, to which shells can be added, or
    	-- -   by adding the shell S to the solid So.
    	--   Warning
    	-- No check is done to verify the conditions of coherence
    	-- of the resulting solid. In particular S must not intersect the solid S0.
    	-- Besides, after all shells have been added using the Add
    	-- function, one of these shells should constitute the outside
    	-- skin of the solid. It may be closed (a finite solid) or open
    	-- (an infinite solid). Other shells form hollows (cavities) in
    	-- the previous ones. Each must bound a closed volume.	
    
    ----------------------------------------------
    -- Auxiliary methods
    ----------------------------------------------

    Add(me : in out; S : Shell from TopoDS)
	---Purpose: Adds the shell to the current solid.
    	--	Warning
    	-- No check is done to verify the conditions of coherence
    	-- of the resulting solid. In particular, S must not intersect
    	-- other shells of the solid under construction.
    	-- Besides, after all shells have been added, one of
    	-- these shells should constitute the outside skin of the
    	-- solid. It may be closed (a finite solid) or open (an
    	-- infinite solid). Other shells form hollows (cavities) in
    	-- these previous ones. Each must bound a closed volume.
    is static;
    
    ----------------------------------------------
    -- Results
    ----------------------------------------------

    IsDone(me) returns Boolean
	---Purpose: Returns true if the solid is built.
    	-- For this class, a solid under construction is always valid.
    	-- If no shell has been added, it could be a whole-space
    	-- solid. However, no check was done to verify the
    	-- conditions of coherence of the resulting solid.
    is redefined;

    Solid(me) returns Solid from TopoDS
	---Purpose: Returns the new Solid.
	--          
	---C++: return const &
	---C++: alias "Standard_EXPORT operator TopoDS_Solid() const;"
 	---Level: Public
    raises
    	NotDone from StdFail
    is static;
 
    IsDeleted (me: in out; S : Shape from TopoDS)
    returns Boolean
    is redefined;

fields  

    myMakeSolid : MakeSolid from BRepLib;

end MakeSolid;
