-- File:	TopoDSToStep_MakeStepFace.cdl
-- Created:	Wed Nov 30 10:14:17 1994
-- Author:	Frederic MAUPAS
--		<fma@bibox>
---Copyright:	 Matra Datavision 1994

class MakeStepFace from TopoDSToStep 
    inherits Root from TopoDSToStep

    ---Purpose: This class implements the mapping between classes 
    --          Face from TopoDS and TopologicalRepresentationItem from
    --          StepShape. 
  
uses Face                          from TopoDS,
     TopologicalRepresentationItem from StepShape,
     Tool                          from TopoDSToStep,
     MakeFaceError                 from TopoDSToStep,
     FinderProcess                 from Transfer
          
raises NotDone from StdFail
     
is 

    Create returns MakeStepFace;
    
    Create (F           : Face from TopoDS;
            T           : in out Tool from TopoDSToStep;
            FP          : mutable FinderProcess from Transfer)
         returns MakeStepFace;
    
    Init(me          : in out;
         F           : Face from TopoDS;
         T           : in out Tool from TopoDSToStep;
         FP          : mutable FinderProcess from Transfer);
	    	    
    Value (me) returns TopologicalRepresentationItem from StepShape
    	raises NotDone
    	is static;
    	---C++: return const&
    
    Error(me) returns MakeFaceError from TopoDSToStep;

fields

    myResult : TopologicalRepresentationItem from StepShape;

    myError  : MakeFaceError from TopoDSToStep;
    
end MakeStepFace;


