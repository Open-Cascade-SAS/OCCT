-- Created on: 1998-10-29
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Hctxee2d from TopOpeBRep inherits TShared from  MMgt

uses

    Shape from TopoDS,
    Edge from TopoDS,
    Surface from BRepAdaptor,
    Face from TopoDS,
    Curve from Geom2dAdaptor,
    CurveType from GeomAbs,
    Domain from IntRes2d
    
is

    Create returns mutable Hctxee2d from TopOpeBRep;
    SetEdges(me:mutable;E1,E2:Edge;BAS1,BAS2:Surface from BRepAdaptor);
    Edge(me;I:Integer) returns Shape;---C++ : return const &
    Curve(me;I:Integer) returns Curve from Geom2dAdaptor; ---C++ : return const &
    Domain(me;I:Integer) returns Domain from IntRes2d; ---C++ : return const &

fields

    myEdge1 : Edge from TopoDS;
    myCurve1 : Curve from Geom2dAdaptor;
    myCurveType1 : CurveType from GeomAbs;
    myDomain1 : Domain from IntRes2d;

    myEdge2 : Edge from TopoDS;
    myCurve2 : Curve from Geom2dAdaptor;
    myCurveType2 : CurveType from GeomAbs;
    myDomain2 : Domain from IntRes2d;

end Hctxee2d from TopOpeBRep;
