-- Created on: 1991-02-20
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



package IntAna2d


    ---Purpose: This package defines the intersection between two elements of
    --          the geometric processor : Line, Circle, Ellipse, Parabola and
    --          Hyperbola; One of these elements is known with his real type,
    --          the other one is known by an implicit quadratic equation (see
    --          class Conic).
    --          A particular case has been made for the intersection between
    --          two Lin2d, two Circ2d, a Lin2d and a Circ2d.

uses

    Standard, TCollection, gp, StdFail

is

    class Conic;

    class AnaIntersection;

    class IntPoint;
     
end IntAna2d;
