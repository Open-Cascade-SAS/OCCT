-- Created on: 1993-06-23
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Point from TopOpeBRepDS

    ---Purpose: A Geom point and a tolerance.

uses

    Pnt from gp,
    Shape from TopoDS
    
is

    Create returns Point from TopOpeBRepDS; 

    Create(P : Pnt from gp; T : Real from Standard)
    returns Point from TopOpeBRepDS; 

    Create(S : Shape from TopoDS)
    returns Point from TopOpeBRepDS;

    IsEqual(me; other : Point from TopOpeBRepDS)
    returns Boolean from Standard
    is static;

    Point(me) returns Pnt from gp
    ---C++: return const &
    is static;
    
    ChangePoint(me : in out) returns Pnt from gp
    ---C++: return &
    is static;
    
    Tolerance(me) returns Real from Standard
    is static;

    Tolerance(me : in out; Tol : Real from Standard)
    is static;

    Keep(me) returns Boolean from Standard
    is static;
    ChangeKeep(me : in out; B : Boolean from Standard)
    is static;

fields

    myPoint     : Pnt from gp;
    myTolerance : Real from Standard;
    myKeep      : Boolean from Standard;
    
end Point from TopOpeBRepDS;
