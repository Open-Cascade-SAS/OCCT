-- Created on: 1993-06-16
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ShellFaceSet from TopOpeBRepBuild 
    inherits ShapeSet from TopOpeBRepBuild

---Purpose: a bound is a shell, a boundelement is a face.
-- The ShapeSet stores :
-- - a list of shell (bounds),
-- - a list of face (boundelements) to start reconstructions,
-- - a map of edge giving the list of face incident to an edge.

uses

    Shape from TopoDS,
    Solid from TopoDS,
    AsciiString from TCollection,
    ListOfShape from TopTools
    
is

    Create returns ShellFaceSet from TopOpeBRepBuild; 
    ---Purpose: Creates a ShellFaceSet to build blocks of faces 
    -- connected by edges.

    Create(S : Shape from TopoDS; Addr : Address from Standard = NULL) 
    returns ShellFaceSet from TopOpeBRepBuild; 
    ---Purpose: Creates a ShellFaceSet to build blocks of faces 
    -- connected by edges.

    Solid(me) returns Solid from TopoDS is static;
    ---C++: return const &

    AddShape(me:in out;S:Shape) is redefined;
    AddStartElement(me:in out;S:Shape) is redefined;
    AddElement(me:in out;S:Shape) is redefined;

    DumpSS(me:in out) is redefined;
    SName(me;S:Shape from TopoDS;sb:AsciiString = "";sa:AsciiString = "")
    returns AsciiString from TCollection is redefined;
    SName(me;S:ListOfShape from TopTools;sb:AsciiString = "";sa:AsciiString = "")
    returns AsciiString from TCollection is redefined;
    SNameori(me;S:Shape;sb:AsciiString = "";sa:AsciiString = "")
    returns AsciiString from TCollection is redefined;
    SNameori(me;S:ListOfShape from TopTools;sb:AsciiString = "";sa:AsciiString = "")
    returns AsciiString from TCollection is redefined;

fields

    mySolid : Solid from TopoDS;

end ShellFaceSet from TopOpeBRepBuild;
