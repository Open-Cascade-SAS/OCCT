-- Created on: 1993-07-27
-- Created by: Jean Louis FRENKEL
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package Image

  ---Purpose: The package Image provides image manipulation classes.

uses

  TCollection,
  TColStd,
  Aspect,
  Quantity,
  gp,
  MMgt

is

  -----------------------------
  ---Category: Imported types:
  -----------------------------

  imported PixMap;
  imported AlienPixMap;
  imported PixMap_Handle;
  imported AlienPixMap_Handle;
  imported Diff;

end Image;
