-- Created on: 1996-05-31
-- Created by: Laurent BUCHARD
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



package IntCurvesFace

----------------------------------------------------------------------
-- This package provide algorithms to  compute the intersection points
-- between a Face [a  Shape] and a set of  curves (The face [shape] is
-- loaded, then for each curve is given to compute the intersection).
-- 
-- Intersector [  ShapeIntersector ] can be  used when the caller have
-- to intersect more than one curve with the face [the shape].
-- 
-- 
-- If there is  only one curve, or  if  the face  has no restrictions,
-- someother algorithms can be called. 
--    
-- see for example the packages : 
-- 
--      ** BRepIntCurveSurface :  ( One Curve   <->   One  Shape )
--      ** IntCurveSurface     :  ( One Curve   <->   One  Surface)
--     
----------------------------------------------------------------------


uses 
    gp              ,
    TopAbs          ,
    TopoDS          ,
    BRepTopAdaptor  ,
    BRepAdaptor     ,
    Adaptor3d         ,
    Bnd             ,
    IntCurveSurface ,
    TColStd         ,
    GeomAbs
    
is

    class Intersector;            -- Intersection between a Face and a set of curves 
    
    class ShapeIntersector;       -- Intersection between a Shape and a set of curves 
                                  -- Note ( has an empty constructor )
    
end;

