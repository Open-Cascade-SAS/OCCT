-- Created on: 1991-01-10
-- Created by: Arnaud BOUZY
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class UnaryExpression from Expr

inherits GeneralExpression from Expr

uses NamedUnknown from Expr

raises OutOfRange from Standard, 
    NumericError from Standard,
    InvalidOperand from Expr

is

    Operand(me)
    ---Purpose: Returns the operand used
    ---C++: inline
    ---C++: return const &
    ---Level : Internal
    returns any GeneralExpression
    is static;

    SetOperand(me : mutable; exp : GeneralExpression)
    ---Purpose: Sets the operand used
    --          Raises InvalidOperand if <exp> contains <me>.
    ---Level : Internal
    raises InvalidOperand
    is static;
    
    CreateOperand(me : mutable; exp : GeneralExpression)
    ---Purpose: Sets the operand used during creation
    ---Level : Internal
    is static protected;
    
    NbSubExpressions(me)
    ---Purpose: Returns the number of sub-expressions contained
    --          in <me> ( >= 0)
    returns Integer
    is static;

    SubExpression(me; I : Integer)
    ---Purpose: Returns the <I>-th sub-expression of <me>.
    --          Raises OutOfRange if <I> > NbSubExpressions(me)
    ---C++: return const &
    returns any GeneralExpression
    raises OutOfRange
    is static;

    ContainsUnknowns(me) 
    ---Purpose: Does <me> contains NamedUnknown ?
    returns Boolean
    is static;

    Contains(me; exp : GeneralExpression)
    ---Purpose: Tests if <exp> is contained in <me>.
    returns Boolean
    is static;

    Replace(me : mutable ; var : NamedUnknown ; with : GeneralExpression)
    ---Purpose: Replaces all occurences of <var> with <with> in <me>
    --          Raises InvalidOperand if <with> contains <me>.
    raises InvalidOperand
    is static;
    
    Simplified(me) 
    ---Purpose: Returns a GeneralExpression after replacement of
    --          NamedUnknowns by an associated expression, and after
    --          values computation.
    returns any GeneralExpression
    raises NumericError;
    
fields

    myOperand : GeneralExpression;

end UnaryExpression;

