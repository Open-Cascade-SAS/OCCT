-- File:	Bisector.cdl
-- Created:	Thu May 19 10:55:33 1994
-- Author:	Yves FRICAUD
--		<yfr@phobox>
---Copyright:	 Matra Datavision 1992

package Bisector 

    --- Purpose : This package provides the bisecting line between two
    --            geometric elements.

uses 
     MMgt,
     Standard,
     TCollection,
     TColStd,	
     TColgp,
     TopAbs,	     
     Geom2d,
     GeomAbs,
     gp,
     math,
     IntCurve,	
     GccInt,
     StdFail,
     IntRes2d
is

    deferred class Curve;
    
   	     class BisecAna;
    	     --- Purpose: This class provides the bisecting line between two
    	     --           geometric elements.The elements are Circles,Lines or
    	     --           Points. 

    	     class BisecPC;
	     ---Purpose: This class provides the bisecting line between a point
	     --          a Curve.
    
    	     class BisecCC;	
	     ---Purpose: This class provides the bisecting line between two
	     --          Curves. 

    class Bisec;
	---Purpose: This class provides the bisecting line between two
	--          geometris  elelements.  The   bisecting   line  is
	--          trimmed by a point, 
    
    class Inter;
    
    class PointOnBis;
    
    class PolyBis;
    
    private class FunctionH;
    
    private class FunctionInter;
    
    IsConvex (Cu : Curve from Geom2d; Sign : Real) 
    returns Boolean from Standard;
    
end Bisector;
