-- Created on: 1993-06-11
-- Created by: Martine LANGLOIS
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package GeomToStep

--- Purpose: Creation des entites geometriques du schema PmsAp2Demo3d a 
--  partir des entites de Geom ou de gp.
--  Update : mise a jour pour traiter le schema StepGeom, pour demo de 94

uses gp, Geom, Geom2d, StepGeom, StdFail, TColgp

is

private deferred class Root;
class MakeCartesianPoint;
class MakeAxis1Placement;
class MakeAxis2Placement2d;
class MakeAxis2Placement3d;
class MakeDirection;
class MakeVector;
class MakeCurve;
class MakeConic;
class MakeBoundedCurve;
class MakeCircle;
class MakeEllipse;
class MakeHyperbola;
class MakeParabola;
class MakeBSplineCurveWithKnots;
class MakeBSplineCurveWithKnotsAndRationalBSplineCurve;
class MakeLine;
class MakePolyline;
class MakePlane;
class MakeSurface;
class MakeBoundedSurface;
class MakeElementarySurface;
class MakeSweptSurface;
class MakeConicalSurface;
class MakeCylindricalSurface;
class MakeRectangularTrimmedSurface;
class MakeSphericalSurface;
class MakeSurfaceOfLinearExtrusion;
class MakeSurfaceOfRevolution;
class MakeToroidalSurface;
class MakeBSplineSurfaceWithKnots;
class MakeBSplineSurfaceWithKnotsAndRationalBSplineSurface;

end GeomToStep;
