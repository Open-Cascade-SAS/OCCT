-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class CurveOnSurface from StepGeom inherits SelectType from StepData

	-- <CurveOnSurface> is an EXPRESS Select Type construct translation.
	-- it gathers : Pcurve, SurfaceCurve, CompositeCurveOnSurface

uses

	Pcurve,
	SurfaceCurve,
	CompositeCurveOnSurface
is

	Create returns CurveOnSurface;
	---Purpose : Returns a CurveOnSurface SelectType

	CaseNum (me; ent : Transient) returns Integer;
	---Purpose: Recognizes a CurveOnSurface Kind Entity that is :
	--        1 -> Pcurve
	--        2 -> SurfaceCurve
	--        3 -> CompositeCurveOnSurface
	--        0 else

	Pcurve (me) returns any Pcurve;
	---Purpose : returns Value as a Pcurve (Null if another type)

	SurfaceCurve (me) returns any SurfaceCurve;
	---Purpose : returns Value as a SurfaceCurve (Null if another type)

	CompositeCurveOnSurface (me) returns any CompositeCurveOnSurface;
	---Purpose : returns Value as a CompositeCurveOnSurface (Null if another type)


end CurveOnSurface;

