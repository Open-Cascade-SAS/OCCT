-- Created on: 2000-08-22
-- Created by: Andrey BETENEV
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class UOperator from ShapeProcess inherits Operator from ShapeProcess

    ---Purpose: Defines operator as container for static function
    --          OperFunc. This allows user to create new operators 
    --          without creation of new classes

uses

    OperFunc from ShapeProcess,
    Context from ShapeProcess

is

    Create (func: OperFunc from ShapeProcess);
    	---Purpose: Creates operator with implementation defined as
	--          OperFunc (static function)

    Perform (me: mutable; context: Context from ShapeProcess) 
    returns Boolean is redefined;
    	---Purpose: Performs operation and records changes in the context

fields

    myFunc: OperFunc from ShapeProcess;

end UOperator;
