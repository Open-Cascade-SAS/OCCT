-- File:        Person.cdl
-- Created:     Mon Dec  4 12:02:28 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWPerson from RWStepBasic

	---Purpose : Read & Write Module for Person

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     Person from StepBasic

is

	Create returns RWPerson;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable Person from StepBasic);

	WriteStep (me; SW : in out StepWriter; ent : Person from StepBasic);

end RWPerson;
