-- Created on: 1998-08-03
-- Created by: Christian CAILLET
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class ToVRML  from SWDRAW

    ---Purpose : Writes a Shape to a File in VRML Format

uses CString, OStream, AsciiString from TCollection, Shape from TopoDS

is

    Create returns ToVRML;

    EmissiveColorRed   (me : in out) returns Real;
    ---C++ : return &
    EmissiveColorGreen (me : in out) returns Real;
    ---C++ : return &
    EmissiveColorBlue  (me : in out) returns Real;
    ---C++ : return &
    DiffuseColorRed    (me : in out) returns Real;
    ---C++ : return &
    DiffuseColorGreen  (me : in out) returns Real;
    ---C++ : return &
    DiffuseColorBlue   (me : in out) returns Real;
    ---C++ : return &
    Transparency       (me : in out) returns Real;
    ---C++ : return &
    AmbientIntensity   (me : in out) returns Real;
    ---C++ : return &
    SpecularColorRed   (me : in out) returns Real;
    ---C++ : return &
    SpecularColorGreen (me : in out) returns Real;
    ---C++ : return &
    SpecularColorBlue  (me : in out) returns Real;
    ---C++ : return &
    Shininess          (me : in out) returns Real;
    ---C++ : return &
    Texture            (me : in out) returns AsciiString;
    ---C++ : return &
    CreaseAngle        (me : in out) returns Real;
    ---C++ : return &
    Deflection         (me : in out) returns Real;
    ---C++ : return &


    Write (me; shape : Shape from TopoDS; filename : CString) returns Boolean;
    ---Purpose : conversion of a Shape into VRML format for 3d visualisation

fields

  myEmissiveColorRed   : Real;  -- def 0.3
  myEmissiveColorGreen : Real;  -- def 0.3
  myEmissiveColorBlue  : Real;  -- def 0.3
  myDiffuseColorRed    : Real;  -- def 0.3
  myDiffuseColorGreen  : Real;  -- def 0.3
  myDiffuseColorBlue   : Real;  -- def 0.5
  myTransparency       : Real;  -- def 0.0
  myAmbientIntensity   : Real;  -- def 0.3
  mySpecularColorRed   : Real;  -- def 0.7
  mySpecularColorGreen : Real;  -- def 0.7
  mySpecularColorBlue  : Real;  -- def 0.8
  myShininess          : Real;  -- def 0.1
  myTexture            : AsciiString;  -- def " [] "
  myCreaseAngle        : Real;  -- def 1.57
  myDeflection         : Real;  -- def 0.005

end ToVRML;
