-- Created on: 1992-02-20
-- Created by: Remy GILET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

generic class FunctionTanCirCu from GccIter (
    TheCurve     as any;
    TheCurveTool as any) -- as CurvePGTool from GccInt(TheCurve)

inherits FunctionWithDerivative from math
         
    ---Purpose: This abstract class describes a Function of 1 Variable 
    --          used to find a line tangent to a curve and a circle.

uses Circ2d from gp    

is

Create (Circ   : Circ2d   from gp ;
    	Curv   : TheCurve         ) returns FunctionTanCirCu from GccIter;

Value (me : in out      ;
       X  :        Real ;
       F  :    out Real ) returns Boolean;
    ---Purpose: Computes the value of the function F for the variable X.
    --          It returns True if the computation is successfully done,
    --          False otherwise.

Derivative (me    : in out      ;
            X     :        Real ;
            Deriv :    out Real ) returns Boolean;
    ---Purpose: Computes the derivative of the function F for the variable X.
    --          It returns True if the computation is successfully done,
    --          False otherwise.

Values (me    : in out      ;
        X     :        Real ;
        F     : out    Real ;
        Deriv : out    Real ) returns Boolean;
    ---Purpose: Computes the value and the derivative of the function F 
    --          for the variable X.
    --          It returns True if the computation is successfully done,
    --          False otherwise.

fields

TheCirc  : Circ2d from gp;
Curve    : TheCurve; 
-- Modified by Sergey KHROMOV - Thu Apr  5 09:50:18 2001 Begin
myWeight : Real;
-- Modified by Sergey KHROMOV - Thu Apr  5 09:50:19 2001 End

end FunctionTanCirCu;
