-- Created on: 1993-01-11
-- Created by: CKY / Contract Toubro-Larsen ( Anand NATRAJAN )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class NodalConstraint from IGESAppli  inherits IGESEntity

        ---Purpose: defines NodalConstraint, Type <418> Form <0>
        --          in package IGESAppli
        --          Relates loads and/or constraints to specific nodes in
        --          the Finite Element Model by creating a relation between
        --          Node entities and Tabular Data Property that contains
        --          the load or constraint data

uses

        TabularData          from IGESDefs,
        Node                 from IGESAppli,
        HArray1OfTabularData from IGESDefs

raises OutOfRange

is

        Create returns mutable NodalConstraint;

        -- Specific Methods pertaining to the class

        Init (me         : mutable;
              aType      : Integer;
              aNode      : Node;
              allTabData : HArray1OfTabularData);
        ---Purpose : This method is used to set the fields of the class
        --           NodalConstraint
        --       - aType      : Loads / Constraints
        --       - aNode      : the Node
        --       - allTabData : Tabular Data Property carrying the load
        --                      or constraint vector

        NbCases (me) returns Integer;
        ---Purpose : returns total number of cases

        Type (me) returns Integer;
        ---Purpose : returns whether Loads (1) or Constraints (2)

        NodeEntity (me) returns Node;
        ---Purpose : returns the Node

        TabularData (me; Index : Integer) returns TabularData
        raises OutOfRange;
        ---Purpose : returns Tabular Data Property carrying load or constraint vector
        -- raises exception if Index <= 0 or Index > NbCases

fields

--
-- Class    : IGESAppli_NodalConstraint
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class NodalConstraint.
--
-- Reminder : A NodalConstraint instance is defined by :
--            - indicator whether Loads or Constraints
--            - a Node
--            - Tabular Data Property carrying load or constraint vector

        theType             : Integer;
        theNode             : Node;
        theTabularDataProps : HArray1OfTabularData;

end NodalConstraint;
