-- Created on: 2000-08-11
-- Created by: Andrey BETENEV
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class AISObject from XCAFPrs inherits Shape from AIS

    ---Purpose: Implements AIS_InteractiveObject functionality
    --          for shape in DECAF document

uses
    Shape from TopoDS,
    PresentationManager3d from PrsMgr,
    Presentation from Prs3d,
    Label from TDF,
    Color from Quantity,
    NameOfMaterial from Graphic3d,
    MaterialAspect from Graphic3d,
    Style from XCAFPrs
    
is

    Create (lab: Label from TDF);
    	---Purpose: Creates an object to visualise the shape label

    SetColor(me:mutable;aColor:Color from Quantity) is redefined virtual;

    UnsetColor(me:mutable) is redefined virtual;
        
    SetMaterial(me:mutable;aName:NameOfMaterial from Graphic3d) is redefined virtual;

    SetMaterial(me:mutable;aName:MaterialAspect from Graphic3d) is redefined virtual;
        
    UnsetMaterial(me:mutable) is redefined virtual;
        
    SetTransparency(me:mutable;aValue : Real from Standard=0.6) is redefined virtual;  
    
    UnsetTransparency(me:mutable) is redefined virtual;
 
    AddStyledItem (me: mutable; style: Style from XCAFPrs;
                   shape: Shape from TopoDS;
                   aPresentationManager : PresentationManager3d from PrsMgr;
                   aPresentation        : mutable Presentation from Prs3d;
    	           aMode                : Integer from Standard = 0) 
    is private;

    Compute (me                   : mutable;
             aPresentationManager : PresentationManager3d from PrsMgr;
             aPresentation        : mutable Presentation from Prs3d;
    	     aMode                : Integer from Standard = 0) 
    is redefined virtual protected;
    	---Purpose: Redefined method to compute presentation

    DefaultStyle (me;
                  aStyle: out Style from XCAFPrs)
    is virtual protected;
    ---Purpose: Fills out a default style object which is used when styles are
    --          not explicitly defined in the document.
    --          By default, the style uses white color for curves and surfaces.

fields
    myLabel : Label from TDF;

end AISObject;
