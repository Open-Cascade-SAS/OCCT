-- File:	MeshAlgo_CircleTool.cdl
-- Created:	Wed May 12 09:30:49 1993
-- Author:	Didier PIFFAULT
--		<dpf@zerox>
---Copyright:	 Matra Datavision 1993


class CircleTool from MeshAlgo 

	---Purpose: Create sort   and  destroy the  circles    used in
	--          triangulation.

uses    Boolean from Standard,
    	Integer from Standard,
    	Real from Standard,
    	XY from gp,
    	Circ2d from gp,
	ListOfInteger from MeshDS,
        CellFilter from MeshAlgo,
	CircleInspector from MeshAlgo,
	BaseAllocator from MeshDS

is      Create (theAlloc : in BaseAllocator from MeshDS)
        returns CircleTool from MeshAlgo;


    	Create     (numberOfComponents : in Integer from Standard;
    	    	    theAlloc : in BaseAllocator from MeshDS)
	---Purpose: Constructs a CircleTool with the maximal dimension
	--          of  the occuped  space and  an  evaluation of  the
	--          number of circles.
    	    returns CircleTool from MeshAlgo;

    	Initialize (me                 : in out;
    	    	    numberOfComponents : in Integer from Standard)
	---Purpose: Constructs a CircleTool with the maximal dimension
	--          of  the occuped  space and  an  evaluation of  the
	--          number of circles.
    	    is static;

        SetCellSize(me                 : in out;
    	    	    theSize            : in Real from Standard)
	---Purpose: Sets new size for cellfilter
       	    is static;

        SetCellSize(me                 : in out;
    	    	    theXSize            : in Real from Standard;
                    theYSize            : in Real from Standard)
	---Purpose: Sets new size for cellfilter
       	    is static;

        SetMinMaxSize(me                 : in out;
    	    	      theMin             : in XY from gp;
                      theMax             : in XY from gp)
	---Purpose: Sets min and max size for circle
       	    is static;

    	Add      (me       : in out;
    	    	  theCirc  : in Circ2d from gp;
    	    	  theIndex : in Integer from Standard)
	---Purpose: Adds and binds circle to the tool.
    	    is static;


    	Add      (me          : in out;
    	    	  p1, p2, p3  : in XY from gp;
    	    	  theIndex    : in Integer from Standard)
	---Purpose: Computes adds and binds circle to the tool.
    	    returns Boolean from Standard is static;
	
	MocAdd   (me          : in out;
	    	  theIndex    : in Integer from Standard);
	---Purpose: Adds implicit zero circle


    	Delete   (me : in out; theIndex : Integer from Standard) 
	---Purpose: Deletes a circle from the tool.
    	    is static;


    	Select   (me : in out; thePnt : XY from gp)
	---Purpose: Select the circles which contains thePnt.
	---C++: return &
	    returns ListOfInteger from MeshDS is static;
	    
fields  Tolerance    : Real from Standard;
        Allocator    : BaseAllocator from MeshDS;
	CellFilter   : CellFilter from MeshAlgo;
        Selector     : CircleInspector from MeshAlgo;
	FaceMax      : XY from gp;
	FaceMin      : XY from gp;

end CircleTool;
