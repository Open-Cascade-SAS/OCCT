-- File     : Prs2d_Repere.cdl
-- Created  : October  2000
-- Author   : Tanya COOL
---Copyright: Matra Datavision 2000

class Repere from Prs2d inherits Dimension from Prs2d

 ---Purpose: Constructs the repere

uses

	Drawer		       from Graphic2d,
	GraphicObject	   from Graphic2d,
	Pnt2d              from gp,
	ExtendedString     from TCollection,
	Array1OfShortReal  from TShort,
    	ArrowSide          from Prs2d,
	TypeOfArrow        from Prs2d,
    	FStream            from Aspect 

is
	Create( aGO           : GraphicObject  from Graphic2d;
	        aPnt1         : Pnt2d          from gp;
            	aPnt2         : Pnt2d          from gp;
		aLenBase      : Real           from Standard; 
		aText         : ExtendedString from TCollection;
       	    	aTxtScale     : Real           from Standard = 1.0;
            	aDrawArrow    : Boolean        from Standard = Standard_False; 
            	anArrAngle    : Real           from Standard = 10.0;
		anArrLength   : Real           from Standard = 10.0;
            	anArrType     : TypeOfArrow    from Prs2d    = Prs2d_TOA_OPENED;
		anArrow       : ArrowSide      from Prs2d    = Prs2d_AS_BOTHAR;
		IsRevArrow    : Boolean        from Standard = Standard_False ) 

	returns mutable Repere from Prs2d;
    	---Level: Public
    	---Purpose: Creates repere 

	-------------------------------------------------
	-- Category: Draw and Pick
	-------------------------------------------------

	Draw( me : mutable; aDrawer: Drawer from Graphic2d ) is static protected;
	---Level: Internal
	---Purpose: Draws the repere <me>.

    	DrawElement( me : mutable; aDrawer: Drawer from Graphic2d;
            	     anIndex: Integer from Standard)
            is redefined protected;
    	---Level: Internal
    	---Purpose: 

    	DrawVertex( me : mutable; aDrawer: Drawer from Graphic2d;
                    anIndex: Integer from Standard)
            is redefined protected;
    	---Level: Internal
    	---Purpose: 

    	Pick( me : mutable; X, Y: ShortReal from Standard;
       	      aPrecision: ShortReal from Standard;
	      aDrawer: Drawer from Graphic2d ) 
    	returns Boolean from Standard is static protected;
	---Level: Internal
	---Purpose: Returns Standard_True if the repere <me> is picked,
	--	    Standard_False if not.

	Save( me; aFStream: in out FStream from Aspect ) is virtual;
													
    	CalcTxtPos(me:mutable; theFromAbs: 
    	    	    Boolean from Standard) 
    	---C++: inline
    	is redefined protected;

fields 
 
    myXVert        : Array1OfShortReal from TShort;
    myYVert        : Array1OfShortReal from TShort;
    myObtuse       : Boolean           from Standard;
    myDrawArrow    : Boolean           from Standard;

end Repere from Prs2d;
