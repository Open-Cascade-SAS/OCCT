-- File:	IGESBasic_ToolName.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolName  from IGESBasic

    ---Purpose : Tool to work on a Name. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses Name from IGESBasic,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolName;
    ---Purpose : Returns a ToolName, ready to work


    ReadOwnParams (me; ent : mutable Name;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : Name;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : Name;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a Name <ent>, from
    --           its specific (own) parameters

    OwnCorrect (me; ent : mutable Name) returns Boolean  is static;
    ---Purpose : Sets automatic unambiguous Correction on a Name
    --           (NbPropertyValues forced to 1)

    DirChecker (me; ent : Name) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : Name;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : Name; entto : mutable Name;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : Name;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolName;
