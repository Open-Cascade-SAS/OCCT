-- Created on: 1992-10-02
-- Created by: Christian CAILLET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class AllConnected  from IFGraph  inherits GraphContent

    	---Purpose : this class gives content of the CONNECTED COMPONANT(S)
    	--           which include specific Entity(ies)

uses Transient, EntityIterator, Graph

is

    Create (agraph : Graph) returns AllConnected;
    ---Purpose : creates an AllConnected from a graph, empty ready to be filled

    Create (agraph : Graph; ent : any Transient)
    	returns AllConnected;
    ---Purpose : creates an AllConnected which memorizes Entities Connected to
    --           a given one, at any level : that is, itself, all Entities
    --           Shared by it and Sharing it, and so on.
    --           In other terms, this is the content of the CONNECTED COMPONANT
    --           which include a specific Entity

    GetFromEntity (me : in out; ent : any Transient);
    ---Purpose : adds an entity and its Connected ones to the list (allows to
    --           cumulate all Entities Connected by some ones)
    --           Note that if "ent" is in the already computed list,, no entity
    --           will be added, but if "ent" is not already in the list, a new
    --           Connected Componant will be cumulated 

    ResetData (me : in out);
    ---Purpose : Allows to restart on a new data set

    	-- --   Results   -- --
    	--   More-Next-Value give all entities noted in Connected Componant,
    	--   including the entities given for construction or to GetFromEntity

    Evaluate (me : in out) is redefined;
    ---Purpose : does the specific evaluation (Connected entities atall levels)

fields

    thegraph : Graph;

end AllConnected;
