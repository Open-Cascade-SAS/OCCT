-- Created on: 1994-03-25
-- Created by: Jean Marc LACHAUME
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class IsoBuilder from DBRep

	---Purpose: Creation of isoparametric curves.

inherits Hatcher from Geom2dHatch

uses

    Face from TopoDS ,
    Face from DBRep ,
    Array1OfReal    from TColStd ,
    Array1OfInteger from TColStd
    

is

    Create (TopologicalFace : Face    from TopoDS ;
    	    Infinite        : Real    from Standard ;
    	    NbIsos          : Integer from Standard)

    	---Purpose: Creates the builder.

    	returns IsoBuilder from DBRep ;


    NbDomains (me)

    	---Purpose: Returns the total number of domains.

    	---C++: inline

    	returns Integer from Standard
    	is static ;


    LoadIsos (me; Face : mutable Face from DBRep)

    	---Purpose: Loading of the isoparametric curves in the
    	--          Data Structure of a drawable face.

    	is static ;


fields

    myInfinite : Real            from Standard ;
    myUMin     : Real            from Standard ;
    myUMax     : Real            from Standard ;
    myVMin     : Real            from Standard ;
    myVMax     : Real            from Standard ;
    myUPrm     : Array1OfReal    from TColStd ;
    myUInd     : Array1OfInteger from TColStd ;    
    myVPrm     : Array1OfReal    from TColStd ;
    myVInd     : Array1OfInteger from TColStd ;    
    myNbDom    : Integer         from Standard ;
    
end IsoBuilder;
