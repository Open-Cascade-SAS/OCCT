-- File:	TColGeom2d.cdl
-- Created:	Thu Apr 15 12:11:39 1993
-- Author:	Philippe DAUTRY
--		<fid@mastox>
-- Copyright:	 Matra Datavision 1993


package TColGeom2d


        ---Purpose : 
-- The package TColGeom2d provides standard and
-- frequently used instantiations of generic classes from
-- the TCollection package with geometric objects from the Geom2d package.

uses TCollection, Geom2d

is


    class Array1OfGeometry 
    	instantiates Array1 from TCollection (Geometry from Geom2d);
    class Array1OfCurve 
    	instantiates Array1 from TCollection (Curve from Geom2d);
    class Array1OfBoundedCurve 
    	instantiates Array1 from TCollection (BoundedCurve from Geom2d);
    class Array1OfBezierCurve 
    	instantiates Array1 from TCollection (BezierCurve from Geom2d);
    class Array1OfBSplineCurve 
    	instantiates Array1 from TCollection (BSplineCurve from Geom2d);

    class HArray1OfGeometry
    	instantiates HArray1 from TCollection (Geometry from Geom2d,
    	    	    	    	Array1OfGeometry from TColGeom2d);
    class HArray1OfCurve
    	instantiates HArray1 from TCollection (Curve from Geom2d,
    	    	    	    	Array1OfCurve from TColGeom2d);
    class HArray1OfBoundedCurve 
    	instantiates HArray1 from TCollection (BoundedCurve from Geom2d,
    	    	    	    	Array1OfBoundedCurve from TColGeom2d);
    class HArray1OfBezierCurve  
    	instantiates HArray1 from TCollection (BezierCurve from Geom2d,
    	    	    	    	Array1OfBezierCurve from TColGeom2d);
    class HArray1OfBSplineCurve 
    	instantiates HArray1 from TCollection (BSplineCurve from Geom2d,
    	    	    	    	Array1OfBSplineCurve from TColGeom2d);


    class SequenceOfGeometry  
    	instantiates Sequence from TCollection (Geometry from Geom2d);
    class SequenceOfCurve  
    	instantiates Sequence from TCollection (Curve from Geom2d);
    class SequenceOfBoundedCurve  
    	instantiates Sequence from TCollection (BoundedCurve from Geom2d);

    class HSequenceOfGeometry  
    	instantiates HSequence from TCollection (Geometry from Geom2d,
    	    	    	    	SequenceOfGeometry from TColGeom2d);
    class HSequenceOfCurve  
    	instantiates HSequence from TCollection (Curve from Geom2d,
    	    	    	    	SequenceOfCurve from TColGeom2d);
    class HSequenceOfBoundedCurve  
    	instantiates HSequence from TCollection (BoundedCurve from Geom2d,
    	    	    	    	SequenceOfBoundedCurve from TColGeom2d);


end TColGeom2d;
