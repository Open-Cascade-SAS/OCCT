-- Created on: 1992-10-22
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



generic class PathPoint from IntStart
    (TheVertex as any;
     TheArc    as any)

	---Purpose: This class describes a point on an arc which
	--          solution intersection between 2 surfaces.

uses Pnt          from gp,
     Vec          from gp,
     Dir2d        from gp

raises DomainError from Standard

is

    Create
    
	returns PathPoint from IntStart;


    Create(P: Pnt from gp; Tol: Real from Standard;
           V: TheVertex; A: TheArc; Parameter: Real from Standard)

    	returns PathPoint from IntStart;
	

    Create(P: Pnt from gp; Tol: Real from Standard;
           A: TheArc; Parameter: Real from Standard)
	
	returns PathPoint from IntStart;


    SetValue(me: in out; P: Pnt from gp; Tol: Real from Standard;
                         V: TheVertex; A: TheArc;
                         Parameter: Real from Standard)

	---C++: inline
    
    	is static;


    SetValue(me: in out; P: Pnt from gp; Tol: Real from Standard;
                         A: TheArc; Parameter: Real from Standard)
	
	---C++: inline
    
	is static;


    Value(me)
    
    	returns Pnt from gp
	---C++: return const&
	---C++: inline
    
	is static;


    Tolerance(me)
    
    	returns Real from Standard
	---C++: inline
    
	is static;


    IsNew(me)
    
    	returns Boolean from Standard
	---C++: inline
    
	is static;
    

    Vertex(me)
    
    	returns any TheVertex
	---C++: return const&
	---C++: inline
    
	raises DomainError from Standard
	is static;


    Arc(me)
    
    	returns any TheArc
	---C++: return const&
	---C++: inline
    
	is static;


    Parameter(me)
    
    	returns Real        from Standard
	---C++: inline
    
	raises  DomainError from Standard
	is static;

fields

    point : Pnt          from gp;
    tol   : Real         from Standard;
    isnew : Boolean      from Standard;
    vtx   : TheVertex;
    arc   : TheArc;
    param : Real         from Standard;

end PathPoint;
