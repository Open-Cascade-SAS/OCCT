-- Created on: 1993-04-26
-- Created by: Jean-Louis Frenkel
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

--   GG  : GER61351 17/11/1999 Change SetColor() with a compatible Quantity_Color instead
--				       the restricted NameOfColor.


class IsoAspect from Prs3d inherits LineAspect from Prs3d
    	---Purpose: A framework to define the display attributes of isoparameters.
    	-- This framework can be used to modify the default
    	-- setting for isoparameters in AIS_Drawer.
        
uses 

    NameOfColor from Quantity,
    Color from Quantity,
    TypeOfLine from Aspect

is
    Create (aColor: NameOfColor from Quantity;
	    aType: TypeOfLine from Aspect;
    	    aWidth: Real from Standard;
          aNumber: Integer from Standard)    
	    returns mutable IsoAspect from Prs3d;
    	---Purpose: Constructs a framework to define display attributes of isoparameters.
    	-- These include:
    	-- -   the color attribute aColor
    	-- -   the type of line aType
    	-- -   the width value aWidth
    	-- -   aNumber, the number of isoparameters to be   displayed.
        
    Create (aColor: Color from Quantity;
	    aType: TypeOfLine from Aspect;
    	    aWidth: Real from Standard;
          aNumber: Integer from Standard)	    
	    returns mutable IsoAspect from Prs3d;
	    

    SetNumber (me: mutable; aNumber: Integer from Standard) 
    	---Purpose: defines the number of U or V isoparametric curves 
    	--         to be drawn for a single face.
    	--          Default value: 10
    is static;

    Number (me) returns Integer from Standard 
    	---Purpose: returns the number of U or V isoparametric curves drawn for a single face.
    is static;
    
fields

    myNumber: Integer from Standard;
    
end IsoAspect from Prs3d;
