-- Created on: 1997-09-18
-- Created by: Christophe MARION
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class BiPoint from BRepMesh

uses
    Address from Standard,
    Real    from Standard,
    Integer from Standard
    
is
    Create
    returns BiPoint from BRepMesh; 
    	---C++: inline
    
    Create(X1,Y1,X2,Y2 : Real    from Standard)
    returns BiPoint from BRepMesh; 
    
    Indices(me) returns Address from Standard
    	---C++: inline
    is static;

    Coordinates(me) returns Address from Standard
    	---C++: inline
    is static;

fields
    myIndices     : Integer from Standard[2];
    myCoordinates : Real    from Standard[6];
    
end BiPoint;
