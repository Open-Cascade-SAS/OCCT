-- Created on: 1997-07-31
-- Created by: Denis PASCAL
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Name from PDataStd inherits Attribute from PDF

uses HExtendedString from PCollection

is

    Create returns mutable Name from  PDataStd;
    
    
    Create (V : HExtendedString from PCollection) 
    returns mutable Name from PDataStd;
    
    
    Get (me) returns HExtendedString from PCollection;
    
    
    Set (me : mutable; V : HExtendedString from PCollection);

    
fields

    myValue : HExtendedString from PCollection;

end Name;
