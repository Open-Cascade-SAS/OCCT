-- Created on: 1997-08-26
-- Created by: Stepan MISHIN
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ApproxSurface from GeomConvert 

        ---Purpose: A framework to convert a surface to a BSpline
    	-- surface. This is done by approximation to a BSpline
    	-- surface within a given tolerance.
        
uses 

    Pnt             from gp,
    Surface         from Geom,
    OffsetSurface   from Geom,
    BSplineSurface  from Geom, 
    HSurface        from Adaptor3d,
    Shape           from GeomAbs,     
    ApproxAFunc2Var from AdvApp2Var, 
    OutOfRange      from Standard 
    
raises OutOfRange from Standard

is
    
    Create(Surf: Surface from Geom;
    	   Tol3d: Real; 
           UContinuity : Shape from GeomAbs;
           VContinuity : Shape from GeomAbs;
           MaxDegU : Integer;
       	   MaxDegV : Integer;	   
    	   MaxSegments: Integer; 
	   PrecisCode : Integer) returns ApproxSurface ;
    	---Purpose: Constructs a surface approximation framework defined by
    	-- -   the conic Surf
    	-- -   the tolerance value Tol3d
    	-- -   the degree of continuity UContinuity, VContinuity
    	--  in the directions of the U and V parameters
    	-- -   the highest degree MaxDegU, MaxDegV which
    	--   the polynomial defining the BSpline curve may
    	--   have in the directions of the U and V parameters
    	-- -   the maximum number of segments MaxSegments
    	--   allowed in the resulting BSpline curve
    	-- -   the index of precision PrecisCode.  
    
    Create(Surf:        HSurface from Adaptor3d;
           Tol3d:       Real;
           UContinuity: Shape from GeomAbs;
           VContinuity: Shape from GeomAbs;
           MaxDegU:     Integer;
           MaxDegV:     Integer;
           MaxSegments: Integer;
           PrecisCode : Integer) returns ApproxSurface ;
        ---Purpose: Constructs a surface approximation framework defined by
        -- -   the Surf
        -- -   the tolerance value Tol3d
        -- -   the degree of continuity UContinuity, VContinuity
        --  in the directions of the U and V parameters
        -- -   the highest degree MaxDegU, MaxDegV which
        --   the polynomial defining the BSpline curve may
        --   have in the directions of the U and V parameters
        -- -   the maximum number of segments MaxSegments
        --   allowed in the resulting BSpline curve
        -- -   the index of precision PrecisCode.  


    Surface(me)   returns BSplineSurface from Geom;
    	---Purpose: Returns the BSpline surface resulting from the approximation algorithm.
    

    IsDone(me)    returns  Boolean  from  Standard; 
    	--- Purpose: Returns Standard_True if the approximation has be done
      
    HasResult(me) returns Boolean;
    	--- Purpose: Returns true if the approximation did come out with a result that
    	--  is not NECESSARILY within the required tolerance or a result
    	--  that is not recognized with the wished continuities. 
    
    MaxError(me)  returns Real  from  Standard;
    	--- Purpose: Returns the greatest distance between a point on the
    	-- source conic surface and the BSpline surface
    	-- resulting from the approximation (>0 when an approximation
        --   has been done, 0 if no  approximation )
     
    Dump(me ; o : in out OStream);
    	---Purpose: Prints on the stream o informations on the current state of the object.

    Approximate(me: in out; 
                theSurf:        HSurface from Adaptor3d;
                theTol3d:       Real;
                theUContinuity: Shape from GeomAbs;
                theVContinuity: Shape from GeomAbs;
                theMaxDegU:     Integer;
                theMaxDegV:     Integer;
                theMaxSegments: Integer;
                thePrecisCode : Integer) is private;
        ---Purpose: Converts a surface to B-spline
             
fields
 
    myIsDone   : Boolean         from Standard; 
    myHasResult: Boolean         from Standard; 
    myBSplSurf : BSplineSurface  from Geom; 
    myMaxError : Real            from Standard;
end;
