-- Created on: 1996-10-17
-- Created by: Odile OLIVIER
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SensitiveWire   from Select3D 
inherits SensitiveEntity from Select3D

	---Purpose: A framework to define selection of a wire owner by an
    	-- elastic wire band.

uses
    Pnt                      from gp,
    Projector                from Select3D,
    Lin                      from gp,
    EntityOwner              from SelectBasics,
    SensitiveEntity          from Select3D,
    SensitiveEntitySequence  from Select3D,
    ListOfBox2d              from SelectBasics,
    PickArgs                 from SelectBasics,
    Array1OfPnt2d            from TColgp,
    Box2d                    from Bnd,
    Location                 from TopLoc

is


    Create (OwnerId      : EntityOwner from SelectBasics;
    	    MaxRect      : Integer = 1)
     returns mutable SensitiveWire;
    	---Purpose: Constructs a sensitive wire object defined by the
    	-- owner OwnerId, and the maximum number of
    	-- sensitive rectangles MaxRect.
    Add (me   :mutable;aSensitive : SensitiveEntity from Select3D)
    is static;
    	---Purpose: Adds the sensitive entity aSensitive to this framework.
    Project (me:mutable;aProjector : Projector from Select3D) 
    is redefined static;
    	---Level: Public 
    	---Purpose: projection of the sensitive primitive in order to
    	--          get 2D boxes for the Sort Algorithm

    Areas   (me:mutable ; boxes : in out ListOfBox2d from SelectBasics) 
    is redefined static;
    	---Level: Public 
    	---Purpose: gives the 2D boxes which represent the segment in the 
    	--          selection process...

    GetConnected(me:mutable;aLocation: Location from TopLoc)
    returns SensitiveEntity from Select3D is redefined static;

    GetEdges(me       : mutable;
	     theEdges : in out SensitiveEntitySequence from Select3D);
	---Level: Public
    	---Purpose: returns the sensitive edges stored in this wire


    SetLocation(me:mutable;aLoc:Location from TopLoc) is redefined static;
    	---Purpose:  propagation of location on all the sensitive inside...
    ResetLocation(me:mutable) is redefined static;
    	---Purpose:  propagation of location on all the sensitive inside...    

    Matches (me : mutable;
             thePickArgs : PickArgs from SelectBasics;
             theMatchDMin, theMatchDepth : out Real from Standard)
    returns Boolean
    is redefined static;
    ---Level: Public
    ---Purpose: Checks whether the sensitive entity matches the picking
    -- detection area (close to the picking line).
    -- For details please refer to base class declaration.

    Matches (me  :mutable; 
             XMin,YMin,XMax,YMax : Real from Standard;
             aTol: Real from Standard) 
    returns Boolean
    is static;
     
    Matches (me  :mutable; 
             Polyline:Array1OfPnt2d from TColgp;
	     aBox:Box2d from Bnd;
             aTol: Real from Standard) 
    returns Boolean
    is redefined virtual;
    	---Level: Public 
    

    MaxBoxes(me) returns Integer is redefined static;    
    	---Level: Public 
    	---Purpose:returns <mymaxrect>
	    
    
    Dump(me; S: in out OStream;FullDump : Boolean from Standard = Standard_True) is redefined virtual; 

    Set(me:mutable;TheOwnerId: EntityOwner from SelectBasics) is redefined static; 
    ---Purpose: Sets the owner for all entities in wire 

    GetLastDetected(me)
    returns SensitiveEntity from Select3D is static; 
    ---Purpose:returns <mymaxrect>

fields
    mysensitive     : SensitiveEntitySequence from Select3D;
    myDetectedIndex : Integer from Standard;
end SensitiveWire;








