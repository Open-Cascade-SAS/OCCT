-- Created on: 1993-06-23
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class FaceBuilder from BRepPrim 

	---Purpose: The  FaceBuilder is an algorithm   to build a BRep
	--          Face from a Geom Surface.
	--          
	--          The  face covers  the  whole surface or  the  area
	--          delimited by UMin, UMax, VMin, VMax

uses
    Surface from Geom,
    Face    from TopoDS,
    Edge    from TopoDS,
    Vertex  from TopoDS,
    Builder from BRep

raises
    ConstructionError from Standard,
    OutOfRange from Standard

is
    Create returns FaceBuilder from BRepPrim;

    Create(B : Builder from BRep;
    	   S : Surface from Geom) returns FaceBuilder from BRepPrim;

    Create(B : Builder from BRep;
    	   S : Surface from Geom;
	   UMin, UMax, VMin, VMax : Real) returns FaceBuilder from BRepPrim 
    raises ConstructionError from Standard; -- if UV are outside the  surface
    
    Init(me : in out;
    	   B : Builder from BRep;
    	   S : Surface from Geom)
    is static;
    
    Init(me : in out;
    	   B : Builder from BRep;
    	   S : Surface from Geom;
	   UMin, UMax, VMin, VMax : Real)
    raises ConstructionError from Standard -- if UV are outside the  surface 
    is static;
    
    Face(me) returns Face from TopoDS
	---C++: return const &
	--      
	---C++: alias "Standard_EXPORT operator TopoDS_Face();"
    is static;
    
    Edge(me; I : Integer) returns Edge from TopoDS
	---Purpose: Returns the edge of index <I>
	--          1 - Edge VMin
	--          2 - Edge UMax
	--          3 - Edge VMax
	--          4 - Edge UMin
	--          
	---C++: return const &
    raises OutOfRange from Standard -- if I < 1 or I > 4
    is static;	
    
    Vertex(me; I : Integer) returns Vertex from TopoDS
	---Purpose: Returns the vertex of index <I>
	--          1 - Vertex UMin,VMin
	--          2 - Vertex UMax,VMin
	--          3 - Vertex UMax,VMax
	--          4 - Vertex UMin,VMax
	--          
	---C++: return const &
    raises OutOfRange from Standard -- if I < 1 or I > 4
    is static;	
    

fields
    myVertex : Vertex from TopoDS [4];
    myEdges  : Edge   from TopoDS [4];
    myFace   : Face   from TopoDS;

end FaceBuilder;
