-- File:	RWStepBasic_RWGroup.cdl
-- Created:	Wed May 10 15:09:07 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class RWGroup from RWStepBasic

    ---Purpose: Read & Write tool for Group

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    Group from StepBasic

is
    Create returns RWGroup from RWStepBasic;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : Group from StepBasic);
	---Purpose: Reads Group

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: Group from StepBasic);
	---Purpose: Writes Group

    Share (me; ent : Group from StepBasic;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWGroup;
