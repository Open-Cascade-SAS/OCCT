
-- File:	Graphic2d_SetOfMarkers.cdl
-- Created:	Thu April 13 16:36:51 1993
-- Author:	Gerard GRAS
--		<gg@stylox>
-- Modified: TCL G002A, 28-11-00, is modified method Values(...)

---Copyright:	 Matra Datavision 1993

class SetOfMarkers from Graphic2d inherits Line from Graphic2d

	---Version:

	---Purpose: The primitive SetOfMarkers
	--  Warning: This primitive must be use as possible for performance
	--	   improvment but is drawn with a global marker attributes
	--	   for all the set.
	--	   NOTE: than the method PickedIndex() permits to known
	--	        the last picked marker in the set.
    	--      SAV : 14/11/01 : Added a set of methods (marked SAV before declaration)
    	--                       to provide highlighting/selection
    	--                       of SetOfMarkers elements. These methods should be redefined
    	--                       for other SetOf<>.
    	--                       
    	--      SAV : 23/05/02 : WARNING!!! method PickByCircle performs only detection
    	--      function. It doesn't cause any visual highlighting.

uses

	Drawer			from Graphic2d,
	GraphicObject		from Graphic2d,
	Length			from Quantity,
	PlaneAngle		from Quantity,
	SequenceOfInteger	from TColStd,
	SequenceOfShortReal	from TShort,
	FStream			from Aspect,
	IFStream		from Aspect,
	PickMode                from Graphic2d,
	MapOfInteger            from TColStd,
	HSequenceOfInteger      from TColStd,
	HArray1OfShortReal      from TShort

raises
	MarkerDefinitionError	from Graphic2d,
	OutOfRange from Standard

is
	-------------------------
	-- Category: Constructors
	-------------------------

	Create (aGraphicObject: GraphicObject from Graphic2d)
	returns mutable SetOfMarkers from Graphic2d;
	---Level: Public
	---Purpose: Creates an empty set of markers in the graphic 
	--         object <aGraphicObject>.
	---Category: Constructors

	Add(me : mutable; X, Y: Length from Quantity);
	---Level: Public
	---Purpose: Add a pixel point marker in the set 
	---Category: Update method

	Add(me : mutable; 
		anIndex: Integer from Standard;
		X, Y: Length from Quantity;
        aWidth: Length from Quantity;
        anHeight: Length from Quantity;
        anAngle: PlaneAngle from Quantity = 0.0)
	---Level: Public
	---Purpose: Add a marker of predefined index <anIndex> in the set 
        --          at position <X>,<Y> and size <aWidth>,<aHeight>.
        --          Angle is measured counterclockwise with 0 radian
        --          at 3 o'clock.
        --  Trigger: Raises MarkerDefinitionError if the
        --          marker index is <= 0 or undefined in the MarkMap,
        --          or the marker size <aWidth,anHeight> is <= 0.
	raises MarkerDefinitionError from Graphic2d;
	---Category: Update method

	Length(me) returns Integer from Standard;
	---Level: Public
	---Purpose: Returns the number of markers in the set.
	---Category: Inquiry method

	Values( me; 
            aRank   :     Integer    from Standard;
            anIndex : out Integer    from Standard;
            X, Y    : out Length     from Quantity;
            aW, aH  : out Length     from Quantity;
            anAngle : out PlaneAngle from Quantity )
	---Level: Public
	---Purpose: Returns the marker type, position, sizes and angle 
    	--          and type from the set at rank <aRank>.
	--  Warning: For the pixel point marker the returned <anIndex> is NULL 
	--  Trigger: Raises OutOfRange if <aRank> is <1 or >Length()
	raises OutOfRange from Standard;
	---Category: Inquiry method

	--------------------------
	-- Category: Draw and Pick
	--------------------------

	Draw (me : mutable; aDrawer: Drawer from Graphic2d)
	is static protected;
	---Level: Internal
	---Purpose: Draws the set of markers <me>.

	DrawElement( me : mutable; aDrawer: Drawer from Graphic2d;
                 anIndex: Integer from Standard)
        is redefined protected;
    	---Level: Internal
    	---Purpose: Draws element <anIndex> of the set <me>.

    	---SAV
	DrawPickedElements(me : mutable; aDrawer: Drawer from Graphic2d )
	is redefined protected;
	---Level: Internal
	---Purpose: Draws the all picked elements of the primitive <me>.

    	---SAV
    	DrawSelectedElements(me : mutable; aDrawer: Drawer from Graphic2d )
	is redefined protected;
	---Level: Internal
	---Purpose: Draws the all selected elements of the primitive <me>.

    	---SAV
    	SetElementsSelected(me : mutable) returns Boolean from Standard
	is redefined;
	---Level: Public
	---Purpose: Declares that previously highlighted elements will be selected ones.

    	---SAV
    	HasSelectedElements(me : mutable)
	returns Boolean from Standard is redefined;
	---Level: Public

    	---SAV
    	DrawElements(me : mutable; aDrawer  : Drawer from Graphic2d;
    	    	    	    	   x,y      : HArray1OfShortReal from TShort)
	is private;
	---Level: Internal

    	---SAV
    	ClearSelectedElements(me : mutable)
	is redefined;
	---Level: Public

    	---SAV
    	GetSelectedElements(me)
	returns MapOfInteger from TColStd;
	---C++: return const &

    	---SAV
    	AddOrRemoveSelected(me : mutable; index : Integer from Standard);
	---Level: Public
	---Purpose: adds/removes marker to/from selection map.

    DrawVertex( me : mutable; aDrawer: Drawer from Graphic2d;
                anIndex: Integer from Standard)
        is redefined protected;
    	---Level: Internal
    	---Purpose: Draws vertex <anIndex> of the set <me>.

	Pick (me : mutable; X, Y: ShortReal from Standard;
		aPrecision: ShortReal from Standard;
		aDrawer: Drawer from Graphic2d)
	returns Boolean from Standard
	is static protected;
	---Level: Internal
        ---Purpose: Returns Standard_True if one marker of the set <me> 
	--	    is picked, Standard_False if not.
	--  Warning: The PickIndex() method returns the rank of the picked
	--	    marker if any.

	----------------------------------------------------------------------

	Save( me; aFStream: in out FStream from Aspect ) is virtual;
--	Retrieve( me; aIFStream: in out IFStream from AIS2D ) is virtual;

    	---SAV
	Pick (me : mutable; X1, Y1, X2, Y2 : ShortReal from Standard;
		    	    aDrawer        : Drawer from Graphic2d;
    	    	    	    aPickMode      : PickMode from Graphic2d)
	returns Boolean from Standard is redefined protected;

    	---SAV
	PickByCircle(me : mutable; x, y, radius : ShortReal from Standard;
		    	    aDrawer      : Drawer from Graphic2d;
    	    	    	    aPickMode    : PickMode from Graphic2d)
	returns Boolean from Standard is redefined protected;
	
	---SAV
	SetHighlightedLimit(me:mutable; number : Integer from Standard);
	---Level: Public
	---Purpose: sets limit of number elements to be highlighted.

    	---SAV
    	SetScaledWidth( me: mutable; width : ShortReal from Standard );
	---Purpose: Changes myScaledWidth field. As this value used in detection
	--          mechanism it should be reset after view transformation.
	
fields

	myType:	    SequenceOfInteger from TColStd;
	myX:	    SequenceOfShortReal from TShort;
	myY:	    SequenceOfShortReal from TShort;
	myWidth:	SequenceOfShortReal from TShort;
	myHeight:	SequenceOfShortReal from TShort;
	myAngle:	SequenceOfShortReal from TShort;
    	mySelIndices    : HSequenceOfInteger from TColStd;
	myMapOfSelected : MapOfInteger from TColStd;
	myHLimit        : Integer from Standard;
	mySuppressHigh  : Boolean from Standard;
	myScaledWidth   : Length from Quantity;

end SetOfMarkers from Graphic2d;
