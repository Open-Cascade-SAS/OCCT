-- Created on: 1996-02-28
-- Created by: Philippe MANGIN
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class MultipleVarFunctionWithHessian from math 
      inherits MultipleVarFunctionWithGradient  from math

	---Purpose: 

uses Matrix from math,
     Vector from math

is
    NbVariables(me)
    	---Purpose: returns the number of variables of the function.

    returns Integer is deferred;


    Value(me: in out; X: Vector; F: out Real)
    	---Purpose: computes the values of the Functions <F> for the 
    	--          variable <X>.
    	--          Returns True if the computation was done successfully, 
    	--          False otherwise.

    returns Boolean is deferred;
    
    
    Gradient(me: in out; X: Vector; G: out Vector)
    	---Purpose:computes the gradient <G> of the functions for the 
    	--         variable <X>.
    	--         Returns True if the computation was done successfully, 
    	--         False otherwise.

    returns Boolean is deferred;
    
    
    Values(me: in out; X: Vector; F: out Real; G: out Vector)
    	---Purpose: computes the value <F> and the gradient <G> of the 
    	--          functions for the variable <X>.
    	--          Returns True if the computation was done successfully, 
    	--          False otherwise.

    returns Boolean is deferred;
    
    Values(me: in out; X: Vector; F: out Real; G: out Vector; H: out Matrix)
    	---Purpose: computes the value  <F>, the gradient <G> and  the
    	--          hessian   <H> of  the functions  for the  variable <X>.
    	--          Returns  True  if  the computation  was  done
    	--          successfully, False otherwise.

    returns Boolean is deferred;

end MultipleVarFunctionWithHessian;
