-- Created on: 1991-10-28
-- Created by: Remi LEQUETTE
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package TopTrans 

	---Purpose: This   package provides  algorithms  to    compute
	--          complex transitions. A transition is the status of
	--          geometry near the boundary of a Shape.  An example
	--          is  the  intersection of  a  curve  and  a surface
	--          enclosing a solid   , the transition  tells if the
	--          parts of the curve just  before and just after the
	--          intersection  are   inside, outside   or   on  the
	--          boundary of the solid.
	--          
	--          The difficulty with transitions arise when dealing
	--          with trimmed geometries like edges and faces. When
	--          the geometric intersections are inside the trimmed
	--          geometry the transition is usually computed by the
	--          intersection algorithms   as the  trimming can  be
	--          safely ignored. If the  intersection  falls on the
	--          trimming  boundaries   one  must   consider    the
	--          neighbouring entities. Consider as  an example the
	--          intersection  of a  curve   and a   solid,  if the
	--          intersection falls on an edge of the solid it does
	--          not falls inside  the  two faces  adjacent to  the
	--          edge, a complex transition occurs.
	--          
	--          This package provides two classes :
	--          
	--              * CurveTransition is  used to compute  complex
	--              transitions with an other curve.
	--              
	--              * SurfaceTransition is used to compute complex
	--              transitions in 3D space.
	--              
        --         The curves and surfaces are  given   by a first  or
        --         second order  approximation around the intersection
        --         point.   For a  curve, the  tangent  vector or  the
        --         osculating circle. For  a surface the normal vector
        --         or the osculating quadric.

uses
    Standard,
    TCollection,
    TColStd,
    gp,
    TopAbs

is
    
    class Array2OfOrientation instantiates 
    	Array2 from TCollection (Orientation from TopAbs);
    
    class CurveTransition;
    
    class SurfaceTransition;

end TopTrans;
