-- Created on: 1995-01-23
-- Created by: Mister rmi
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package SelectBasics 

	---Purpose:  kernel of dynamic selection:
	--           - contains the algorithm to sort the sensitive areas
	--           before the selection action;->quick selection of
	--           an item in a set of items...
	--           - contains the entities able to give the algorithm
	--             sensitive areas .

uses
    Bnd,
    TCollection,
    TColStd,
    Standard,
    MMgt,
    gp,
    TColgp,
    TopLoc
    

is


    deferred class EntityOwner;
    ---Purpose: entity able to set multiple owners for a SensitiveEntity;

    class SortAlgo; 
    ---Purpose: sort algorithm for 2D rectangles.

    class BasicTool;
    ---Purpose: give Tools for sorting Selection results
    --          (example : sensitive entities matching)

    class ListOfBox2d instantiates List from TCollection 
    (Box2d from Bnd);
    

    class SequenceOfOwner instantiates Sequence from TCollection 
    (EntityOwner);
    


    deferred class SensitiveEntity;
    ---Purpose: general entity able to give sensitive areas 


    class ListOfSensitive instantiates List from TCollection 
    (SensitiveEntity);

    imported PickArgs;
    ---Purpose: Structure to provide all-in-one information on picking arguments
    -- for "Matches" method of SelectBasics_SensitiveEntity.

    MaxOwnerPriority returns Integer;
    
    MinOwnerPriority returns Integer;


end SelectBasics;
