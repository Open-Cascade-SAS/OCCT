-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package StepGeom 

    ---Purpose : AP214 CC1 , Revision 4  for Geom (Part42, geometric)
    --           Upgrading from Revision 2 to Revision 4 : 26 Mar 1997

uses


	TCollection, TColStd, StepData, Interface, MMgt,
	StepBasic, StepRepr

is


enumeration BSplineCurveForm is     -- reordered from Rev2 to Rev4

	bscfPolylineForm,
	bscfCircularArc,
	bscfEllipticArc,
	bscfParabolicArc,
	bscfHyperbolicArc,
	bscfUnspecified
end;

enumeration BSplineSurfaceForm is   -- reordered from Rev2 to Rev4

	bssfPlaneSurf,
	bssfCylindricalSurf,
	bssfConicalSurf,
	bssfSphericalSurf,
	bssfToroidalSurf,
	bssfSurfOfRevolution,
	bssfRuledSurf,
	bssfGeneralisedCone,
	bssfQuadricSurf,
	bssfSurfOfLinearExtrusion,
	bssfUnspecified
end;

enumeration KnotType is     -- reordered from Rev2 to Rev4

	ktUniformKnots,
	ktUnspecified,
	ktQuasiUniformKnots,
	ktPiecewiseBezierKnots
end;

enumeration PreferredSurfaceCurveRepresentation is   -- reordered Rev2 to Rev4

	pscrCurve3d,
	pscrPcurveS1,
	pscrPcurveS2
end;

-- Removed from Rev2 to Rev4 :enumeration TextPath

enumeration TransitionCode is   -- reordered from Rev2 to Rev4

	tcDiscontinuous,
	tcContinuous,
	tcContSameGradient,
	tcContSameGradientSameCurvature
end;

enumeration TrimmingPreference is   -- reordered from Rev2 to Rev4

	tpCartesian,
	tpParameter,
	tpUnspecified
end;

class Axis2Placement;		-- Select Type for

	-- Axis2Placement2d
	-- Axis2Placement3d


class CurveOnSurface;		-- Select Type for

	-- Pcurve
	-- SurfaceCurve
	-- CompositeCurveOnSurface

class PcurveOrSurface;		-- Select Type for

	-- Pcurve
	-- Surface


class TrimmingSelect;		-- Select Type for

	-- CartesianPoint
	-- ParameterValue i.e. Real (TrimmingMember)

class TrimmingMember;

class VectorOrDirection;		-- Select Type for

	-- Vector
	-- Direction


--class Protocol;


class CompositeCurveSegment;
	class ReparametrisedCompositeCurveSegment;
--class RepresentationContext;
	class GeometricRepresentationContext;
	class GeometricRepresentationContextAndGlobalUnitAssignedContext;
    	-- Hand Made by FMA :
	class GeomRepContextAndGlobUnitAssCtxAndGlobUncertaintyAssCtx;     
    	-- Hand Made by FMA :
	class GeometricRepresentationContextAndParametricRepresentationContext;
--class RepresentationItem;
	class GeometricRepresentationItem;
		class CartesianTransformationOperator;
			class CartesianTransformationOperator2d;
			class CartesianTransformationOperator3d;
		class Curve;
			class BoundedCurve;
				class BSplineCurve;
					class BSplineCurveWithKnots;
					class BezierCurve;
					class QuasiUniformCurve;
					class RationalBSplineCurve;
					class UniformCurve;
					class UniformCurveAndRationalBSplineCurve;
					class BSplineCurveWithKnotsAndRationalBSplineCurve;
					class QuasiUniformCurveAndRationalBSplineCurve;
					class BezierCurveAndRationalBSplineCurve;
				class CompositeCurve;
					class CompositeCurveOnSurface;
						class BoundaryCurve;
							class OuterBoundaryCurve;
				class Polyline;
				class TrimmedCurve;
			class Conic;
				class Circle;
				class Ellipse;
				class Hyperbola;
				class Parabola;
			class CurveReplica;
			class Line;
			class OffsetCurve3d;
			class Pcurve;
			class SurfaceCurve;
				class IntersectionCurve;
				class SeamCurve;
			    class SurfaceCurveAndBoundedCurve;
		class Direction;
		class Placement;
			class Axis1Placement;
			class Axis2Placement2d;
			class Axis2Placement3d;
--V		class PlanarExtent;
--V			class PlanarBox;
		class Point;
			class CartesianPoint;
			class DegeneratePcurve;
				class EvaluatedDegeneratePcurve;
			class PointOnCurve;
			class PointOnSurface;
			class PointReplica;
		class Surface;
			class BoundedSurface;
				class BSplineSurface;
					class BSplineSurfaceWithKnots;
					class BezierSurface;
					class QuasiUniformSurface;
					class RationalBSplineSurface;
					class UniformSurface;
					class BSplineSurfaceWithKnotsAndRationalBSplineSurface;
					class UniformSurfaceAndRationalBSplineSurface;
					class QuasiUniformSurfaceAndRationalBSplineSurface;
					class BezierSurfaceAndRationalBSplineSurface;
				class CurveBoundedSurface;
				class RectangularCompositeSurface;
				class RectangularTrimmedSurface;
			class ElementarySurface;
				class ConicalSurface;
				class CylindricalSurface;
				class Plane;
				class SphericalSurface;
				class ToroidalSurface;
					class DegenerateToroidalSurface;
			class OffsetSurface;
			class SurfaceReplica;
			class SweptSurface;
				class SurfaceOfLinearExtrusion;
				class SurfaceOfRevolution;
			class OrientedSurface; --  Added from AP214 DIS to IS 4.01.2002
		class Vector;
class SurfacePatch;
class SurfaceBoundary;


imported Array1OfCurve;
imported transient class HArray1OfCurve;

imported Array1OfCartesianPoint;
imported transient class HArray1OfCartesianPoint;

imported Array2OfCartesianPoint;
imported transient class HArray2OfCartesianPoint;

imported Array1OfCompositeCurveSegment;
imported transient class HArray1OfCompositeCurveSegment;

imported Array1OfBoundaryCurve;
imported transient class HArray1OfBoundaryCurve;

imported Array2OfSurfacePatch;
imported transient class HArray2OfSurfacePatch;

imported Array1OfSurfaceBoundary;
imported transient class HArray1OfSurfaceBoundary;

imported Array1OfPcurveOrSurface;
imported transient class HArray1OfPcurveOrSurface;

imported Array1OfTrimmingSelect;
imported transient class HArray1OfTrimmingSelect;

--	Protocol returns Protocol from StepGeom;

end StepGeom;

