-- Created on: 1996-12-16
-- Created by: Christian CAILLET
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SelectNamed  from StepData    inherits SelectMember

    ---Purpose : This select member can be of any kind, and be named
    --           But its takes more memory than some specialised ones
    --           This class allows one name for the instance

uses CString, Logical, AsciiString from TCollection,  Field from StepData

is

    Create  returns mutable SelectNamed;

    HasName (me) returns Boolean  is redefined;

    Name (me) returns CString  is redefined;

    SetName (me : mutable; name : CString)  returns Boolean  is redefined;
    -- redefined to accept any name

    Field (me) returns Field;
    ---C++ : return const &

    CField (me : mutable) returns Field;
    ---C++ : return &


    Kind (me) returns Integer  is redefined;
    --  see Field for Kind (same codes)

    SetKind  (me : mutable; kind : Integer)  is redefined;
    --  called by various Set*

    Int (me) returns Integer  is redefined;
    ---Purpose : This internal method gives access to a value implemented by an
    --           Integer (to read it)

    SetInt (me : mutable; val : Integer)  is redefined;
    ---Purpose : This internal method gives access to a value implemented by an
    --           Integer (to set it)

    Real (me) returns Real  is redefined;

    SetReal (me : mutable; val : Real)  is redefined;

    String (me) returns CString  is redefined;

    SetString (me : mutable; val : CString)  is redefined;

fields

    thename : AsciiString;
    theval  : Field from StepData;

end SelectNamed;
