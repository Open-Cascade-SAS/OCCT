-- Created on: 1997-12-08
-- Created by: Serguei ZARITCHNY
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class FilletRadiusPresentation from DsgPrs

        ---Purpose: A framework for displaying radii of fillets.
uses
    Presentation from Prs3d,
    Pnt from gp,
    Dir from gp,
    Drawer from Prs3d,
    ExtendedString from TCollection,
    ArrowSide from DsgPrs,
    TrimmedCurve from Geom,
    Circle  from Geom,
    Ax1 from gp
is
    Add( myclass; aPresentation : Presentation from Prs3d;
    	    	  aDrawer       : Drawer from Prs3d;
		  thevalue      : Real from Standard;
		  aText         : ExtendedString from TCollection;
		  aPosition     : Pnt from gp;
		  aNormalDir    : Dir from gp;
		  aBasePnt      : Pnt from gp;
		  aFirstPoint   : Pnt from gp;
		  aSecondPoint  : Pnt from gp;
		  aCenter       : Pnt from gp;
		  ArrowPrs      : ArrowSide from DsgPrs; 
		  drawRevers    : Boolean from Standard; 
    	    	  DrawPosition  : out Pnt from gp;
    	    	  EndOfArrow    : out Pnt from gp;
    	    	  TrimCurve     : out TrimmedCurve from Geom;
    	    	  HasCircle     : out Boolean from Standard);
    	---Purpose: Adds a display of the radius of a fillet to the
    	-- presentation aPresentation. The display ttributes
    	-- defined by the attribute manager aDrawer. the value
    	-- specifies the length of the radius.
		  
end FilletRadiusPresentation;
