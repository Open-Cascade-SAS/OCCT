-- Created on: 1991-11-21
-- Created by: NW,JPB,CAL
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PickDescriptor from Visual3d

	---Version:

	---Purpose: This class contains the pick information.
	--	    It contains a certain number of PickPaths.

	---Keywords: Pick Descriptor, Path, Structure, PickId

	---Warning:
	---References:

uses

	Structure		from Graphic3d,
	ContextPick		from Visual3d,
	PickPath		from Visual3d,
	HSequenceOfPickPath	from Visual3d

raises

	PickError		from Visual3d

is

	Create ( CTX : ContextPick from Visual3d )
		returns PickDescriptor from Visual3d;
	---Level: Public
	---Purpose: Creates a PickDescriptor <me>.

	---------------------------------------------------
	-- Category: Methods to modify the class definition
	---------------------------------------------------

	AddPickPath ( me	: in out;
		      APickPath	: PickPath from Visual3d )
		is static;
	---Level: Public
	---Purpose: Adds a PickPath to PickDescriptor <me>.
	---Category: Methods to modify the class definition

	Clear ( me : in out )
		is static;
	---Level: Public
	---Purpose: Erases all the information in <me>.
	---Category: Methods to modify the class definition

	----------------------------
	-- Category: Inquire methods
	----------------------------

	Depth ( me )
		returns Integer from Standard
		is static;
	---Level: Public
	---Purpose: Returns the pick depth, that is the
	--	    number of PickPaths available in the PickDescriptor.
	---Category: Inquire methods

	PickPath ( me )
		returns HSequenceOfPickPath from Visual3d
		is static;
	---Level: Internal
	---Purpose: Returns the group of PickPaths of <me>.
	---Category: Inquire methods

	TopStructure ( me )
		returns Structure from Graphic3d
	---Level: Public
	---Purpose: Returns the root structure.
	--	    If the pick order was of the type TOO_TOPFIRST
	--	    then it's the first structure.
	--	    If the pick order was of the type TOO_BOTTOMFIRST
	--	    Then it's the last structure.
	--	    The pick order is set by the method SetOrder
	--	    from ContextPick.
	--  Category: Inquire methods
	--  Warning: Raises PickError if Depth == 0 (no picked structure).
	raises PickError from Visual3d is static;

	TopPickId ( me )
		returns Integer from Standard
	---Level: Public
	---Purpose: Returns the root structure pickid.
	--	    If the pick order was of the type TOO_TOPFIRST
	--	    then it's the first pickid.
	--	    If the pick order was of the type TOO_BOTTOMFIRST
	--	    then it's the last pickid.
	--	    The pick order is set by the method SetOrder
	--	    from ContextPick.
	--  Category: Inquire methods
	--  Warning: Raises PickError if Depth == 0 (no picked structure).
	raises PickError from Visual3d is static;

	TopElementNumber ( me )
		returns Integer from Standard
	---Level: Public
	---Purpose: Returns the root structure element number.
	--	    If the pick order was of the type TOO_TOPFIRST
	--	    then it's the first element number.
	--	    If the pick order was of the type TOO_BOTTOMFIRST
	--	    then it's the last element number.
	--	    The pick order is set by the method SetOrder
	--	    from ContextPick.
	--  Category: Inquire methods
	--  Warning: Raises PickError if Depth == 0 (no picked structure).
	raises PickError from Visual3d is static;

--

fields

--
-- Class	:	Visual3d_PickDescriptor
--
-- Purpose	:	Declaration of variables specific to the class
--			describing a pick.
--
-- Reminders 	: 	A pick return is defined by:
--			- a sequence of (Elem_number, Pick_Id, Struct_Id)
--			- a depth

	-- pick sequence
	MyPickPathSequence	:	HSequenceOfPickPath from Visual3d;

	-- context associated to a pick
	MyContext		:	ContextPick from Visual3d;

end PickDescriptor;
