-- Created on: 1993-07-12
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class MakeFace from BRepLib inherits MakeShape from BRepLib 

	---Purpose: Provides methods to build faces.
	--          
	--          A face may be built :
	--          
	--          * From a surface.
	--          
	--             - Elementary surface from gp.
	--             
	--             - Surface from Geom.
	--             
	--          * From a surface and U,V values.
	--          
	--          * From a wire.
	--            
	--            - Find the surface automatically if possible.
	--          
	--          * From a surface and a wire.
	--          
	--            - A flag Inside is given, when this flag is True
	--            the  wire is  oriented to bound a finite area on
	--            the surface.
	--          
	--          * From a face and a wire.
	--            
	--            - The new wire is a perforation.

uses
    Pln       from gp,
    Cylinder  from gp,
    Cone      from gp,
    Sphere    from gp,
    Torus     from gp,
    Surface   from Geom,
    Face      from TopoDS,
    Wire      from TopoDS,
    FaceError from BRepLib
    
raises
    NotDone    from StdFail

is

    Create  
	---Purpose: Not done.
	---Level: Public
    returns MakeFace from BRepLib;
    
    Create(F : Face from TopoDS)  
	---Purpose: Load a face. Usefull to add wires.
	---Level: Public
    returns MakeFace from BRepLib;

    ----------------------------------------------
    -- From a surface
    ----------------------------------------------

    Create(P : Pln from gp)
	---Purpose: Make a face from a plane.
	---Level: Public
    returns MakeFace from BRepLib;

    Create(C : Cylinder from gp)
	---Purpose: Make a face from a cylinder.
	---Level: Public
    returns MakeFace from BRepLib;

    Create(C : Cone from gp)
	---Purpose: Make a face from a cone.
	---Level: Public
    returns MakeFace from BRepLib;

    Create(S : Sphere from gp)
	---Purpose: Make a face from a sphere.
	---Level: Public
    returns MakeFace from BRepLib;

    Create(C : Torus from gp)
	---Purpose: Make a face from a torus.
	---Level: Public
    returns MakeFace from BRepLib;

    Create(S : Surface from Geom; TolDegen : Real)
    ---Purpose: Make a face from a Surface. Accepts tolerance value (TolDegen)
    --          for resolution of degenerated edges.
    ---Level: Public
    returns MakeFace from BRepLib;

    ----------------------------------------------
    -- From a surface and U,V values
    ----------------------------------------------

    Create(P : Pln from gp; UMin, UMax, VMin, VMax : Real)
	---Purpose: Make a face from a plane.
	---Level: Public
    returns MakeFace from BRepLib;

    Create(C : Cylinder from gp; UMin, UMax, VMin, VMax : Real)
	---Purpose: Make a face from a cylinder.
	---Level: Public
    returns MakeFace from BRepLib;

    Create(C : Cone from gp; UMin, UMax, VMin, VMax : Real)
	---Purpose: Make a face from a cone.
	---Level: Public
    returns MakeFace from BRepLib;

    Create(S : Sphere from gp; UMin, UMax, VMin, VMax : Real)
	---Purpose: Make a face from a sphere.
	---Level: Public
    returns MakeFace from BRepLib;

    Create(C : Torus from gp; UMin, UMax, VMin, VMax : Real)
	---Purpose: Make a face from a torus.
	---Level: Public
    returns MakeFace from BRepLib;

    Create(S : Surface from Geom; UMin, UMax, VMin, VMax, TolDegen : Real)
    ---Purpose: Make a face from a Surface. Accepts min & max parameters
    --          to construct the face's bounds. Also accepts tolerance value (TolDegen)
    --          for resolution of degenerated edges.
    ---Level: Public
    returns MakeFace from BRepLib;

    ----------------------------------------------
    -- From a wire
    ----------------------------------------------

    Create(W         : Wire    from TopoDS;
    	   OnlyPlane : Boolean from Standard = Standard_False)
	---Purpose: Find a surface from the wire and make a face.
	--          if <OnlyPlane> is true, the computed surface will be
	--          a plane. If it is not possible to find a plane, the
	--          flag NotDone will be set.
	---Level: Public
    returns MakeFace from BRepLib;

    ----------------------------------------------
    -- From a surface and a wire
    ----------------------------------------------

    Create(P : Pln from gp; W : Wire from TopoDS;
    	   Inside : Boolean = Standard_True)
	---Purpose: Make a face from a plane and a wire.
	---Level: Public
    returns MakeFace from BRepLib;

    Create(C : Cylinder from gp; W : Wire from TopoDS;
    	   Inside : Boolean = Standard_True)
	---Purpose: Make a face from a cylinder and a wire.
	---Level: Public
    returns MakeFace from BRepLib;

    Create(C : Cone from gp; W : Wire from TopoDS;
    	   Inside : Boolean = Standard_True)
	---Purpose: Make a face from a cone and a wire.
	---Level: Public
    returns MakeFace from BRepLib;

    Create(S : Sphere from gp; W : Wire from TopoDS;
    	   Inside : Boolean = Standard_True)
	---Purpose: Make a face from a sphere and a wire.
	---Level: Public
    returns MakeFace from BRepLib;

    Create(C : Torus from gp; W : Wire from TopoDS;
    	   Inside : Boolean = Standard_True)
	---Purpose: Make a face from a torus and a wire.
	---Level: Public
    returns MakeFace from BRepLib;

    Create(S : Surface from Geom; W : Wire from TopoDS;
    	   Inside : Boolean = Standard_True)
	---Purpose: Make a face from a Surface and a wire.
	---Level: Public
    returns MakeFace from BRepLib;

    ----------------------------------------------
    -- From face and wire.
    ----------------------------------------------

    Create(F : Face from TopoDS; W : Wire from TopoDS)
	---Purpose: Adds the wire <W> in the face <F>
	---Level: Public
    returns MakeFace from BRepLib;
    
    ----------------------------------------------
    -- Auxiliary methods
    ----------------------------------------------

    Init(me : in out; F : Face from TopoDS)
	---Purpose: Load the face.
	---Level: Public
    is static;

    Init(me : in out; S : Surface from Geom; Bound : Boolean; TolDegen : Real)
    ---Purpose: Creates the face  from the  surface. If Bound is
    --          True a wire is made from the natural bounds.
    --          Accepts tolerance value (TolDegen) for resolution
    --          of degenerated edges.
    ---Level: Public
    is static;

    Init(me : in out; S : Surface from Geom; UMin, UMax, VMin, VMax, TolDegen : Real) 
    ---Purpose: Creates the face from the surface and the min-max
    --          values. Accepts tolerance value (TolDegen) for resolution
    --          of degenerated edges.
    ---Level: Public
    is static;

    Add(me : in out; W : Wire from TopoDS)
	---Purpose: Adds the wire <W> in the current face.
	---Level: Public
    is static;

    ----------------------------------------------
    -- Auxiliary methods
    ----------------------------------------------

    CheckInside(me : in out)
	---Purpose: Reorient the current face if  the boundary  is not
	--          finite.
	---Level: Public
    is static private;

    ----------------------------------------------
    -- Results
    ----------------------------------------------

    Error(me) returns FaceError from BRepLib
	---Level: Public
    is static;

    Face(me) returns Face from TopoDS
	---Purpose: Returns the new face.
	--          
	---C++: return const &
	---C++: alias "Standard_EXPORT operator TopoDS_Face() const;"
	---Level: Public
    raises 
    	NotDone from StdFail
    is static;
    
fields
    myError    : FaceError from BRepLib;
end MakeFace;
