-- Created on: 1997-12-09
-- Created by: Jean-Louis Frenkel
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


private class ReadWriter_1 from PCDM inherits ReadWriter from PCDM

uses
    ExtendedString from TCollection,  
    AsciiString from TCollection, 
    Data from Storage, 
    Document from CDM, 
    MessageDriver from CDM, 
    SequenceOfExtendedString from TColStd, 
    SequenceOfReference from PCDM

is

    Create returns mutable ReadWriter_1 from PCDM;
   
    Version(me) returns AsciiString from TCollection;
    ---Purpose: returns PCDM_ReadWriter_1.
   
    WriteReferenceCounter(me; aData: mutable Data from Storage; aDocument: Document from CDM);

    WriteReferences(me; aData: mutable Data from Storage; aDocument: Document from CDM; theReferencerFileName: ExtendedString from TCollection);

    
    WriteExtensions(me; aData: mutable Data from Storage; aDocument: Document from CDM);

    
    WriteVersion(me; aData: mutable Data from Storage; aDocument: Document from CDM);

    
    ReadReferenceCounter(me; aFileName: ExtendedString from TCollection; theMsgDriver: MessageDriver from CDM)
    returns Integer from Standard;

    ReadReferences(me; aFileName: ExtendedString from TCollection; theReferences: in out  SequenceOfReference from PCDM; theMsgDriver: MessageDriver from CDM);

    
    ReadExtensions(me; aFileName: ExtendedString from TCollection; theExtensions: in out  SequenceOfExtendedString from TColStd; theMsgDriver: MessageDriver from CDM);

    ReadUserInfo(myclass; aFileName: ExtendedString from TCollection; Start, End: AsciiString from TCollection; theUserInfo:in  out SequenceOfExtendedString from TColStd;theMsgDriver: MessageDriver from CDM)
    is private;

    ReadDocumentVersion(me; aFileName: ExtendedString from TCollection; theMsgDriver: MessageDriver from CDM)
    returns Integer from Standard;


end ReadWriter_1 from PCDM;
