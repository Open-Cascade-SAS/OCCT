-- Created on: 1992-10-08
-- Created by: Isabelle GRIGNON
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



package GeomAdaptor 

	---Purpose: this package contains the  geometric definition of
	--          curve and surface necessary to use algorithmes.

uses 
    Geom,
    GeomAbs,
    Adaptor3d,
    gp,
    Standard,
    TColStd,
    Geom2dAdaptor,
    TColgp,
    Precision

is
      class Curve; 
        ---Purpose: creation of the loaded curve the curve is C1 by piece.
        --          Inherits  Curve from Adaptor3d 

      class Surface;
        ---Purpose: creation of the loaded surface the surface is C1 by piece 
        --          Inherits  Surface from Adaptor3d 

      private class GHSurface instantiates GenHSurface from Adaptor3d
      	    (Surface from GeomAdaptor);
	    
      class HSurface;
	---Purpose: Inherited  from    GHSurface.   Provides a  surface
	--          handled by reference.

      private class GHCurve instantiates GenHCurve from Adaptor3d
            (Curve from GeomAdaptor);
      
      class HCurve;
	---Purpose: Inherited  from    GHCurve.   Provides a  curve
	--          handled by reference.

    
      MakeCurve( C : Curve from Adaptor3d)
	---Purpose: Build a Geom_Curve using the informations from the 
	--          Curve from Adaptor3d
      returns Curve from Geom;
      
      MakeSurface( S : Surface from Adaptor3d)
	---Purpose: Build a Geom_Surface using the informations from the 
	--          Surface from Adaptor3d
      returns Surface from Geom;
      
end GeomAdaptor;
