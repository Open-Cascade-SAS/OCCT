-- Created on: 1993-06-03
-- Created by: Bruno DUMORTIER
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Curve from Geom2dAdaptor inherits Curve2d from Adaptor2d

        ---Purpose: An interface between the services provided by any
    	-- curve from the package Geom2d and those required
    	-- of the curve by algorithms which use it.
        
uses Vec2d                  from gp,
     Pnt2d                  from gp,
     Circ2d                 from gp,
     Elips2d                from gp,
     Hypr2d                 from gp,
     Parab2d                from gp,
     Lin2d                  from gp,
     Array1OfReal           from TColStd,
     Curve                  from Geom2d,
     BezierCurve            from Geom2d,
     BSplineCurve           from Geom2d,
     CurveType              from GeomAbs,
     Shape                  from GeomAbs,
     HCurve2d               from Adaptor2d,
     Cache                  from BSplCLib
     
     
raises NoSuchObject from Standard,
       ConstructionError from Standard,
       OutOfRange  from Standard,
       DomainError from Standard


is

    Create returns Curve from Geom2dAdaptor;

    Create(C : Curve from Geom2d) returns Curve from Geom2dAdaptor;

    Create(C : Curve from Geom2d; UFirst,ULast : Real)
    returns Curve from Geom2dAdaptor
    raises 
    	ConstructionError from Standard;
    	---Purpose: ConstructionError is raised if Ufirst>Ulast
   
    Load(me : in out; C : Curve from Geom2d);
    	---C++: inline
   
    Load(me : in out; C : Curve from Geom2d; UFirst,ULast : Real)
    raises 
    	ConstructionError from Standard;
    	---C++: inline
    	---Purpose: ConstructionError is raised if Ufirst>Ulast

    Curve(me) returns Curve from Geom2d
        ---C++: return const& 
    	---C++: inline
    is static;



    FirstParameter(me) returns Real
	---C++: inline
    is redefined static;

    LastParameter(me) returns Real
	---C++: inline
    is redefined static;     

    Continuity(me) returns Shape from GeomAbs
    is redefined static;

    NbIntervals(me; S : Shape from GeomAbs) returns Integer
	---Purpose: If necessary,  breaks the  curve in  intervals  of
	--          continuity  <S>.    And  returns   the number   of
	--          intervals.
    is redefined static;

    Intervals(me; T : in out Array1OfReal from TColStd; 
    	          S : Shape from GeomAbs)
	---Purpose: Stores in <T> the  parameters bounding the intervals
	--          of continuity <S>.
	--          
	--          The array must provide  enough room to  accomodate
	--          for the parameters. i.e. T.Length() > NbIntervals()
    raises
    	OutOfRange from Standard 
    is redefined static;
    
    Trim(me; First, Last, Tol : Real) returns HCurve2d from Adaptor2d
	---Purpose: Returns    a  curve equivalent   of  <me>  between
	--          parameters <First>  and <Last>. <Tol>  is used  to
	--          test for 3d points confusion.
    raises
    	OutOfRange from Standard
	---Purpose: If <First> >= <Last> 
    is redefined static;
    
    IsClosed(me) returns Boolean
    is redefined static;
    
    IsPeriodic(me) returns Boolean
    is redefined static;

    Period(me) returns Real
    raises
    	DomainError from Standard -- if the curve is not periodic
    is redefined static;

    
    Value(me; U : Real) returns Pnt2d from gp
        --- Purpose : Computes the point of parameter U on the curve 
    is redefined static;

    ValueBSpline(me; U: Real) returns Pnt2d from gp
        --- Purpose : Computes the point of parameter U on the B-spline curve
    is private;

    ValueOffset(me; U: Real) returns Pnt2d from gp
        --- Purpose : Computes the point of parameter U on the offset curve
    is private;

    D0 (me; U : Real; P : out Pnt2d from gp)
        --- Purpose : Computes the point of parameter U.
    is redefined static;

    D0BSpline(me; theU : Real; theP : out Pnt2d from gp)
        --- Purpose : Computes the point of parameter U on the B-spline curve
    is private;

    D0Offset(me; theU : Real; theP : out Pnt2d from gp)
        --- Purpose : Computes the point of parameter U on the offset curve
    is private;

    D1 (me; U : Real; P : out Pnt2d from gp ; V : out Vec2d from gp)
        --- Purpose : Computes the point of parameter U on the curve with its
        --  first derivative.
    raises 
       DomainError from Standard
        --- Purpose : Raised if the continuity of the current interval
        --  is not C1.
    is redefined static;

    D1BSpline(me; theU : Real; theP : out Pnt2d from gp ; theV : out Vec2d from gp)
        --- Purpose : Computes the point of parameter U on the B-spline curve
        --  and its derivative
    is private;

    D1Offset(me; theU : Real; theP : out Pnt2d from gp ; theV : out Vec2d from gp)
        --- Purpose : Computes the point of parameter U on the offset curve
        --  and its derivative
    is private;
    
    D2 (me; U : Real; P : out Pnt2d from gp; V1, V2 : out Vec2d from gp)
        --- Purpose :
        --  Returns the point P of parameter U, the first and second
        --  derivatives V1 and V2.
    raises 
       DomainError from Standard
        --- Purpose : Raised if the continuity of the current interval
        --  is not C2.
    is redefined static;

    D2BSpline(me; theU : Real; theP : out Pnt2d from gp; theV1, theV2 : out Vec2d from gp)
        --- Purpose : Computes the point of parameter U on the B-spline curve
        --  and its first and second derivatives
    is private;

    D2Offset(me; theU : Real; theP : out Pnt2d from gp; theV1, theV2 : out Vec2d from gp)
        --- Purpose : Computes the point of parameter U on the offset curve
        --  and its first and second derivatives
    is private;

    D3 (me; U : Real; P : out Pnt2d from gp; V1, V2, V3 : out Vec2d from gp)
        --- Purpose :
        --  Returns the point P of parameter U, the first, the second 
        --  and the third derivative.
    raises 
    	DomainError from Standard
        --- Purpose : Raised if the continuity of the current interval
        --  is not C3.
    is redefined static;

    D3BSpline(me; theU : Real; theP : out Pnt2d from gp; theV1, theV2, theV3 : out Vec2d from gp)
        --- Purpose : Computes the point of parameter U on the B-spline curve
        --  and its first, second and third derivatives
    is private;

    D3Offset(me; theU : Real; theP : out Pnt2d from gp; theV1, theV2, theV3 : out Vec2d from gp)
        --- Purpose : Computes the point of parameter U on the offset curve
        --  and its first, second and third derivatives
    is private;
        
    DN (me; U : Real; N : Integer)   returns Vec2d from gp
        --- Purpose :
        --  The returned vector gives the value of the derivative for the 
        --  order of derivation N.
    raises  
    	DomainError from Standard,
        --- Purpose : Raised if the continuity of the current interval
        --  is not CN.
        OutOfRange from Standard
        --- Purpose : Raised if N < 1.            
    is redefined static;

    DNBSpline(me; theU : Real; N : Integer) returns Vec2d from gp
        --- Purpose :
        --  The returned vector gives the value of the derivative for the 
        --  order of derivation N.
    is private;

    DNOffset(me; theU : Real; N : Integer) returns Vec2d from gp
        --- Purpose :
        --  The returned vector gives the value of the derivative for the 
        --  order of derivation N.
    is private;


    Resolution(me; Ruv :Real) returns Real
        ---Purpose : returns the parametric resolution
    is redefined static;   
   

    GetType(me) returns CurveType from GeomAbs
    	---C++: inline
    is redefined static;

    Line(me) returns Lin2d from gp
    raises 
    	NoSuchObject from Standard
    is redefined static;
   
    Circle(me) returns Circ2d from gp
    raises 
    	NoSuchObject from Standard
    is redefined static;

    Ellipse(me) returns Elips2d from gp
    raises 
    	NoSuchObject from Standard
    is redefined static;

    Hyperbola(me) returns  Hypr2d from gp
    raises 
    	NoSuchObject from Standard
    is redefined static;

    Parabola(me) returns Parab2d from gp
    raises 
    	NoSuchObject from Standard
    is redefined static;

     
     Degree(me) returns Integer
     raises 
    	NoSuchObject from Standard
     is redefined static;
     
     IsRational(me) returns Boolean
     raises 
    	NoSuchObject from Standard
     is redefined static;
     
     NbPoles(me) returns Integer
     raises 
    	NoSuchObject from Standard
     is redefined static;

  
     NbKnots(me) returns Integer
     raises 
    	NoSuchObject from Standard
     is redefined static;     
          
    NbSamples(me) returns Integer from Standard is redefined;

    Bezier(me) returns BezierCurve from Geom2d
    raises 
    	NoSuchObject from Standard
    is redefined static;
    
    BSpline(me) returns BSplineCurve from Geom2d
    raises 
    	NoSuchObject from Standard
    is redefined static;
    
    LocalContinuity(me; U1, U2 : Real) returns Shape from GeomAbs 
    is static private;

    load(me : in out; C : Curve from Geom2d; UFirst,ULast : Real)
    is private;
    
    RebuildCache(me; theParameter : Real)
    ---Purpose: Rebuilds B-spline cache
    -- \param theParameter the value on the knot axis which identifies the caching span
    is static private;
   
fields 

  myCurve             : Curve            from Geom2d ;
  myTypeCurve         : CurveType        from GeomAbs ;
  myFirst             : Real             from Standard ;
  myLast              : Real             from Standard;
  myCurveCache        : Cache            from BSplCLib;
  myOffsetBaseCurveAdaptor : HCurve2d    from Adaptor2d;
  
end Curve;

