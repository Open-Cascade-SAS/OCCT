-- Created on: 2002-12-12
-- Created by: data exchange team
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class Volume3dElementDescriptor from StepElement
inherits ElementDescriptor from StepElement

    ---Purpose: Representation of STEP entity Volume3dElementDescriptor

uses
    ElementOrder from StepElement,
    HAsciiString from TCollection,
    HArray1OfVolumeElementPurposeMember from StepElement,
    Volume3dElementShape from StepElement

is
    Create returns Volume3dElementDescriptor from StepElement;
	---Purpose: Empty constructor

    Init (me: mutable; aElementDescriptor_TopologyOrder: ElementOrder from StepElement;
                       aElementDescriptor_Description: HAsciiString from TCollection;
                       aPurpose: HArray1OfVolumeElementPurposeMember from StepElement;
                       aShape: Volume3dElementShape from StepElement);
	---Purpose: Initialize all fields (own and inherited)

    Purpose (me) returns HArray1OfVolumeElementPurposeMember from StepElement;
	---Purpose: Returns field Purpose
    SetPurpose (me: mutable; Purpose: HArray1OfVolumeElementPurposeMember from StepElement);
	---Purpose: Set field Purpose

    Shape (me) returns Volume3dElementShape from StepElement;
	---Purpose: Returns field Shape
    SetShape (me: mutable; Shape: Volume3dElementShape from StepElement);
	---Purpose: Set field Shape

fields
    thePurpose: HArray1OfVolumeElementPurposeMember from StepElement;
    theShape: Volume3dElementShape from StepElement;

end Volume3dElementDescriptor;
