-- Created on: 1993-08-10
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package HLRTopoBRep

	---Purpose: This     Package  provides  some       topological
	--          reconstruction services needed  by the Hidden Line
	--          Removal Algorithms   using OutLine  and    IsoLine
	--          facilities, applied  to an object represented by a
	--          BRep data structure.

uses
    Standard,
    MMgt,
    TCollection,
    TColStd,
    TopoDS,
    TopTools,
    TopExp,
    gp,
    Geom2d,
    IntSurf,
    BRepAdaptor,
    BRepTopAdaptor,
    Contap,
    HLRAlgo
    
is
    class VData;

    class ListOfVData            instantiates List    from TCollection 
    	(VData from HLRTopoBRep);

    class MapOfShapeListOfVData  instantiates DataMap from TCollection
    	(Shape          from TopoDS,
         ListOfVData    from HLRTopoBRep,
         ShapeMapHasher from TopTools);

    class FaceData;

    class DataMapOfShapeFaceData instantiates DataMap from TCollection
    	(Shape          from TopoDS,
	 FaceData       from HLRTopoBRep,
	 ShapeMapHasher from TopTools);
					
    class Data;

    class FaceIsoLiner;
    
    class OutLiner;

    class DSFiller;

end HLRTopoBRep;
