-- Created on: 1998-07-08
-- Created by: Stephanie HUMEAU
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


deferred  class TrihedronWithGuide from GeomFill  
inherits TrihedronLaw from GeomFill

	---Purpose: To define Trihedron along one Curve with a guide
	--          
	--          
	--          
      
uses 
    HCurve from  Adaptor3d, 
    Real  from  Standard 

raises 
    OutOfRange,  NotImplemented   

is  
     
    Guide(me) 
    returns  HCurve  from  Adaptor3d 
    is  deferred;  
     
    Origine(me  :  mutable; 
    	    Param1  :  Real; 
    	    Param2  :  Real) 
    is deferred;
          
fields 
    myGuide  :  HCurve  from  Adaptor3d  is  protected; 
    myTrimG  :  HCurve  from  Adaptor3d  is  protected; 

end TrihedronWithGuide;
    
