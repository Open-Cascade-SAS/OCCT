-- Created on: 2003-06-04
-- Created by: Galina KULIKOVA
-- Copyright (c) 2003-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class ShapeToleranceSelect from StepDimTol
inherits SelectType from StepData

    ---Purpose: Representation of STEP SELECT type ShapeToleranceSelect

uses
    GeometricTolerance from StepDimTol,
    PlusMinusTolerance from StepShape

is
    Create returns ShapeToleranceSelect from StepDimTol;
	---Purpose: Empty constructor

    CaseNum (me; ent: Transient) returns Integer;
	---Purpose: Recognizes a kind of ShapeToleranceSelect select type
	--          1 -> GeometricTolerance from StepDimTol
	--          2 -> PlusMinusTolerance from StepShape
	--          0 else

    GeometricTolerance (me) returns GeometricTolerance from StepDimTol;
	---Purpose: Returns Value as GeometricTolerance (or Null if another type)

    PlusMinusTolerance (me) returns PlusMinusTolerance from StepShape;
	---Purpose: Returns Value as PlusMinusTolerance (or Null if another type)

end ShapeToleranceSelect;
