-- Created on: 1995-07-18
-- Created by: Modelistation
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



generic class   GenExtPC from Extrema (Curve   as any; 
    	    	    	    	       Tool    as any;   --as ToolCurve(Curve)
				       POnC    as any; 
                                       Pnt     as any;
                                       Vec     as any)
				     
    	---Purpose: It calculates all the distances between a point
    	--          and a curve.
    	--          These distances can be minimum or maximum.


raises  NotDone      from StdFail,
    	OutOfRange   from Standard,
	TypeMismatch from Standard
	
private class PCF instantiates FuncExtPC from Extrema (Curve, Tool, POnC, Pnt, Vec);
	
is

    Create returns GenExtPC;
    

    Create (P: Pnt; C: Curve; NbU: Integer; TolU,TolF: Real)
    	returns GenExtPC;
      	---Purpose: It calculates all the distances.
        --          The function F(u)=distance(P,C(u)) has an extremum
        --          when g(u)=dF/du=0. The algorithm searchs all the
        --          zeros inside the definition range of the curve.
      	--          NbU is used to locate the close points to 
      	--          find the zeros.
      	--          Tol and TolU are used to decide to stop the 
      	--          iterations according to the following condition:
      	--          if n is the number of iterations,
      	--           abs(Un-Un-1) < TolU and abs(F(Un)-F(Un-1)) < Tol.


    Create (P: Pnt; C: Curve; NbU: Integer; Umin, Usup: Real; TolU,TolF: Real)
    	returns GenExtPC;
      	---Purpose: It calculates all the distances.
        --          The function F(u)=distance(P,C(u)) has an extremum
        --          when g(u)=dF/du=0. The algorithm searchs all the
        --          zeros inside the definition range of the curve.
      	--          NbU is used to locate the close points to 
      	--          find the zeros.
      	--          Zeros are searched between umin and usup.
      	--          Tol and TolU are used to decide to stop the 
      	--          iterations according to the following condition:
      	--          if n is the number of iterations,
      	--           abs(Un-Un-1) < TolU and abs(F(Un)-F(Un-1)) < Tol.



    Initialize(me: in out; C: Curve; NbU: Integer; TolU, TolF: Real)
    	---Purpose: sets the fields of the algorithm.
    is static;


    Initialize(me: in out; C: Curve; NbU: Integer; 
               Umin, Usup: Real; TolU, TolF: Real)
    	---Purpose: sets the fields of the algorithm.
    is static;

    Initialize(me: in out; C: Curve)
    	---Purpose: sets the fields of the algorithm.
    is static;

    Initialize(me: in out; NbU: Integer; Umin, Usup: Real; TolU, TolF: Real)
    	---Purpose: sets the fields of the algorithm.
    is static;


    Perform(me: in out; P: Pnt)
        ---Purpose: the algorithm is done with the point P.
        --          An exception is raised if the fields have not
        --          been initialized.  
    raises TypeMismatch from Standard
    is static;
    
    
    IsDone (me) returns Boolean
    	---Purpose: True if the distances are found.
    raises TypeMismatch from Standard
    is static;

    NbExt (me) returns Integer
    	---Purpose: Returns the number of extremum distances.
    raises TypeMismatch from Standard,
           NotDone from StdFail
	    	-- if IsDone(me)=False.
    	is static;
    
    SquareDistance (me; N: Integer) returns Real
    	---Purpose: Returns the value of the Nth extremum square distance.
    raises TypeMismatch from Standard,
    	   NotDone from StdFail,
	    	-- if IsDone(me)=False.
    	   OutOfRange from Standard
	    	-- if N < 1 or N > NbPoints(me).
    is static;


    IsMin (me; N: Integer) returns Boolean
    	---Purpose: Returns True if the Nth extremum distance is a
    	--          minimum.
    raises TypeMismatch from Standard,
    	   NotDone from StdFail,
	    	-- if IsDone(me)=False.
    	   OutOfRange from Standard
	    	-- if N < 1 or N > NbPoints(me).
    is static;


    Point (me; N: Integer) returns POnC
        ---C++: return const &
    	---Purpose: Returns the point of the Nth extremum distance.
    raises TypeMismatch from Standard,
    	   NotDone from StdFail,
	    	-- if IsDone(me)=False.
    	   OutOfRange from Standard
	    	-- if N < 1 or N > NbPoints(me).
    is static;



fields
    myDone :    Boolean;
    myInit:     Boolean;
    mynbsample: Integer;
    myumin:     Real;
    myusup:     Real;
    mytolu:     Real;
    mytolF:     Real;
    myF   :     PCF;

end GenExtPC;

