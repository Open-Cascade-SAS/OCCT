-- Created on: 1998-01-21
-- Created by: Kernel
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class AVLBaseNode from TCollection
    inherits TShared from MMgt
    uses AVLBaseNodePtr from TCollection,
    	 Side from TCollection
    is
    	Create(L,R : AVLBaseNodePtr from TCollection) returns mutable AVLBaseNode from TCollection;
	---C++: inline

    	SetChild(me : mutable; theNode : AVLBaseNodePtr from TCollection; theSide : Side from TCollection);
	---C++: inline

    	Height(myclass; ANode : AVLBaseNodePtr from TCollection) returns Integer;
    	RecursiveExtent(myclass;  ANode : AVLBaseNodePtr from TCollection) returns Integer;
	RecursiveTotalExtent(myclass;  ANode : AVLBaseNodePtr from TCollection) returns Integer;

    	Right(me) returns AVLBaseNodePtr from TCollection;
	---C++: inline
	---C++: return &

    	Left(me) returns AVLBaseNodePtr from TCollection;
	---C++: inline
	---C++: return &

    	Count(me) returns Integer;
	---C++: inline
	---C++: return &

    fields
      myLeft : AVLBaseNodePtr from TCollection is protected;
      myRight : AVLBaseNodePtr from TCollection is protected;
      myCount : Integer from Standard is protected;      
    end;
    
