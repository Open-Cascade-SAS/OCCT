-- Created on: 1992-02-18
-- Created by: Christophe MARION
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package HLRAlgo 
--- Purpose:        In order to have the precision required in
-- industrial design, drawings need to offer the
-- possibility of removing lines, which are hidden
-- in a given projection. To do this, the Hidden
-- Line Removal component provides two
 --   algorithms: HLRBRep_Algo and HLRBRep_PolyAlgo.
-- These algorithms remove or indicate lines
-- hidden by surfaces. For a given projection, they
-- calculate a set of lines characteristic of the
-- object being represented. They are also used
-- in conjunction with extraction utilities, which
-- reconstruct a new, simplified shape from a
-- selection of calculation results. This new shape
-- is made up of edges, which represent the lines
-- of the visualized shape in a plane. This plane is the projection plane.
-- HLRBRep_Algo takes into account the shape
-- itself. HLRBRep_PolyAlgo works with a
-- polyhedral simplification of the shape. When
-- you use HLRBRep_Algo, you obtain an exact
-- result, whereas, when you use
-- HLRBRep_PolyAlgo, you reduce computation
-- time but obtain polygonal segments.
uses
    Standard,
    StdFail,
    MMgt,
    TCollection,
    TColStd,
    TColgp,
    Intrv,
    gp,
    GeomAbs,
    TopAbs,
    TopBas,
    TopCnx,
    TopLoc,
    IntRes2d,
    IntCurveSurface

is
    class BiPoint;
    
    imported ListOfBPoint;
    
    imported ListIteratorOfListOfBPoint;

    class PolyShellData;

    class PolyInternalData;

    class PolyInternalSegment;

    class PolyInternalNode;

    class PolyData;

    class PolyHidingData;

    class TriangleData;

    imported Array1OfPHDat;
	
    imported transient class HArray1OfPHDat;
	
    imported Array1OfPISeg;
	
    imported transient class HArray1OfPISeg;
	
    imported Array1OfPINod;
	
    imported transient class HArray1OfPINod;
	
    imported Array1OfTData;
	
    imported transient class HArray1OfTData;
	
    class PolyAlgo;

    class EdgeStatus;

    class Projector;

    class Intersection;

    class Coincidence;

    class Interference             instantiates Interference from TopBas
    	(Intersection from HLRAlgo, 
	 Coincidence  from HLRAlgo);

    imported InterferenceList;

    imported ListIteratorOfInterferenceList;
	
    class EdgesBlock;

    class WiresBlock;

    class EdgeIterator;
	---Purpose: Iterator  on the  visible or  hidden  parts of  an
	--          EdgeStatus.
    
    UpdateMinMax (x,y,z : Real    from Standard;
                  Min   : Address from Standard;
                  Max   : Address from Standard);

    EnlargeMinMax (tol : Real    from Standard;
                   Min : Address from Standard;
                   Max : Address from Standard);

    InitMinMax (Big : Real    from Standard;
                Min : Address from Standard;
                Max : Address from Standard);

    EncodeMinMax (Min    : Address from Standard;
                  Max    : Address from Standard;
                  MinMax : Address from Standard);

    SizeBox (Min    : Address from Standard;
             Max    : Address from Standard)
    returns Real from Standard;

    DecodeMinMax (MinMax : Address from Standard;
                  Min    : Address from Standard;
                  Max    : Address from Standard);

    CopyMinMax (IMin : Address from Standard;
                IMax : Address from Standard;
                OMin : Address from Standard;
                OMax : Address from Standard);

    AddMinMax (IMin : Address from Standard;
               IMax : Address from Standard;
               OMin : Address from Standard;
               OMax : Address from Standard);

end HLRAlgo;
