-- File:	RWStepShape_RWNonManifoldSurfaceShapeRepresentation.cdl
-- Created:	Fri Dec 28 16:02:02 2001 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class RWNonManifoldSurfaceShapeRepresentation from RWStepShape

    ---Purpose: Read & Write tool for NonManifoldSurfaceShapeRepresentation

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    NonManifoldSurfaceShapeRepresentation from StepShape

is
    Create returns RWNonManifoldSurfaceShapeRepresentation from RWStepShape;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : NonManifoldSurfaceShapeRepresentation from StepShape);
	---Purpose: Reads NonManifoldSurfaceShapeRepresentation

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: NonManifoldSurfaceShapeRepresentation from StepShape);
	---Purpose: Writes NonManifoldSurfaceShapeRepresentation

    Share (me; ent : NonManifoldSurfaceShapeRepresentation from StepShape;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWNonManifoldSurfaceShapeRepresentation;
