-- Created on: 1993-01-09
-- Created by: CKY / Contract Toubro-Larsen ( TCD )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class HighLight from IGESGraph  inherits IGESEntity

        ---Purpose: defines IGESHighLight, Type <406> Form <20>
        --          in package IGESGraph
        --
        --          Attaches information that an entity is to be
        --          displayed in some system dependent manner

uses  Integer  -- no one specific type


is

        Create returns mutable HighLight;

        -- Specific Methods pertaining to the class

        Init (me               : mutable;
              nbProps          : Integer;
              aHighLightStatus : Integer);
        ---Purpose : This method is used to set the fields of the class
        --           HighLight
        --      - nbProps          : Number of property values (NP = 1)
        --      - aHighLightStatus : HighLight Flag

        NbPropertyValues(me) returns Integer;
        ---Purpose : returns the number of property values in <me>

        HighLightStatus(me) returns Integer;
        ---Purpose : returns 0 if <me> is not highlighted(default),
        --         1 if <me> is highlighted

        IsHighLighted(me) returns Boolean;
        ---Purpose : returns True if entity is highlighted

fields

--
-- Class    : IGESGraph_HighLight
--
-- Purpose  : Declaration of the variables specific to a
--            HighLight property.
--
-- Reminder : A HighLight property is defined by :
--                  - Number of property values (NP=1)
--                  - Flag
--

        theNbPropertyValues : Integer;

        theHighLight        : Integer;

end HighLight;
