-- Created on: 1992-10-19
-- Created by: Laurent BUCHARD
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

generic class Polygon2dGen from IntCurve ( 
    TheCurve         as any;
    TheCurveTool     as any) -- as CurveTool from IntCurve(TheCurve)

	---Purpose: Describe a polyline  as  a topology to compute the
	--          interference beetween two polylines 2 dimension.

        ---Level: Internal

inherits Polygon2d from Intf

uses    Pnt2d              from gp,
    	Box2d              from Bnd,
    	Array1OfPnt2d      from TColgp,
        Array1OfReal       from TColStd,
        Array1OfInteger    from TColStd,
        Domain             from IntRes2d

raises  OutOfRange from Standard

is  

    Create         (Curve       : TheCurve;
    	    	    NbPnt       : Integer  from Standard;
		    Domain      : Domain   from IntRes2d;
    	    	    Tol         : Real     from Standard) 
		    
		    ---Purpose: Compute a polygon on the domain of the curve.
		    
		    
    	    	    returns Polygon2dGen from IntCurve;

    Create         (Curve       : TheCurve;
    	    	    NbPnt       : Integer  from Standard;
		    Domain      : Domain   from IntRes2d;
    	    	    Tol         : Real     from Standard;
		    OtherBox    : Box2d    from Bnd)
		    
		    ---Purpose: Compute a polygon on the domain of the
		    --          curve.   parameters of  the  begin and
		    --          end of the curve (and its polygon) are
		    --          adjusted to lie in the OtherBox.
		    
    	    	    returns Polygon2dGen from IntCurve;


    ComputeWithBox(me       : in out; 
                   Curve    : TheCurve;
		   OtherBox : Box2d  from Bnd)
		   
		   ---Purpose: The current polygon is modified if most
		   --          of the  points of the  polygon  are are
		   --          outside  the  box  <OtherBox>.  In this
		   --          situation, bounds are computed to build
		   --          a polygon inside or near the OtherBox.
                   is static;

    DeflectionOverEstimation(me)
		   returns Real from Standard
		   ---C++: inline
		   is redefined virtual;

    SetDeflectionOverEstimation(me: in out; x:Real from Standard)
                    ---C++: inline
		    is static;

    Closed         (me : in out; clos : Boolean from Standard)
    	            ---C++: inline
		    is static;

    NbSegments     (me)
    	    	    returns Integer
		    ---C++: inline
    	    	    is redefined virtual;
    ---Purpose: Give the number of Segments in the polyline.

    Segment (me; theIndex : in Integer from Standard;
                 theBegin, theEnd : in out Pnt2d from gp)
        raises OutOfRange from Standard is redefined virtual;
    ---Purpose: Returns the points of the segment <Index> in the Polygon.

-- Implementation : 


   InfParameter(me) 
   
    	---Purpose: Returns the parameter (On the curve)
    	--          of the first point of the Polygon
   
    	returns Real from Standard
	---C++: inline
	is static;

   SupParameter(me) 

       	---Purpose: Returns the parameter (On the curve)
    	--          of the last point of the Polygon
   
    	returns Real from Standard
	---C++: inline
	is static;


   AutoIntersectionIsPossible(me) 
       returns Boolean from Standard
       is static;

   ApproxParamOnCurve(me; 
                      Index       : in  Integer from Standard;
		      ParamOnLine : in  Real    from Standard)
    	    	      
                      returns Real      from Standard
    	    	     
		      raises OutOfRange from Standard
    	    	      is static;

            ---Purpose: Give an approximation of the parameter on the curve 
            --          according to the discretization of the Curve.

     
    CalculRegion  (me; 
    	    	   x  :  Real  from  Standard  ; 
		   y  :  Real  from  Standard  ;
    	    	   x1 :  Real  from  Standard  ; 
    	    	   x2 :  Real  from  Standard  ; 
		   y1 :  Real  from  Standard  ;
		   y2 :  Real  from  Standard  ) 
	returns  Integer  from  Standard  ;	   
	---C++: inline
		 	
    Dump           (me)
    	is static;


fields  TheDeflection : Real                 from Standard;
    	NbPntIn       : Integer              from Standard;
        TheMaxNbPoints: Integer              from Standard;
    	ThePnts       : Array1OfPnt2d        from TColgp;
        TheParams     : Array1OfReal         from TColStd;
        TheIndex      : Array1OfInteger      from TColStd;
        ClosedPolygon : Boolean              from Standard;

	--- To compute an approximate parameter on the Curve
	--  
	Binf          : Real                 from Standard;
	Bsup          : Real                 from Standard;

end Polygon2dGen;
