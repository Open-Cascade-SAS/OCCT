-- Created on: 1993-06-22
-- Created by: Jean Louis FRENKEL, Gerard Gras.
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


package GGraphic2d

	---Version:

	---Purpose: This package permits the creation of 2d graphic curves
	--          and set of curves in a   in a visualiser.
	--	    It moved from the Graphic2d package to this package
	--	    since it required services from the UL GEOMETRY
	--	    

	---Keywords: Drawer, View, Graphic Object, Primitive, Line,
	--	     Circle, Polyline, Ellips, Curve, Image, Text, HidingText,
	--	     FramedText, Paragraph
	---Warning:
	---References:

uses
        Graphic2d,
	Aspect,
	Geom2d,
	Image,
	MMgt,
	gp,
	OSD,
	Quantity,
	TCollection,
	TColStd,
	TShort,
	TColGeom2d

is
        class Curve ;
	---Category: Set of primitive curves
	--           
	class SetOfCurves;
	---Category: Set Of Graphic primitives


	-----------------------
	-- Category: Exceptions
	-----------------------


	exception CurveDefinitionError inherits OutOfRange;	
	---Category: Exceptions
		
end GGraphic2d;

