-- Created by: DAUTRY Philippe
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

--      	----------------------------

---Version:	0.0
--Version	Date		Purpose
--		0.0	Aug 27 1997	Creation


class XLinkIterator from TDocStd 

	---Purpose: Iterates on Reference attributes.

uses Document from TDocStd,
     XLink     from TDocStd,
     XLinkPtr  from TDocStd

raises

    NoMoreObject from Standard

is

    Create
    returns XLinkIterator from TDocStd;
	---Purpose: Returns an empty iterator;

    Create (D : Document from TDocStd)
    returns XLinkIterator from TDocStd;
    	---Purpose: Creates an iterator on Reference of <D>.
    
    Initialize (me  : in out; D : Document from TDocStd);
    	---Purpose: Restarts an iteration with <D>.
    
    More (me) returns Boolean;
	---Purpose: Returns True if there is a current Item in the
	--          iteration.
	--          
	---C++: inline
    
    Next (me : in out)
    	raises NoMoreObject from Standard;
    	---Purpose: Move to the next item; raises if there is no more item.
    
    Value (me) returns XLinkPtr from TDocStd;
	---Purpose: Returns the current item; a null handle if there is none.
	--          
	---C++: inline

    Init (me : in out; D : Document from TDocStd) is private;


fields

    myValue : XLinkPtr from TDocStd;

end XLinkIterator;
