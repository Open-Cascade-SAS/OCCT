-- File:        ProductDefinition.cdl
-- Created:     Mon Dec  4 12:02:29 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWProductDefinition from RWStepBasic

	---Purpose : Read & Write Module for ProductDefinition

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     ProductDefinition from StepBasic,
     EntityIterator from Interface

is

	Create returns RWProductDefinition;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable ProductDefinition from StepBasic);

	WriteStep (me; SW : in out StepWriter; ent : ProductDefinition from StepBasic);

	Share(me; ent : ProductDefinition from StepBasic; iter : in out EntityIterator);

end RWProductDefinition;
