-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class CsgSelect from StepShape 

    -- inherits SelectType from StepData

	-- <CsgSelect> is an EXPRESS Select Type construct translation.
	-- it gathers : BooleanResult, CsgPrimitive

uses

	BooleanResult,
	CsgPrimitive
is

	Create returns CsgSelect;
	---Purpose : Returns a CsgSelect SelectType

    	SetTypeOfContent(me : in out; aTypeOfContent : Integer);

	TypeOfContent(me) returns Integer;
	--        1 -> BooleanResult
	--        2 -> CsgPrimitive
	--        0 else
	
	BooleanResult (me) returns any BooleanResult;
	---Purpose : returns Value as a BooleanResult (Null if another type)

    	SetBooleanResult (me : in out;aBooleanResult : BooleanResult from StepShape);
	
	CsgPrimitive (me) returns CsgPrimitive;
	---Purpose : returns Value as a CsgPrimitive (Null if another type)

    	SetCsgPrimitive (me : in out; aCsgPrimitive : CsgPrimitive from StepShape);
	
fields

    theBooleanResult : BooleanResult from StepShape;
    theCsgPrimitive  : CsgPrimitive  from StepShape;  -- a Select Type
    theTypeOfContent : Integer       from Standard;

end CsgSelect;

