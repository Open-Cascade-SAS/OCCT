-- Created on: 2006-08-07
-- Created by: Galina KULIKOVA
-- Copyright (c) 2006-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class FaceDivideArea from ShapeUpgrade inherits FaceDivide from ShapeUpgrade

	---Purpose: Divides face by max area criterium.

uses
    Face from TopoDS

is

    Create returns FaceDivideArea from ShapeUpgrade; 
        ---Purpose: Creates empty  constructor.

    Create (F : Face from TopoDS) returns FaceDivideArea from ShapeUpgrade;
    
    Perform (me: mutable) returns Boolean is redefined;
        ---Purpose: Performs splitting and computes the resulting shell
	--          The context is used to keep track of former splittings
    
    MaxArea(me: mutable) returns Real;
    ---C++: inline
    ---C++: return &
    ---Purpose:Set max area allowed for faces
     
fields

    myMaxArea : Real;

end FaceDivideArea;
