-- File:        TopologicalRepresentationItem.cdl
-- Created:     Mon Dec  4 12:02:32 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWTopologicalRepresentationItem from RWStepShape

	---Purpose : Read & Write Module for TopologicalRepresentationItem

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     TopologicalRepresentationItem from StepShape

is

	Create returns RWTopologicalRepresentationItem;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable TopologicalRepresentationItem from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : TopologicalRepresentationItem from StepShape);

end RWTopologicalRepresentationItem;
