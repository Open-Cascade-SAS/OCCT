-- File:	BOPTColStd_ShapeWithRank.cdl
-- Created:	Fri Jun  8 17:12:40 2001
-- Author:	Peter KURNEV
--		<pkv@irinox>
---Copyright:	 Matra Datavision 2001


class ShapeWithRank from BOPTColStd 

	---Purpose: 
    	--  The auxiliary class provides structure to store a shape 
    	--  and its rank 
    	--- 
uses
    Shape from TopoDS

--raises

is 
    Create   
    	returns ShapeWithRank from BOPTColStd; 
    ---Purpose:   
    -- Empty constructor
    ---     
    SetShape(me:out;   
    	aS: Shape from TopoDS); 
    ---Purpose:   
    -- Modifier
    ---      
    SetRank(me:out; 
	aR:  Integer from Standard); 
    ---Purpose:   
    -- Modifier
    ---   
    Shape(me) 
    	returns Shape from TopoDS;   	    	    	
    ---C++: return  const & 
    ---Purpose:   
    -- Selector
    --- 
    Rank(me) 
	returns Integer from Standard; 
    ---Purpose:   
    -- Selector
    --- 
    HashCode(me; 
    	    Upper:Integer from Standard) 
    	returns Integer from Standard; 
    ---Purpose: Returns a HasCode value  for  the  Key <K>  in the
    --          range 0..Upper.
    -- 
    IsEqual(me; 
    	    Other:ShapeWithRank from BOPTColStd)		 
    	returns Boolean from Standard;	     
    ---Purpose: Returns True  when the two  keys are the same. Two
    --          same  keys  must   have  the  same  hashcode,  the
    --          contrary is not necessary.
    -- 
     
fields 
    myShape :  Shape from TopoDS; 
    myRank  :  Integer from Standard; 
     
end ShapeWithRank;
