-- Created on: 1999-04-15
-- Created by: Denis PASCAL
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package MDocStd 

	---Purpose: Drivers for TDocStd_Document

uses TColStd, TCollection, PCollection, PTColStd,
     CDM, PCDM,  
     TDF, PDF, MDF,
     TDocStd, PDocStd

is

    ---Purpose: Standard CAF Document drivers
    --          =============================


    class DocumentStorageDriver;
     
    class DocumentRetrievalDriver;
    
    
    ---Purpose: External Reference Attribute  drivers
    --          =====================================

    class XLinkStorageDriver;
    
    class XLinkRetrievalDriver;
    
--    class PersistentMap instantiates Map from TCollection( Persistent from Standard,
--    	                                                   MapPersistentHasher from PTColStd);

--    class DocEntryList instantiates List from TCollection (AsciiString from TCollection);
    

    AddStorageDrivers(aDriverSeq : ASDriverHSequence from MDF; theMessageDriver : MessageDriver from CDM);
	---Purpose: Adds the attribute storage driver(s) to <aDriverSeq>.

    AddRetrievalDrivers(aDriverSeq : ARDriverHSequence from MDF; theMessageDriver : MessageDriver from CDM);
	---Purpose: Adds the attribute retrieval driver(s) to <aDriverSeq>.
    
    
--    WeightWatcher(aSource : Data from TDF;
--                  aReloc   : SRelocationTable from MDF;
--                  aEntry : DocEntryList from MDocStd);
--    ---Purpose: suppresses the geometries  of the shapes from the XLink
--    --          associated to  <aEntry>

    ---Purpose: Factory method
    --          ==============
    
    Factory(aGUID: GUID from Standard)
    returns Transient from Standard;

end MDocStd;
