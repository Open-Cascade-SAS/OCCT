-- Created on: 2002-12-12
-- Created by: data exchange team
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class CurveElementSectionDerivedDefinitions from StepElement
inherits CurveElementSectionDefinition from StepElement

    ---Purpose: Representation of STEP entity CurveElementSectionDerivedDefinitions

uses
    HAsciiString from TCollection,
    HArray1OfMeasureOrUnspecifiedValue from StepElement,
    HArray1OfReal from TColStd,
    MeasureOrUnspecifiedValue from StepElement,
    HArray1OfMeasureOrUnspecifiedValue from StepElement

is
    Create returns CurveElementSectionDerivedDefinitions from StepElement;
	---Purpose: Empty constructor

    Init (me: mutable; aCurveElementSectionDefinition_Description: HAsciiString from TCollection;
                       aCurveElementSectionDefinition_SectionAngle: Real;
                       aCrossSectionalArea: Real;
                       aShearArea: HArray1OfMeasureOrUnspecifiedValue from StepElement;
                       aSecondMomentOfArea: HArray1OfReal from TColStd;
                       aTorsionalConstant: Real;
                       aWarpingConstant: MeasureOrUnspecifiedValue from StepElement;
                       aLocationOfCentroid: HArray1OfMeasureOrUnspecifiedValue from StepElement;
                       aLocationOfShearCentre: HArray1OfMeasureOrUnspecifiedValue from StepElement;
                       aLocationOfNonStructuralMass: HArray1OfMeasureOrUnspecifiedValue from StepElement;
                       aNonStructuralMass: MeasureOrUnspecifiedValue from StepElement;
                       aPolarMoment: MeasureOrUnspecifiedValue from StepElement);
	---Purpose: Initialize all fields (own and inherited)

    CrossSectionalArea (me) returns Real;
	---Purpose: Returns field CrossSectionalArea
    SetCrossSectionalArea (me: mutable; CrossSectionalArea: Real);
	---Purpose: Set field CrossSectionalArea

    ShearArea (me) returns HArray1OfMeasureOrUnspecifiedValue from StepElement;
	---Purpose: Returns field ShearArea
    SetShearArea (me: mutable; ShearArea: HArray1OfMeasureOrUnspecifiedValue from StepElement);
	---Purpose: Set field ShearArea

    SecondMomentOfArea (me) returns HArray1OfReal from TColStd;
	---Purpose: Returns field SecondMomentOfArea
    SetSecondMomentOfArea (me: mutable; SecondMomentOfArea: HArray1OfReal from TColStd);
	---Purpose: Set field SecondMomentOfArea

    TorsionalConstant (me) returns Real;
	---Purpose: Returns field TorsionalConstant
    SetTorsionalConstant (me: mutable; TorsionalConstant: Real);
	---Purpose: Set field TorsionalConstant

    WarpingConstant (me) returns MeasureOrUnspecifiedValue from StepElement;
	---Purpose: Returns field WarpingConstant
    SetWarpingConstant (me: mutable; WarpingConstant: MeasureOrUnspecifiedValue from StepElement);
	---Purpose: Set field WarpingConstant

    LocationOfCentroid (me) returns HArray1OfMeasureOrUnspecifiedValue from StepElement;
	---Purpose: Returns field LocationOfCentroid
    SetLocationOfCentroid (me: mutable; LocationOfCentroid: HArray1OfMeasureOrUnspecifiedValue from StepElement);
	---Purpose: Set field LocationOfCentroid

    LocationOfShearCentre (me) returns HArray1OfMeasureOrUnspecifiedValue from StepElement;
	---Purpose: Returns field LocationOfShearCentre
    SetLocationOfShearCentre (me: mutable; LocationOfShearCentre: HArray1OfMeasureOrUnspecifiedValue from StepElement);
	---Purpose: Set field LocationOfShearCentre

    LocationOfNonStructuralMass (me) returns HArray1OfMeasureOrUnspecifiedValue from StepElement;
	---Purpose: Returns field LocationOfNonStructuralMass
    SetLocationOfNonStructuralMass (me: mutable; LocationOfNonStructuralMass: HArray1OfMeasureOrUnspecifiedValue from StepElement);
	---Purpose: Set field LocationOfNonStructuralMass

    NonStructuralMass (me) returns MeasureOrUnspecifiedValue from StepElement;
	---Purpose: Returns field NonStructuralMass
    SetNonStructuralMass (me: mutable; NonStructuralMass: MeasureOrUnspecifiedValue from StepElement);
	---Purpose: Set field NonStructuralMass

    PolarMoment (me) returns MeasureOrUnspecifiedValue from StepElement;
	---Purpose: Returns field PolarMoment
    SetPolarMoment (me: mutable; PolarMoment: MeasureOrUnspecifiedValue from StepElement);
	---Purpose: Set field PolarMoment

fields
    theCrossSectionalArea: Real;
    theShearArea: HArray1OfMeasureOrUnspecifiedValue from StepElement;
    theSecondMomentOfArea: HArray1OfReal from TColStd;
    theTorsionalConstant: Real;
    theWarpingConstant: MeasureOrUnspecifiedValue from StepElement;
    theLocationOfCentroid: HArray1OfMeasureOrUnspecifiedValue from StepElement;
    theLocationOfShearCentre: HArray1OfMeasureOrUnspecifiedValue from StepElement;
    theLocationOfNonStructuralMass: HArray1OfMeasureOrUnspecifiedValue from StepElement;
    theNonStructuralMass: MeasureOrUnspecifiedValue from StepElement;
    thePolarMoment: MeasureOrUnspecifiedValue from StepElement;

end CurveElementSectionDerivedDefinitions;
