-- Created on: 2002-02-07
-- Created by: Igor FEOKTISTOV
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ReShaper from QANewModTopOpe inherits TShared from  MMgt 
    	---Purpose: to remove  "floating" objects from compound.
	-- "floating" objects are wires, edges, vertices that do not belong
	-- solids, shells or faces.

uses 
    Shape from TopoDS, 
    HSequenceOfShape  from  TopTools, 
    MapOfShape  from  TopTools 
is 
 
    Create(TheInitialShape  :  Shape from TopoDS) 
     
    returns  mutable  ReShaper; 
     
    Create(TheInitialShape  :  Shape from TopoDS;   
    	   TheMap  :  MapOfShape  from  TopTools) 
     
    returns  mutable  ReShaper; 
     
    Create(TheInitialShape  :  Shape from TopoDS;   
           TheShapeToBeRemoved  : HSequenceOfShape  from  TopTools) 
     
    returns  mutable  ReShaper; 
     
    Remove(me  :  mutable;  TheS  :  Shape from TopoDS); 
     
    Perform(me  :  mutable); 
     
    Clear(me  :  mutable);  
    ---Purpose:  to  clear  all  added  for  removing  shapes  from  inner  map.
     
    GetResult(me)  returns  Shape  from  TopoDS; 
	---C++: return const &
	---C++: alias "Standard_EXPORT operator TopoDS_Shape() const;"
     
fields 
 
    myInitShape  :  Shape  from  TopoDS; 
    myResult     :  Shape  from  TopoDS;  
    myMap        :  MapOfShape  from  TopTools;  
    
end;    
