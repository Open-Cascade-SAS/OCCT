-- Created on: 1999-08-31
-- Created by: Pavel DURANDIN
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



private class Tool from ShapeUpgrade inherits TShared from MMgt

	---Purpose: Tool is a root class for splitting classes
	--          Provides context for recording changes, basic 
    	--          precision value and limit (minimal and maximal) 
    	--          values for tolerances

uses

    ReShape from ShapeBuild

is

    Create returns Tool from ShapeUpgrade;
    	---Purpose: Empty constructor
	    
    Set (me: mutable; tool: Tool from ShapeUpgrade);
    	---Purpose: Copy all fields from another Root object
	
    SetContext (me: mutable; context : ReShape from ShapeBuild);
	---Purpose: Sets context
	---C++: inline
	
    Context (me) returns ReShape from ShapeBuild;
    	---Purpose: Returns context 
	---C++: inline
	
    SetPrecision (me: mutable; preci: Real);
    	---Purpose: Sets basic precision value
	---C++: inline
    
    Precision (me) returns Real;
    	---Purpose: Returns basic precision value
	---C++: inline
	
    SetMinTolerance (me: mutable; mintol: Real);
    	---Purpose: Sets minimal allowed tolerance
	---C++: inline
    
    MinTolerance (me) returns Real;
    	---Purpose: Returns minimal allowed tolerance
	---C++: inline
	
    SetMaxTolerance (me: mutable; maxtol: Real);
    	---Purpose: Sets maximal allowed tolerance
	---C++: inline
    
    MaxTolerance (me) returns Real;
    	---Purpose: Returns maximal allowed tolerance
	---C++: inline
    
    LimitTolerance (me; toler: Real) returns Real;
    	---Purpose: Returns tolerance limited by [myMinTol,myMaxTol]
	---C++: inline

fields

    myContext  : ReShape from ShapeBuild;
    myPrecision: Real;       -- basic precision
    myMinTol   : Real;       -- minimal allowed tolerance
    myMaxTol   : Real;       -- maximal allowed tolerance

end Tool;
