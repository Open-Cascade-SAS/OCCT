-- Created on: 1994-09-02
-- Created by: Frederic MAUPAS
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class MakeEllipse from GeomToStep inherits Root from GeomToStep

    ---Purpose: This class implements the mapping between classes 
    --          Ellipse from Geom, and Circ from gp, and the class
    --          Ellipse from StepGeom which describes a Ellipse from
    --          Prostep. 
  
uses Elips from gp,
     Elips2d from gp,
     Ellipse from Geom,
     Ellipse from Geom2d,
     Ellipse from StepGeom
     
raises NotDone from StdFail
     
is 

Create ( C : Elips from gp ) returns MakeEllipse;

Create ( C : Ellipse from Geom ) returns MakeEllipse;

Create ( C : Ellipse from Geom2d ) returns MakeEllipse;

Value (me) returns Ellipse from StepGeom
    raises NotDone
    is static;
    ---C++: return const&
  
fields

    theEllipse : Ellipse from StepGeom;
    	-- The solution from StepGeom
    	
end MakeEllipse;


