-- Created on: 1994-02-17
-- Created by: Bruno DUMORTIER
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Generator from GeomFill inherits Profiler from GeomFill

        ---Purpose: Create a surface using generating lines.  Inherits
        --          profiler.  The  surface will be  a  BSplineSurface
        --          passing  by   all  the  curves  described  in  the
        --          generator. The VDegree of the resulting surface is
        --          1.


uses
    Surface from Geom


raises
    NotDone     from StdFail,
    DomainError from Standard

is
    Create returns Generator from GeomFill;
    
    Perform(me   : in out ;
            PTol : in Real from Standard)
	---Purpose: Converts all curves to BSplineCurves.
	--          Set them to the common profile.
	--          Compute the surface (degv = 1).
	--          <PTol> is used to compare 2 knots.
    is redefined;
    
    Surface(me)
    returns Surface from Geom
    	---C++: return const&
    	---C++: inline
    is static;
    
    
fields
    mySurface : Surface from Geom;

end Generator;
