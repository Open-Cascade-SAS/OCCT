-- Created by: DAUTRY Philippe
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

--      	--------------

---Version:	0.0
--Version	Date		Purpose
--		0.0	Mar 13 1997	Creation


class Tool from MDF

	---Purpose: A tool to translate...

uses

    Label                  from TDF,
    Data                   from TDF,
    Data                   from PDF,
    HAttributeArray1       from PDF,
    TypeARDriverMap        from MDF,
    TypeASDriverMap        from MDF,
    ARDriverTable          from MDF,
    ASDriverTable          from MDF,
    RRelocationTable       from MDF,
    SRelocationTable       from MDF,
    Integer                from Standard,
    HArray1OfInteger       from PColStd,
    TransientPersistentMap from PTColStd

-- raises

is

    WriteLabels(myclass;
    	  aSource : Data from TDF;
	  aTarget : Data from PDF;
	  aDriverMap    : TypeASDriverMap from MDF;
	  aReloc        : SRelocationTable from MDF);
	---Purpose: Writes the labels with empty attributes.

    WriteLabels(myclass;
    	  aSourceLab    : Label from TDF;
	  theLabels     : HArray1OfInteger from PColStd;
	  theAttributes : HAttributeArray1 from PDF;
	  aDriverMap    : TypeASDriverMap from MDF;
	  aReloc        : SRelocationTable from MDF;
	  labAlloc      : in out Integer from Standard;
	  attAlloc      : in out Integer from Standard);
	---Purpose: Used for recursivity.

    WriteAttributes(myclass;
	aDriverMap    : TypeASDriverMap from MDF;
    	aReloc        : SRelocationTable from MDF);
	---Purpose: Writes attributes content.



    ReadLabels(myclass;
    	  aSource : Data from PDF;
	  aTarget : Data from TDF;
	  aDriverMap    : TypeARDriverMap from MDF;
	  aReloc        : RRelocationTable from MDF);
	---Purpose:  Reads the labels abd adds empty attributes to them.

    ReadLabels(myclass;
    	  anIns         : in out Label from TDF;
	  theLabels     : HArray1OfInteger from PColStd;
	  theAttributes : HAttributeArray1 from PDF;
	  aDriverMap    : TypeARDriverMap from MDF;
	  aReloc        : RRelocationTable from MDF;
	  labRead       : in out Integer from Standard;
	  attRead       : in out Integer from Standard);
	---Purpose: Used for recursivity.

    ReadAttributes(myclass;
	aDriverMap    : TypeARDriverMap from MDF;
    	aReloc        : RRelocationTable from MDF);
	---Purpose: Reads attributes content and paste them.

end Tool;
