-- Created on: 2001-01-06
-- Created by: OCC Team
-- Copyright (c) 2001-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class PrinterOStream from Message inherits Printer from Message

    ---Purpose: Implementation of a message printer associated with an ostream
    --          The ostream may be either externally defined one (e.g. cout),
    --          or file stream maintained internally (depending on constructor).

uses

    Address        from Standard,
    OStream        from Standard,
    Gravity        from Message,
    AsciiString    from TCollection,
    ExtendedString from TCollection    

is

    Create (theTraceLevel: Gravity from Message = Message_Info)
    returns PrinterOStream from Message;
    	---Purpose: Empty constructor, defaulting to cout
    
    Create (theFileName: CString; theDoAppend: Boolean;
            theTraceLevel: Gravity from Message = Message_Info)
    returns PrinterOStream from Message;
    	---Purpose: Create printer for output to a specified file.
    	--          The option theDoAppend specifies whether file should be
    	--          appended or rewritten.
    	--          For specific file names (cout, cerr) standard streams are used
    
    Close (me: mutable);
        ---C++: alias ~
    	---Purpose: Flushes the output stream and destroys it if it has been
    	--          specified externally with option doFree (or if it is internal
        --          file stream)
	
    GetTraceLevel (me) returns Gravity from Message;
    	---C++: inline
    	---Purpose: Return trace level used for filtering messages;
	--          messages with lover gravity will be ignored.

    SetTraceLevel (me: mutable; theTraceLevel: Gravity from Message);
    	---C++: inline
    	---Purpose: Set trace level used for filtering messages.
    	--          By default, trace level is Message_Info, so that 
    	--          all messages are output

    GetUseUtf8 (me) returns Boolean;
    	---Purpose: Returns option to convert non-Ascii symbols to UTF8 encoding
    	---C++: inline

    SetUseUtf8 (me: mutable; useUtf8: Boolean);
    	---Purpose: Sets option to convert non-Ascii symbols to UTF8 encoding
    	---C++: inline

    GetStream (me) returns OStream;
    	---Purpose: Returns reference to the output stream
	---C++: return &
    	---C++: inline
    
    Send (me; theString : CString; theGravity: Gravity from Message;
	      putEndl: Boolean = Standard_True) is redefined;
    	---Purpose: Puts a message to the current stream
	--          if its gravity is equal or greater
	--          to the trace level set by SetTraceLevel()
	      
    Send (me; theString : AsciiString from TCollection;
              theGravity: Gravity from Message;
	      putEndl: Boolean = Standard_True) is redefined;
    	---Purpose: Puts a message to the current stream
	--          if its gravity is equal or greater
	--          to the trace level set by SetTraceLevel()
	      
    Send (me; theString : ExtendedString from TCollection;
              theGravity: Gravity from Message;
	      putEndl: Boolean = Standard_True) is redefined;
    	---Purpose: Puts a message to the current stream
	--          if its gravity is equal or greater
	--          to the trace level set by SetTraceLevel()
	--          Non-Ascii symbols are converted to UTF-8 if UseUtf8
        --          option is set, else replaced by symbols '?'
	      
fields

    myTraceLevel: Gravity from Message;
    myStream:     Address from Standard; -- pointer to OStream 
    myIsFile:     Boolean from Standard;
    myUseUtf8:    Boolean from Standard;

end PrinterOStream;
