-- Created on: 1997-07-29
-- Created by: Denis PASCAL
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class NoteBook from TDataStd inherits Attribute from TDF

    	---Purpose: NoteBook Object attribute


uses Attribute       from TDF,
     Label           from TDF,
     Real            from TDataStd,
     Integer         from TDataStd,
     GUID            from Standard,
     DataSet         from TDF,
     RelocationTable from TDF

is  

    ---Purpose: class methods
    --          =============
    
    Find (myclass; current : Label from TDF; N : in out NoteBook from TDataStd)
    ---Purpose: try to retrieve a NoteBook attribute at <current> label
    --           or in  fathers  label of  <current>. Returns True  if
    --          found and set <N>.
    returns Boolean from Standard;
    
    New (myclass; label : Label from TDF)   
    ---Purpose:  Create  an  enpty   NoteBook attribute,  located  at
    --          <label>. Raises if <label> has attribute
    returns NoteBook from TDataStd;
    
    GetID (myclass)   
    ---C++: return const &  
    returns GUID from Standard;
    ---Purpose: NoteBook methods
    --          ===============

    Create
    returns mutable NoteBook from TDataStd; 
    

    Append (me : mutable; value  : Real    from Standard; 
                          isExported : Boolean from Standard = Standard_False)    
    ---Purpose:  Tool to Create  an  Integer  attribute from  <value>,
    --          Insert it in   a  new son  label   of <me>. The   Real
    --          attribute is returned.
    returns Real from TDataStd;
    
    Append (me : mutable; value  : Integer from Standard; 
                          isExported : Boolean from Standard = Standard_False)    
    ---Purpose: Tool to Create  an Real attribute from <value>, Insert
    --          it  in a new son label  of <me>. The Integer attribute
    --          is returned.
    returns Integer from TDataStd;

    
    ---Category: methodes de TDF_Attribute
    --           =========================

    ID (me)
    ---C++: return const & 
    returns GUID from Standard;

    Restore (me: mutable; with : Attribute from TDF);

    NewEmpty (me)
    returns mutable Attribute from TDF;

    Paste (me; into : mutable Attribute from TDF;
	       RT   : mutable RelocationTable from TDF);    

    Dump(me; anOS : in out OStream from Standard)
    	returns OStream from Standard
    	is redefined;
	---C++: return &
    
end NoteBook;
