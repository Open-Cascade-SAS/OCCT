-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class BooleanResult from StepShape 

inherits GeometricRepresentationItem from StepGeom

uses

	BooleanOperator from StepShape, 
	BooleanOperand from StepShape, 
	HAsciiString from TCollection
is

	Create returns mutable BooleanResult;
	---Purpose: Returns a BooleanResult


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aOperator : BooleanOperator from StepShape;
	      aFirstOperand : BooleanOperand from StepShape;
	      aSecondOperand : BooleanOperand from StepShape) is virtual;

	-- Specific Methods for Field Data Access --

	SetOperator(me : mutable; aOperator : BooleanOperator);
	Operator (me) returns BooleanOperator;
	SetFirstOperand(me : mutable; aFirstOperand : BooleanOperand);
	FirstOperand (me) returns BooleanOperand;
	SetSecondOperand(me : mutable; aSecondOperand : BooleanOperand);
	SecondOperand (me) returns BooleanOperand;

fields

	anOperator : BooleanOperator from StepShape; -- an Enumeration
	firstOperand : BooleanOperand from StepShape; -- a SelectType
	secondOperand : BooleanOperand from StepShape; -- a SelectType

end BooleanResult;
