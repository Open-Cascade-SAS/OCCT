-- File:	MDataStd_ExpressionStorageDriver.cdl
-- Created:	Thu Aug  7 17:09:27 1997
-- Author:	PASCAL Denis
---Copyright:	 Matra Datavision 1997

class ExpressionStorageDriver from MDataStd inherits ASDriver from MDF

	---Purpose: 

uses SRelocationTable from MDF,
     Attribute        from TDF,
     Attribute        from PDF, 
     MessageDriver    from CDM


is

    Create(theMessageDriver : MessageDriver from CDM) 
    returns mutable ExpressionStorageDriver from MDataStd;


    VersionNumber(me) returns Integer from Standard;
	---Purpose: Returns the version number from which the driver
	--          is available: 0.

    SourceType(me) returns Type from Standard;
	---Purpose: Returns the type: Integer from TDataStd.

    NewEmpty (me) returns mutable Attribute from PDF;


    Paste(me; Source     :         Attribute from TDF;
    	      Target     : mutable Attribute from PDF;
    	      RelocTable : SRelocationTable from MDF);


end ExpressionStorageDriver;

