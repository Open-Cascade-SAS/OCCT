-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class CurveStyleFontSelect from StepVisual inherits SelectType from StepData

	-- <CurveStyleFontSelect> is an EXPRESS Select Type construct translation.
	-- it gathers : CurveStyleFont, PreDefinedCurveFont, ExternallyDefinedCurveFont

uses

	CurveStyleFont,
	PreDefinedCurveFont,
	ExternallyDefinedCurveFont
is

	Create returns CurveStyleFontSelect;
	---Purpose : Returns a CurveStyleFontSelect SelectType

	CaseNum (me; ent : Transient) returns Integer;
	---Purpose: Recognizes a CurveStyleFontSelect Kind Entity that is :
	--        1 -> CurveStyleFont
	--        2 -> PreDefinedCurveFont
	--        3 -> ExternallyDefinedCurveFont
	--        0 else

	CurveStyleFont (me) returns any CurveStyleFont;
	---Purpose : returns Value as a CurveStyleFont (Null if another type)

	PreDefinedCurveFont (me) returns any PreDefinedCurveFont;
	---Purpose : returns Value as a PreDefinedCurveFont (Null if another type)

	ExternallyDefinedCurveFont (me) returns any ExternallyDefinedCurveFont;
	---Purpose : returns Value as a ExternallyDefinedCurveFont (Null if another type)


end CurveStyleFontSelect;

