-- File:	StepRepr_PropertyDefinitionRelationship.cdl
-- Created:	Thu Dec 12 16:04:59 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class PropertyDefinitionRelationship from StepRepr
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity PropertyDefinitionRelationship

uses
    HAsciiString from TCollection,
    PropertyDefinition from StepRepr

is
    Create returns PropertyDefinitionRelationship from StepRepr;
	---Purpose: Empty constructor

    Init (me: mutable; aName: HAsciiString from TCollection;
                       aDescription: HAsciiString from TCollection;
                       aRelatingPropertyDefinition: PropertyDefinition from StepRepr;
                       aRelatedPropertyDefinition: PropertyDefinition from StepRepr);
	---Purpose: Initialize all fields (own and inherited)

    Name (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Name
    SetName (me: mutable; Name: HAsciiString from TCollection);
	---Purpose: Set field Name

    Description (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Description
    SetDescription (me: mutable; Description: HAsciiString from TCollection);
	---Purpose: Set field Description

    RelatingPropertyDefinition (me) returns PropertyDefinition from StepRepr;
	---Purpose: Returns field RelatingPropertyDefinition
    SetRelatingPropertyDefinition (me: mutable; RelatingPropertyDefinition: PropertyDefinition from StepRepr);
	---Purpose: Set field RelatingPropertyDefinition

    RelatedPropertyDefinition (me) returns PropertyDefinition from StepRepr;
	---Purpose: Returns field RelatedPropertyDefinition
    SetRelatedPropertyDefinition (me: mutable; RelatedPropertyDefinition: PropertyDefinition from StepRepr);
	---Purpose: Set field RelatedPropertyDefinition

fields
    theName: HAsciiString from TCollection;
    theDescription: HAsciiString from TCollection;
    theRelatingPropertyDefinition: PropertyDefinition from StepRepr;
    theRelatedPropertyDefinition: PropertyDefinition from StepRepr;

end PropertyDefinitionRelationship;
