-- Created on: 1992-03-06
-- Created by: Isabelle GRIGNON
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred generic class ISurfaceTool from IntImp
       ( ImplicitSurface as any)
                                        
	---Purpose: Template class for a tool on an
	--          implicit surface.


uses Vec from gp


is

    Value(myclass; Is: ImplicitSurface;
          X, Y, Z: Real from Standard)
	  
    	---Purpose: Returns the value of the function.

    	returns Real from Standard;

    
    Gradient(myclass; Is: ImplicitSurface;
             X, Y, Z: Real from Standard ; V: out Vec from gp);
	     
    	---Purpose: Returns the gradient of the function.



    ValueAndGradient(myclass; Is: ImplicitSurface; 
                     X, Y, Z: Real from Standard;
                     Val: out Real from Standard; Grad: out Vec from gp);
		     
    	---Purpose: Returns the value and the gradient.


    Tolerance(myclass; Is: ImplicitSurface )
    
	---Purpose: returns the tolerance of the zero of the implicit function

    	returns Real from Standard; 

    
end ISurfaceTool;
