-- Created on: 1996-10-17
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class SurfaceExplorer from TopOpeBRepDS

uses

    DataStructure from TopOpeBRepDS,
    Surface from TopOpeBRepDS
    
is

    Create returns SurfaceExplorer from TopOpeBRepDS;
    Create(DS : DataStructure from TopOpeBRepDS;
           FindOnlyKeep : Boolean from Standard = Standard_True)
    returns SurfaceExplorer from TopOpeBRepDS;
    
    Init(me : in out;
    	 DS : DataStructure from TopOpeBRepDS;
         FindOnlyKeep : Boolean from Standard = Standard_True);
    
    More(me) returns Boolean  is static;
    Next(me : in out) is static;
    Surface(me) returns Surface from TopOpeBRepDS
    ---C++: return const &
    is static;

    IsSurface(me; I : Integer ) 
    returns Boolean  is static;
    IsSurfaceKeep(me; I : Integer ) returns Boolean  is static;
    Surface(me; I : Integer ) 
    returns Surface from TopOpeBRepDS
    ---C++: return const &
    is static;
    NbSurface(me : in out) returns Integer
    is static;

    Index(me) returns Integer 
    is static;

    Find(me : in out) is static private;
        
fields

    myIndex   : Integer ;
    myMax     : Integer ;
    myDS      : Address ; -- (TopOpeBRepDS_DataStructure*)
    myFound   : Boolean ;
    myEmpty   : Surface from TopOpeBRepDS;
    myFindKeep : Boolean;
    
end SurfaceExplorer from TopOpeBRepDS;
