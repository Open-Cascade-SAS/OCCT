-- File:	Scale2d.cdl
-- Created:	Wed Aug 26 14:35:24 1992
-- Author:	Remi GILET
--		<reg@topsn3>
---Copyright:	 Matra Datavision 1992

class MakeScale2d

from gce

    ---Purpose: This class implements an elementary construction algorithm for
    -- a scaling transformation in 2D space. The result is a gp_Trsf2d transformation.
    -- A MakeScale2d object provides a framework for:
    -- -   defining the construction of the transformation,
    -- -   implementing the construction algorithm, and
    -- -   consulting the result.

uses Pnt2d  from gp,
     Trsf2d from gp,
     Real   from Standard
     
is

Create(Point : Pnt2d from gp      ;
       Scale : Real  from Standard) returns MakeScale2d;
    --- Purpose:
    -- Constructs a scaling transformation with:
    -- -   Point as the center of the transformation, and
    -- -   Scale as the scale factor.
        
Value(me) returns Trsf2d from gp
    is static;
    ---C++: return const&
    ---Purpose: Returns the constructed transformation.

Operator(me) returns Trsf2d from gp
    is static;
    ---C++: return const&
    ---C++: alias "Standard_EXPORT operator gp_Trsf2d() const;"

fields

    TheScale2d : Trsf2d from gp;

end MakeScale2d;

