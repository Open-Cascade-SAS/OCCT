-- Created on: 1992-08-13
-- Created by: Remi LEQUETTE
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

generic class Interference from TopBas (TheSubShape as any;
    	    	    	    	    	TheShape    as any)

	---Purpose: An  Interference  is an   Intersection on a  Shape
	--          called  the Reference, it contains :
	--          
	--          * The  Intersection : The  SubShape describing the
	--          intersection. For example a Vertex.
	--          
	--          * The   Boundary : The  Shape  that  generated the
	--          intersection with the referrence.  For  example an
	--          Edge.
	--          
	--          *   The  Orientation  :  The  orientation  of  the
	--          Intersection relative to the Boundary.
	--          
	--          * The Transition : How the referrence  crosses the
	--          Boundary at the Intersection.
	--          
	--          * The  BoundaryTransition  : How the Referrence is
	--          on the boundary at the Intersection.
	--          
	--          *    Next : The    Next Interference  on  the same
	--          Reference. Used to make lists.


uses
    Orientation from TopAbs
    
is
   Create returns Interference;

   Create(Inters : TheSubShape;
   	  Bound  : TheShape;
	  Orient : Orientation from TopAbs;
	  Trans  : Orientation from TopAbs;
	  BTrans : Orientation from TopAbs) returns Interference; 
	   
   Intersection(me : in out; I : TheSubShape)
    	---C++: inline
   is static;
   
   Boundary(me : in out; B : TheShape)
    	---C++: inline
   is static;
   
   Orientation(me : in out; O : Orientation from TopAbs)
    	---C++: inline
   is static;
   
   Transition(me : in out; Tr : Orientation from TopAbs)
    	---C++: inline
   is static;
   
   BoundaryTransition(me : in out; BTr : Orientation from TopAbs)
    	---C++: inline
   is static;
   
   Intersection(me) returns TheSubShape
    	---C++: inline
	---C++: return const &
   is static;
   
   ChangeIntersection(me : in out) returns TheSubShape
    	---C++: inline
	---C++: return &
   is static;
   
   Boundary(me) returns TheShape
    	---C++: inline
	---C++: return const &
   is static;
   
   ChangeBoundary(me : in out) returns TheShape
    	---C++: inline
	---C++: return &
   is static;
   
   Orientation(me) returns Orientation from TopAbs
    	---C++: inline
   is static;
   
   Transition(me) returns Orientation from TopAbs
    	---C++: inline
   is static;
   
   BoundaryTransition(me) returns Orientation from TopAbs
    	---C++: inline
   is static;
   
fields
    myIntersection : TheSubShape;
    myBoundary     : TheShape;
    myOrientation  : Orientation from TopAbs;
    myTransition   : Orientation from TopAbs;
    myBTransition  : Orientation from TopAbs;

end Interference;
