-- Created on: 1999-03-10
-- Created by: data exchange team
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class AppliedSecurityClassificationAssignment from StepAP214 
inherits SecurityClassificationAssignment from StepBasic
	

uses
    	HArray1OfSecurityClassificationItem from StepAP214, 
	SecurityClassificationItem from StepAP214, 
	SecurityClassification from StepBasic


is
    	Create returns mutable AppliedSecurityClassificationAssignment;
	---Purpose: Returns a AppliedSecurityClassificationAssignment


	Init (me : mutable;
	      aAssignedSecurityClassification : mutable SecurityClassification from StepBasic) is redefined;

	Init (me : mutable;
	      aAssignedSecurityClassification : mutable SecurityClassification from StepBasic;
	      aItems : mutable HArray1OfSecurityClassificationItem from StepAP214) is virtual;

	-- Specific Methods for Field Data Access --

	SetItems(me : mutable; aItems : mutable HArray1OfSecurityClassificationItem from StepAP214);
	Items (me) returns mutable HArray1OfSecurityClassificationItem from StepAP214;
	ItemsValue (me; num : Integer) returns SecurityClassificationItem;
	---C++: return const &
	NbItems (me) returns Integer;
    

fields

    items :  HArray1OfSecurityClassificationItem from StepAP214;

end AppliedSecurityClassificationAssignment;
