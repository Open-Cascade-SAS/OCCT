-- Created on: 1999-10-11
-- Created by: Atelier CAS2000
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package  BRepFilletAPI 

uses    
    TColgp, 
    GeomAbs, 
    Geom,
    TopoDS,
    TopTools,
    BRepBuilderAPI, 
    ChFiDS,
    ChFi3d,
    ChFi2d, 
    TopOpeBRepBuild,
    Law 
     
is   

    -- 
    -- Local Operations
    --      
    deferred  class  LocalOperation  ;  ---  inherits  MakeShape  from BRepBuilderAPI
 
    class  MakeFillet    ;    ---  inherits  LocalOperation from BRepFilletAPI

    class  MakeChamfer   ;    ---  inherits  LocalOperation from BRepFilletAPI
     
    class  MakeFillet2d  ;    ---  inherits  inherits MakeShape from BRepBuilderAPI

end;
