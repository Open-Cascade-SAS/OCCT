-- Created on: 1998-07-14
-- Created by: data exchange team
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Curve from ShapeConstruct 

	---Purpose: Adjusts curve to have start and end points at the given
	--          points (currently works on lines and B-Splines only)

uses

    Pnt   from gp,
    Pnt2d from gp,
    Curve from Geom,
    Curve from Geom2d,
    BSplineCurve from Geom,
    BSplineCurve from Geom2d,
    HArray1OfReal from TColStd,
    Array1OfReal  from TColStd

is

    AdjustCurve (me; C3D: Curve from Geom;
    	    	     P1, P2: Pnt from gp;
    	    	     take1, take2: Boolean = Standard_True)
    returns Boolean;
    	---Purpose : Modifies a curve in order to make its bounds confused with
    	--           given points.
	--           Works only on lines and B-Splines, returns True in this case,
    	--           else returns False.           
	--           For line considers both bounding points, for B-Splines only
	--           specified.
    	--           
    	--  Warning : Does not check if curve should be reversed

    AdjustCurveSegment (me; C3D: Curve from Geom;
    	    	    	    P1, P2: Pnt from gp;
    	    	    	    U1, U2: Real)
    returns Boolean;
    	---Purpose : Modifies a curve in order to make its bounds confused with
    	--           given points.
	--           Works only on lines and B-Splines.
	--
	--           For lines works as previous method, B-Splines are segmented
	--           at the given values and then are adjusted to the points.

    AdjustCurve2d (me; C2D: Curve from Geom2d;
    	    	       P1, P2: Pnt2d from gp;
    	    	       take1, take2: Boolean = Standard_True)
    returns Boolean;
    	---Purpose : Modifies a curve in order to make its bounds confused with
    	--           given points.
	--           Works only on lines and B-Splines, returns True in this case,
    	--           else returns False.
    	--           
	--           For line considers both bounding points, for B-Splines only
	--           specified.
    	--           
    	--  Warning : Does not check if curve should be reversed

    ConvertToBSpline (me; C: Curve from Geom; first, last: Real; prec: Real) 
    returns BSplineCurve from Geom;
    	---Purpose: Converts a curve of any type (only part from first to last) 
        --          to bspline. The method of conversion depends on the type
	--          of original curve:
	--          BSpline -> C.Segment(first,last)
	--          Bezier and Line -> GeomConvert::CurveToBSplineCurve(C).Segment(first,last)
	--          Conic and Other -> Approx_Curve3d(C[first,last],prec,C1,9,1000)

    ConvertToBSpline (me; C: Curve from Geom2d; first, last: Real; prec: Real) 
    returns BSplineCurve from Geom2d;
    	---Purpose: Converts a curve of any type (only part from first to last) 
        --          to bspline. The method of conversion depends on the type
	--          of original curve:
	--          BSpline -> C.Segment(first,last)
	--          Bezier and Line -> GeomConvert::CurveToBSplineCurve(C).Segment(first,last)
	--          Conic and Other -> Approx_Curve2d(C[first,last],prec,C1,9,1000)
	
    FixKnots (myclass; knots: in out HArray1OfReal from TColStd) returns Boolean;
    FixKnots (myclass; knots: in out  Array1OfReal from TColStd) returns Boolean;
        ---Purpose: Fix bspline knots to ensure that there is enough
	--          gap between neighbouring values
	--          Returns True if something fixed (by shifting knot)


end Curve;
