-- Created on: 1994-02-03
-- Created by: Jean Marc LACHAUME
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Grid from Draw inherits Drawable3D from Draw

uses
    Display from Draw

is

    Create
     
    	---Purpose: Creates a grid.

	returns mutable Grid from Draw ;


    Steps (me : mutable; StepX, StepY, StepZ : Real from Standard)
    
    	---Purpose: Sets the steps along the X, Y & Z axis.

    	is static ;


    StepX (me)
    
    	---Purpose: Returns the step along the X axis.

	---C++: inline

    	returns Real from Standard
    	is static ;


    StepY (me)
    
    	---Purpose: Returns the step along the Y axis.

	---C++: inline

    	returns Real from Standard
    	is static ;


    StepZ (me)
    
    	---Purpose: Returns the step along the Z axis.

	---C++: inline

    	returns Real from Standard
    	is static ;


    IsActive (me)

    	---Purpose: Returns if the grid is active or not.

	---C++: inline

    	returns Boolean from Standard
	is static ;


    DrawOn (me; Out : in out Display from Draw)

    	---Purpose: Displays the grid.

    	is static ;


fields

  myStepX    : Real    from Standard ;
  myStepY    : Real    from Standard ;
  myStepZ    : Real    from Standard ;
  myIsActive : Boolean from Standard ;

end Grid ;
