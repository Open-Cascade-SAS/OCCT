-- Created on: 2000-05-10
-- Created by: Andrey BETENEV
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1

class IdentificationAssignment from StepBasic
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity IdentificationAssignment

uses
    HAsciiString from TCollection,
    IdentificationRole from StepBasic

is
    Create returns IdentificationAssignment from StepBasic;
	---Purpose: Empty constructor

    Init (me: mutable; aAssignedId: HAsciiString from TCollection;
                       aRole: IdentificationRole from StepBasic);
	---Purpose: Initialize all fields (own and inherited)

    AssignedId (me) returns HAsciiString from TCollection;
	---Purpose: Returns field AssignedId
    SetAssignedId (me: mutable; AssignedId: HAsciiString from TCollection);
	---Purpose: Set field AssignedId

    Role (me) returns IdentificationRole from StepBasic;
	---Purpose: Returns field Role
    SetRole (me: mutable; Role: IdentificationRole from StepBasic);
	---Purpose: Set field Role

fields
    theAssignedId: HAsciiString from TCollection;
    theRole: IdentificationRole from StepBasic;

end IdentificationAssignment;
