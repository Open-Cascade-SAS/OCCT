-- Created on: 1997-04-09
-- Created by: VAUTHIER Jean-Claude
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Real from PDataStd inherits Attribute from PDF

	---Purpose: 

uses Real from Standard

is

    Create returns mutable Real from PDataStd;

    
    Create (Value     : Real from Standard;
            Dimension : Integer from Standard)
    returns mutable Real from PDataStd;
    
    Get (me) returns Real from Standard;

    Set (me : mutable; V : Real from Standard);
    
    SetDimension (me : mutable; DIM : Integer from Standard);
    
    GetDimension (me)
    returns Integer from Standard;

fields

    myValue     : Real    from Standard;
    myDimension : Integer from Standard;

end Real;
