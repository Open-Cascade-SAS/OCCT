-- Created on: 1993-07-22
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class MakeOneAxis from BRepPrimAPI inherits MakeShape from BRepBuilderAPI

	---Purpose: The abstract class MakeOneAxis is the root class of
    	-- algorithms used to construct rotational primitives.

uses
    Address from Standard,
    Face    from TopoDS,
    Shell   from TopoDS,
    Solid   from TopoDS

raises
    NotDone     from StdFail

is
    OneAxis(me : in out) returns Address from Standard
	---Purpose: The inherited commands should provide the algorithm.
	--          Returned as a pointer.
	---Level: Public
    is deferred;
    
    Build(me : in out)
	---Purpose: Stores the solid in myShape.
	---Level: Public
    is redefined;

    Face(me : in out) 
	---Purpose: Returns the lateral face of the rotational primitive.
	--          
	---C++: return const &
	---C++: alias "Standard_EXPORT operator TopoDS_Face();" 
	---Level: Public
    returns Face from TopoDS
    is static;

    Shell(me : in out) 
	---Purpose: Returns the constructed rotational primitive as a shell.
    	---C++: return const &
	---C++: alias "Standard_EXPORT operator TopoDS_Shell();" 
    returns Shell from TopoDS
    is static;

    Solid(me : in out) 
	---Purpose: Returns the constructed rotational primitive as a solid.
	---C++: return const &
	---C++: alias "Standard_EXPORT operator TopoDS_Solid();" 
    returns Solid from TopoDS 
    is static;


end MakeOneAxis;
