-- Created on: 1999-02-11
-- Created by: Pavel DURANDIN
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Counter from STEPSelections

	---Purpose: 

uses
   
    Graph from Interface,
    MapOfTransient from TColStd,
    ConnectedFaceSet from StepShape,
    CompositeCurve from StepGeom
  
is
    Create returns Counter from STEPSelections;
    
    Count(me: in out;graph: Graph from Interface;
    	            start: Transient);
	  
    Clear(me: in out);
    
    NbInstancesOfFaces(me)  returns Integer;
    	---C++: inline
    	---Purpose:
    
    POP(me)  returns Integer;
    	---C++: inline
    	---Purpose:
    
    POP2(me)  returns Integer
    	---C++: inline
	;
    	---Purpose:
    
    NbInstancesOfShells(me) returns Integer;
    	---C++: inline
    	---Purpose:
    
    NbInstancesOfSolids(me) returns Integer;
    	---C++: inline
    	---Purpose:
    
    NbInstancesOfEdges(me) returns Integer;
    	---C++: inline
	---Purpose:
    
    NbInstancesOfWires(me) returns Integer;
    	---C++: inline
	---Purpose:
	
    NbSourceFaces(me)  returns Integer;
    	---C++: inline
    	---Purpose:
    
    NbSourceShells(me) returns Integer;
    	---C++: inline
    	---Purpose:
    
    NbSourceSolids(me) returns Integer;
    	---C++: inline
    	---Purpose:
	
    NbSourceEdges(me) returns Integer;
    	---C++: inline
	---Purpose:
	
    NbSourceWires(me) returns Integer;
    	---C++: inline
	---Purpose:
	
   AddShell(me: in out; cfs: ConnectedFaceSet from StepShape) is private;
   
   AddCompositeCurve(me: in out; ccurve: CompositeCurve from StepGeom) is private;

fields

    myNbFaces : Integer;
    myNbShells: Integer;
    myNbSolids: Integer;
    myNbEdges : Integer;
    myNbWires : Integer;
    
    myMapOfFaces : MapOfTransient from TColStd;
    myMapOfShells: MapOfTransient from TColStd;
    myMapOfSolids: MapOfTransient from TColStd;  
    myMapOfEdges : MapOfTransient from TColStd;
    myMapOfWires : MapOfTransient from TColStd;

end Counter;
