-- Created on: 1995-03-16
-- Created by: Christian CAILLET
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Functions  from XSDRAW

    ---Purpose : Defines additionnal commands for XSDRAW to :
    --           - control of initialisation (xinit, xnorm, newmodel)
    --           - analyse of the result of a transfer (recorded in a
    --             TransientProcess for Read, FinderProcess for Write) :
    --             statistics, various lists (roots,complete,abnormal), what
    --             about one specific entity, producing a model with the
    --             abnormal result
    --             
    --           This appendix of XSDRAW is compiled separately to distinguish
    --           basic features from user callable forms

uses CString

is

    Init (myclass);
    ---Purpose : Defines and loads all basic functions for XSDRAW (as ActFunc)

end Functions;
