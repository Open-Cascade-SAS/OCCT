-- Created on: 1999-08-11
-- Created by: Roman LYGIN
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class TransferResultInfo from TransferBRep inherits TShared from MMgt 

    ---Purpose: Data structure for storing information on transfer result.
    --          At the moment it dispatches information for the following types:
    --          - result,
    --          - result + warning(s),
    --          - result + fail(s),
    --          - result + warning(s) + fail(s)
    --          - no result,
    --          - no result + warning(s),
    --          - no result + fail(s),
    --          - no result + warning(s) + fail(s),

is

    Create returns TransferResultInfo from TransferBRep;
    	---Purpose: Creates object with all fields nullified.
	
    Clear (me: mutable);
    	---Purpose: Resets all the fields.
	
    Result (me: mutable) returns Integer;
    	---C++: inline
    	---C++: return &
	
    ResultWarning (me: mutable) returns Integer;
    	---C++: inline
    	---C++: return &
	
    ResultFail (me: mutable) returns Integer;
    	---C++: inline
    	---C++: return &
	
    ResultWarningFail (me: mutable) returns Integer;
    	---C++: inline
    	---C++: return &
	
    NoResult (me: mutable) returns Integer;
    	---C++: inline
    	---C++: return &
	
    NoResultWarning (me: mutable) returns Integer;
    	---C++: inline
    	---C++: return &
	
    NoResultFail (me: mutable) returns Integer;
    	---C++: inline
    	---C++: return &
	
    NoResultWarningFail (me: mutable) returns Integer;
    	---C++: inline
    	---C++: return &
	
fields

    myR,  myRW,  myRF,  myRWF,
    myNR, myNRW, myNRF, myNRWF: Integer;
    
end TransferResultInfo;
