-- Created on: 1992-02-19
-- Created by: Jean Pierre TIRAULT
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

generic class HSingleList from PCollection (Item as Storable) 
inherits PManaged 

raises
    NoSuchObject from Standard

is

	---Purpose: Definition of a single linked list.

	Create returns mutable HSingleList;
		---Creation of an empty list.

	IsEmpty(me) returns Boolean from Standard;
                ---Level: Public
		---Purpose: Returns True if the list contains no element.


	Construct(me; T : Item) returns mutable 
		HSingleList;
                ---Level: Public
		---Purpose: add T at the begining of me
		---Example: before
		--   me = (A B C) 
                -- after
		--   me = (A B C)
		-- returns 
		--   (T A B C)

	Value(me) returns any Item
                raises NoSuchObject from Standard;
                ---Level: Public
		---Purpose: Returns the value of the first node of me.
		-- Raises an exception if me is empty.
		---Example: before
		--   me = (A B C) 
                -- after
		--   me = (A B C)
		-- returns 
		--   A

	Tail(me) returns any HSingleList
                raises NoSuchObject from Standard;
                ---Level: Public
		---Purpose: End of the list me.
		-- Raises an exception if me is empty.
		---Example: before
		--   me = (A B C) 
                -- after
		--   me = (A B C)
		-- returns 
		--   (B C)

	SwapTail(me : mutable; WithList : in out any HSingleList)
	   	raises NoSuchObject from Standard;
                ---Level: Public
		---Purpose: Exchanges the end of <me> with the list WithList.
		-- Raises an exception if me is empty.
		---Example: before
		--   me = (A B C)
		--   WithList = (D E)
		-- after
		--   me = (A D E)
		--   WithList = (B C)
		
	SetValue(me : mutable; T : Item)
                raises NoSuchObject from Standard ;
                ---Level: Public
		---Purpose: Changes the value of the first node of me.
		-- Raises an exception if me is empty.
		---Example: before
		--   me = (A B C) 
                -- after
		--   me = (T B C)

	ChangeForwardPointer(me : mutable; ForwardPointer : HSingleList);
                ---Level: Public
		---Purpose: Modification of the node link.

fields 
           Data : 	Item;
           Next : 	HSingleList;

end HSingleList;
