-- Created on: 1992-10-13
-- Created by: Laurent BUCHARD
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.





generic class ProjPCurGen from IntCurve (
    TheCurve         as any;
    TheCurveTool     as any) -- as CurveTool from IntCurve(TheCurve)

    ---Purpose: this class provide a tool which computes the parameter
    --          of a point near a parametric curve.

    ---Level: Internal

uses Pnt2d     from gp,
     Vec2d     from gp,
     POnCurv2d from Extrema
     
     

    class TheCurveLocator instantiates CurveLocator from Extrema (
    	TheCurve,
	TheCurveTool,
	TheCurve,
	TheCurveTool,
	POnCurv2d       from Extrema,
	Pnt2d           from gp);
	
    class TheLocateExtPC instantiates GenLocateExtPC from Extrema (
	TheCurve,
	TheCurveTool,
	POnCurv2d      from Extrema,
	Pnt2d          from gp,
	Vec2d          from gp);



is
		 
    FindParameter(myclass; C:   TheCurve;
    	    	           Pnt: Pnt2d  from gp;
			   Tol: Real   from Standard)
			   
	--- Purpose: Returns the parameter V of the point on the 
	--           parametric curve corresponding to the Point Pnt.
	--           The Correspondance between Pnt and the point P(V) 
	--           on the parametric curve must be coherent with the 
	--           way of determination of the signed distance 
	--           between a point and the implicit curve.
	--           Tol is the tolerance on the distance between a point
	--           and the parametrised curve.
	--           In that case, no bounds are given. The research of
	--           the rigth parameter has to be made on the natural
	--           parametric domain of the curve.
			   
    	returns Real from Standard;

	
    FindParameter(myclass; C:   TheCurve;
    	    	           Pnt: Pnt2d  from gp;
			   LowParameter,HighParameter,Tol: Real from Standard)
			   
	--- Purpose: Returns the parameter V of the point on the 
	--           parametric curve corresponding to the Point Pnt.
	--           The Correspondance between Pnt and the point P(V) 
	--           on the parametric curve must be coherent with the 
	--           way of determination of the signed distance 
	--           between a point and the implicit curve.
	--           Tol is the tolerance on the distance between a point
	--           and the parametrised curve.
	--           LowParameter and HighParameter give the 
	--           boundaries of the interval in wich the parameter 
	--           certainly lies. These parameters are given to
	--           implement a more efficient algoritm. So, it is not
	--           necessary to check that the returned value verifies 
	--                LowParameter <= Value <= HighParameter.
			   
    	returns Real from Standard;
	
end ProjPCurGen;



