-- Created on: 1993-06-23
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Surface from TopOpeBRepDS

    ---Purpose: A Geom poimt and a tolerance.

uses

    Surface from Geom

is

    Create returns Surface from TopOpeBRepDS; 
    
    Create(P : Surface from Geom; T : Real from Standard)
    returns Surface from TopOpeBRepDS; 
     
--modified by NIZNHY-PKV Tue Oct 30 09:27:32 2001  f    
    Create  (Other :Surface from TopOpeBRepDS) 
    	returns Surface from TopOpeBRepDS; 
	 
    Assign(me :out;  
    	    Other: Surface from TopOpeBRepDS);  
    ---C++: alias operator=
--modified by NIZNHY-PKV Tue Oct 30 09:27:25 2001  t     

    Surface(me) returns Surface from Geom
	---C++: return const &
    is static;
    
    Tolerance(me) returns Real from Standard
    is static;

    Tolerance(me : in out; tol : Real)
    ---Purpose: Update the tolerance
    is static;
	
    Keep(me) returns Boolean from Standard
    is static;
    ChangeKeep(me : in out; B : Boolean from Standard)
    is static;

fields

    mySurface   : Surface from Geom;
    myTolerance : Real from Standard;
    myKeep      : Boolean from Standard;

end Surface from TopOpeBRepDS;
