-- Created on: 1995-09-01
-- Created by: Bruno DUMORTIER
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class OffsetAncestors from BRepFill 

	---Purpose: this class is used to find the generating shapes
	--          of an OffsetWire.

uses
    OffsetWire          from BRepFill,
    Shape               from TopoDS,
    Edge                from TopoDS,	
    DataMapOfShapeShape from TopTools
    
raises
    NotDone from StdFail
    
is
    Create returns OffsetAncestors from BRepFill;
    
    Create ( Paral : in out OffsetWire from BRepFill)
    returns OffsetAncestors from BRepFill;
    
    Perform ( me : in out; Paral : in out OffsetWire from BRepFill)
    is static;
    
    IsDone( me)
    returns Boolean from Standard
    is static;

    HasAncestor (me; S1 : Edge from TopoDS)	    
    returns Boolean from Standard
    is static;

    Ancestor    (me ; S1 : Edge from TopoDS)
	---Purpose: may return a Null Shape if S1 is not a subShape
	--          of <Paral>;
	---C++: return const &
    returns Shape from TopoDS
    raises
    	NotDone from StdFail
	---Purpose: if Perform is not done.
    is static;
    
fields

    myIsPerform : Boolean             from Standard;
    myMap       : DataMapOfShapeShape from TopTools;
    
end OffsetAncestors;
