-- Created on: 1996-01-09
-- Created by: Laurent PAINNOT
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

private class FuncExtSS from Extrema

 inherits FunctionSetWithDerivatives from math
    ---Purpose: Function to find extrema of the 
    --          distance between two surfaces.

uses    POnSurf           from Extrema,
	SequenceOfPOnSurf from Extrema,
	SequenceOfReal    from TColStd,
	Pnt               from gp,
	Vector            from math,
	Matrix            from math,
	Surface           from Adaptor3d,
    	SurfacePtr        from Adaptor3d

raises  OutOfRange from Standard

is
    Create returns FuncExtSS;

    Create (S1, S2: Surface from Adaptor3d) returns FuncExtSS;
    	---Purpose:

    Initialize(me: in out; S1, S2: Surface from Adaptor3d)
    	---Purpose: sets the field mysurf of the function.
    is static;
    
    ------------------------------------------------------------
    -- In all next methods, an exception is raised if the fields 
    -- were not initialized.

    NbVariables (me) returns Integer;

    NbEquations (me) returns Integer;

    Value (me: in out; UV: Vector; F: out Vector) returns Boolean;
    	---Purpose: Calculate Fi(U,V).

    Derivatives (me: in out; UV: Vector; DF: out Matrix)
    	returns Boolean;
    	---Purpose: Calculate Fi'(U,V).

    Values (me: in out; UV: Vector; F: out Vector; DF: out Matrix)
    	returns Boolean;
    	---Purpose: Calculate Fi(U,V) and Fi'(U,V).

    GetStateNumber (me: in out) returns Integer
    	---Purpose: Save the found extremum.
    	is redefined;

    NbExt (me) returns Integer;
    	---Purpose: Return the number of found extrema.

    SquareDistance (me; N: Integer) returns Real
    	---Purpose: Return the value of the Nth distance.
    	raises  OutOfRange;
	    	-- if N < 1 or N > NbExt(me).

    PointOnS1 (me; N: Integer) returns POnSurf
        ---C++: return const &
    	---Purpose: Return the Nth extremum on S1.
    	raises  OutOfRange;
	    	-- if N < 1 or N > NbExt(me).

    PointOnS2 (me; N: Integer) returns POnSurf
        ---C++: return const &
    	---Purpose: Renvoie le Nieme extremum sur S2.
    	raises  OutOfRange;
	    	-- si N < 1 ou N > NbExt(me).

    Bidon(me) returns SurfacePtr from Adaptor3d
    is static private;


fields
    myS1   : SurfacePtr from Adaptor3d;
    myS2   : SurfacePtr from Adaptor3d;
    
    myP1   : Pnt from gp;
    myP2   : Pnt from gp;

    myU1    : Real;          -- current value of U on S1
    myV1    : Real;          -- current value of V on S1
    myU2    : Real;          -- current value of U on S2
    myV2    : Real;          -- current value of V on S2

    mySqDist:  SequenceOfReal    from TColStd;
    myPoint1: SequenceOfPOnSurf from Extrema;
    myPoint2: SequenceOfPOnSurf from Extrema;
    
    myS1init: Boolean;
    myS2init: Boolean;

end FuncExtSS;
