-- Created by: Peter KURNEV
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class EdgeSet from BOPTools 


uses 
    Shape from TopoDS, 
    Edge from TopoDS,
    ShapeEnum from TopAbs,  
    BaseAllocator from BOPCol, 
    MapOfShape from BOPCol, 
    ListOfShape from BOPCol 
    
--raises

is 
    Create 
    	returns EdgeSet from BOPTools;  
    ---C++: alias "virtual ~BOPTools_EdgeSet();"  
    ---C++: inline 
     
    Create (theAllocator: BaseAllocator from BOPCol)
    	returns EdgeSet from BOPTools; 
    ---C++: inline   
     
    SetShape(me:out; 
    	    theS:Shape from TopoDS); 
    ---C++: inline  
     
    Shape(me) 
    	 returns Shape from TopoDS; 
    ---C++: return const & 
    ---C++: inline  
    
    AddEdge(me:out; 
    	    theEdge:Edge from TopoDS); 
    ---C++: inline 

    AddEdges(me:out; 
    	    theLS:ListOfShape from BOPCol);  

    AddEdges(me:out; 
    	    theFace:Shape from TopoDS); 
    ---C++: inline 
     
    Clear(me:out);
    ---C++: inline 
    
    Get(me; 
	    theLS:out ListOfShape from BOPCol);     
    ---C++: inline 
    
    Contains(me; 
	    theSet:EdgeSet from BOPTools) 
    	returns Boolean from Standard; 
    ---C++: inline
    
     
fields  
    myShape  : Shape from TopoDS is protected;   
    myMap    : MapOfShape from BOPCol is protected;   
    myEdges : ListOfShape from BOPCol is protected;   
	    
end EdgeSet; 
