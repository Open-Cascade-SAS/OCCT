-- Created on: 1995-03-09
-- Created by: Laurent PAINNOT
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




deferred class GCurve from BRep inherits CurveRepresentation from BRep

	---Purpose: Root   class    for    the    geometric     curves
	--          representation. Contains a range.

uses

    Location from TopLoc,
    Pnt      from gp

is

    Initialize(L : Location from TopLoc; First, Last : Real);

    SetRange(me : mutable; First, Last : Real)
	---C++: inline
    is static;
    
    Range(me; First, Last : out Real)
	---C++: inline
    is static;
    
    First(me) returns Real
	---C++: inline
    is static;

    Last(me) returns Real
	---C++: inline
    is static;

    First(me : mutable; F : Real)
	---C++: inline
    is static;

    Last(me : mutable; L : Real)
	---C++: inline
    is static;


    D0(me; U : Real; P : out Pnt from gp)
	---Purpose: Computes the point at parameter U.
    is deferred;
    

    Update(me : mutable)
	---Purpose: Recomputes any derived data after a modification.
	--          This is called when the range is modified.
    is virtual;

fields
    myFirst    : Real;
    myLast     : Real;

end GCurve;
