-- Created on: 2001-07-25
-- Created by: Julia DOROVSKIKH
-- Copyright (c) 2001-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class DocumentRetrievalDriver from XmlDrivers inherits DocumentRetrievalDriver from XmlLDrivers

uses

    ADriverTable		from XmlMDF, 
    ADriver                     from XmlMDF, 
    Element                     from XmlObjMgt,
    MessageDriver               from CDM

is
    Create returns mutable DocumentRetrievalDriver from XmlDrivers;
    -- Constructor

    AttributeDrivers	(me : mutable; theMsgDriver: MessageDriver from CDM)
	returns ADriverTable from XmlMDF
	is redefined virtual; 
	 
    ReadShapeSection (me:mutable; thePDoc  :  Element from XmlObjMgt; 
                                  theMsgDriver : MessageDriver from CDM) 
        returns ADriver from XmlMDF
        is redefined virtual; 
	 
    ShapeSetCleaning(me:mutable; theDriver : ADriver from XmlMDF) 
        is redefined virtual;
	
    PropagateDocumentVersion(me:mutable; theDocVersion : Integer from Standard) 
        is redefined virtual;  
	 
end DocumentRetrievalDriver;
