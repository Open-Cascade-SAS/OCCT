-- File:        BRepMesh_Triangle.cdl
-- Created:     Wed Sep 22 18:11:52 1993
-- Author:      Didier PIFFAULT
--              <dpf@zerox>
---Copyright:    Matra Datavision 1993


class Triangle from BRepMesh 

  ---Purpose: 

uses    Boolean from Standard,
        Integer from Standard,
        DegreeOfFreedom from BRepMesh



is        Create  returns Triangle from BRepMesh;


          Create         (e1, e2, e3 : Integer from Standard;
                          o1, o2, o3 : Boolean from Standard;
                          canMove : DegreeOfFreedom from BRepMesh)
            returns Triangle from BRepMesh;


          Initialize     (me : in out;
                          e1, e2, e3 : Integer from Standard;
                          o1, o2, o3 : Boolean from Standard;
                          canMove : DegreeOfFreedom from BRepMesh)
            is static;


          Edges          (me;
                          e1, e2, e3 : out Integer from Standard;
                          o1, o2, o3 : out Boolean from Standard)
            is static;


          Movability     (me)
            ---C++: inline
            returns DegreeOfFreedom from BRepMesh
            is static;


          SetMovability  (me   : in out;
                          Move : DegreeOfFreedom from BRepMesh)
            is static;


          HashCode       (me;
                          Upper : Integer from Standard)
            returns Integer from Standard
            ---C++: function call
            is static;


          IsEqual        (me; Other : Triangle from BRepMesh)
            returns Boolean from Standard
            ---C++: alias operator ==
            is static;


        fields  Edge1        : Integer from Standard;
                Orientation1 : Boolean from Standard;
                Edge2        : Integer from Standard;
                Orientation2 : Boolean from Standard;
                Edge3        : Integer from Standard;
                Orientation3 : Boolean from Standard;
                myMovability : DegreeOfFreedom from BRepMesh;

end Triangle;
