-- Created on: 1994-04-18
-- Created by: Modelistation
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Text2D from Draw inherits Drawable2D from Draw

	---Purpose: 

uses Pnt2d from gp,
    Color from Draw,
    Display from Draw,
    AsciiString from TCollection

is

    Create(p : Pnt2d; T : CString; col : Color)
    returns mutable Text2D from Draw;
    
    Create(p : Pnt2d; T : CString; col : Color;
    	   moveX : Integer; moveY : Integer)
    returns mutable Text2D from Draw;
    
    SetPnt2d(me : mutable; p : Pnt2d);

    DrawOn(me; dis : in out Display);

fields

    myPoint : Pnt2d        from gp;
    myColor : Color        from Draw;
    myText  : AsciiString  from TCollection;
    mymoveX : Integer      from Standard;
    mymoveY : Integer      from Standard;
    
end Text2D;
