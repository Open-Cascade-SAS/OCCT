-- File:	RWStepRepr_RWMaterialPropertyRepresentation.cdl
-- Created:	Thu Dec 12 17:15:59 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWMaterialPropertyRepresentation from RWStepRepr

    ---Purpose: Read & Write tool for MaterialPropertyRepresentation

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    MaterialPropertyRepresentation from StepRepr

is
    Create returns RWMaterialPropertyRepresentation from RWStepRepr;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : MaterialPropertyRepresentation from StepRepr);
	---Purpose: Reads MaterialPropertyRepresentation

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: MaterialPropertyRepresentation from StepRepr);
	---Purpose: Writes MaterialPropertyRepresentation

    Share (me; ent : MaterialPropertyRepresentation from StepRepr;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWMaterialPropertyRepresentation;
