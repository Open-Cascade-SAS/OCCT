-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class SurfaceStyleElementSelect from StepVisual inherits SelectType from StepData

	-- <SurfaceStyleElementSelect> is an EXPRESS Select Type construct translation.
	-- it gathers : SurfaceStyleFillArea, SurfaceStyleBoundary, SurfaceStyleSilhouette, SurfaceStyleSegmentationCurve, SurfaceStyleControlGrid, SurfaceStyleParameterLine
	-- Rev4 : only remain SurfaceStyleFillArea, SurfaceStyleBoundary, SurfaceStyleParameterLine

uses

	SurfaceStyleFillArea,
	SurfaceStyleBoundary,
--	SurfaceStyleSilhouette,
--	SurfaceStyleSegmentationCurve,
--	SurfaceStyleControlGrid,
	SurfaceStyleParameterLine
is

	Create returns SurfaceStyleElementSelect;
	---Purpose : Returns a SurfaceStyleElementSelect SelectType

	CaseNum (me; ent : Transient) returns Integer;
	---Purpose: Recognizes a SurfaceStyleElementSelect Kind Entity that is :
	--        1 -> SurfaceStyleFillArea
	--        2 -> SurfaceStyleBoundary
	--        3 -> SurfaceStyleParameterLine
	--        4 -> SurfaceStyleSilhouette
	--        5 -> SurfaceStyleSegmentationCurve
	--        6 -> SurfaceStyleControlGrid
	--        0 else

	SurfaceStyleFillArea (me) returns any SurfaceStyleFillArea;
	---Purpose : returns Value as a SurfaceStyleFillArea (Null if another type)

	SurfaceStyleBoundary (me) returns any SurfaceStyleBoundary;
	---Purpose : returns Value as a SurfaceStyleBoundary (Null if another type)

	SurfaceStyleParameterLine (me) returns any SurfaceStyleParameterLine;
	---Purpose : returns Value as a SurfaceStyleParameterLine (Null if another type)


end SurfaceStyleElementSelect;

