-- Created on: 1997-07-28
-- Created by: Pierre CHALAMET
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Texture1Dmanual from Graphic3d

inherits Texture1D from Graphic3d

---Purpose: This class provides the implementation of a manual 1D texture.
-- you MUST provides texture coordinates on your facets if you want to see your texture. 

uses

  NameOfTexture1D from Graphic3d,
  AsciiString     from TCollection,
  PixMap_Handle   from Image

is

  Create (theFileName : AsciiString from TCollection) returns mutable Texture1Dmanual from Graphic3d;
  ---Purpose: Creates a texture from the file FileName.

  Create (theNOT : NameOfTexture1D from Graphic3d) returns mutable Texture1Dmanual from Graphic3d;
  ---Purpose: Create a texture from a predefined texture name set.

  Create (thePixMap : PixMap_Handle from Image) returns mutable Texture1Dmanual from Graphic3d;
  ---Purpose: Creates a texture from the pixmap.

end Texture1Dmanual;
