-- File:	StepFEA_NodeGroup.cdl
-- Created:	Thu Dec 12 17:51:06 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class NodeGroup from StepFEA
inherits FeaGroup from StepFEA

    ---Purpose: Representation of STEP entity NodeGroup

uses
    HAsciiString from TCollection,
    FeaModel from StepFEA,
    HArray1OfNodeRepresentation from StepFEA

is
    Create returns NodeGroup from StepFEA;
	---Purpose: Empty constructor

    Init (me: mutable; aGroup_Name: HAsciiString from TCollection;
                       aGroup_Description: HAsciiString from TCollection;
                       aFeaGroup_ModelRef: FeaModel from StepFEA;
                       aNodes: HArray1OfNodeRepresentation from StepFEA);
	---Purpose: Initialize all fields (own and inherited)

    Nodes (me) returns HArray1OfNodeRepresentation from StepFEA;
	---Purpose: Returns field Nodes
    SetNodes (me: mutable; Nodes: HArray1OfNodeRepresentation from StepFEA);
	---Purpose: Set field Nodes

fields
    theNodes: HArray1OfNodeRepresentation from StepFEA;

end NodeGroup;
