-- Created on: 1993-09-07
-- Created by: Bruno DUMORTIER
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ComputeApprox from ProjLib 


uses
     HCurve       from Adaptor3d,
     HSurface     from Adaptor3d,
     BSplineCurve from Geom2d,
     BezierCurve  from Geom2d
is

    Create(C   : HCurve   from Adaptor3d ; 
           S   : HSurface from Adaptor3d;
    	   Tol : Real     from Standard) 
    	---Purpose: <Tol>    is   the   tolerance   with  which    the
    	--          approximation is performed.
    returns ComputeApprox from ProjLib;
    
    BSpline(me) returns BSplineCurve from Geom2d ;

    Bezier(me)  returns BezierCurve  from Geom2d ;
    
    Tolerance(me) returns Real from Standard;
    	---Purpose: returns the reached Tolerance.
    
fields

    myTolerance : Real         from Standard;    
    myBSpline   : BSplineCurve from Geom2d ;
    myBezier    : BezierCurve  from Geom2d ;

end ComputeApprox;
