-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Reducer from TopOpeBRepDS 

---Purpose: reduce interferences of a data structure (HDS)
--          used in topological operations.

uses

    DataMapOfShapeListOfShapeOn1State from TopOpeBRepDS,
    HDataStructure from TopOpeBRepDS

is

    Create(HDS:HDataStructure from TopOpeBRepDS) returns Reducer from TopOpeBRepDS;
    ProcessFaceInterferences(me:out;M:DataMapOfShapeListOfShapeOn1State);
    ProcessEdgeInterferences(me:out);

fields

    myHDS : HDataStructure from TopOpeBRepDS;
    
end Reducer from TopOpeBRepDS;
