-- File:	StepBasic_ExternalSource.cdl
-- Created:	Wed May 10 15:09:06 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class ExternalSource from StepBasic
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity ExternalSource

uses
    SourceItem from StepBasic

is
    Create returns ExternalSource from StepBasic;
	---Purpose: Empty constructor

    Init (me: mutable; aSourceId: SourceItem from StepBasic);
	---Purpose: Initialize all fields (own and inherited)

    SourceId (me) returns SourceItem from StepBasic;
	---Purpose: Returns field SourceId
    SetSourceId (me: mutable; SourceId: SourceItem from StepBasic);
	---Purpose: Set field SourceId

fields
    theSourceId: SourceItem from StepBasic;

end ExternalSource;
