-- Created on: 1995-01-27
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package GeomInt

	---Purpose: Provides intersections on between two surfaces of Geom.
	--          The result are curves from Geom.


uses StdFail,
     TCollection,
     TColStd,
     TopAbs,
     
     gp,
     Geom,
     Geom2d,
     TColGeom,
     TColGeom2d,     
     Adaptor3d,
     GeomAdaptor,

     IntSurf,
     IntPatch,
     ApproxInt

is

    class IntSS;

    class LineConstructor;

    class LineTool;

    class WLApprox instantiates Approx from ApproxInt
    	(HSurface     from Adaptor3d,
	 HSurfaceTool from Adaptor3d,
	 Quadric      from IntSurf,
	 QuadricTool  from IntSurf,
	 WLine        from IntPatch);

    private class ParameterAndOrientation;

    private class SequenceOfParameterAndOrientation instantiates
    	Sequence from TCollection(ParameterAndOrientation);

end GeomInt;
