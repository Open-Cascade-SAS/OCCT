-- Created on: 1997-02-19
-- Created by: Alexander BRIVIN
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


---Purpose: WFDeflectionShape -   computes    the    wireframe
--          presentation of compound set  of faces,  edges and
--          vertices by displaying a  given number of U and/or
--          V isoparametric  curves,   converts this  one into  VRML
--          objects and writes (adds) them into anOStream.
--          All requested properties of the representation are
--          specify in aDrawer. 
--          This kind of the presentation  is  converted  into
--          IndexedLineSet and PointSet ( VRML ).

--          The isoparametric curves are drawn  with respect to
--          a given maximal chordial deviation.

class WFDeflectionShape from VrmlConverter 

uses
 
    Shape            from TopoDS,
    Length           from Quantity,
    Drawer           from VrmlConverter

is
 
    Add(myclass; anOStream: in out OStream from Standard;
    	    	 aShape       : Shape        from TopoDS;
                 aDrawer      : Drawer       from VrmlConverter);
	
	 
end WFDeflectionShape;
