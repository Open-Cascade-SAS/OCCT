-- Created on: 1993-02-09
-- Created by: Mireille MERCIEN
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package PCollection

uses 
    Standard,
    DBC,
    MMgt,
    PMMgt,
    TCollection
 
is
          
        enumeration AccessMode is
    	    Read,
	    Update
        end AccessMode;

    
        generic class HArray1, FieldOfHArray1 ;   

        generic class HArray2, FieldOfHArray2 ;   

	generic class HSequence,SeqNode,SeqExplorer;

		---Purpose: Generic sequence of elements
		-- indexed by an integer in the range 1..N.

	
        class HAsciiString;

	class HExtendedString;
	
	
end PCollection;


