-- Created on: 1995-03-09
-- Created by: Laurent PAINNOT
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Polygon3D from BRep inherits CurveRepresentation from BRep

	---Purpose: 

uses
    Polygon3D           from Poly,
    CurveRepresentation from BRep,
    Location            from TopLoc

raises DomainError from Standard

is

    Create(P: Polygon3D from Poly;
    	   L: Location  from TopLoc) 
    	---Purpose:

    returns Polygon3D from BRep;
    
    
    IsPolygon3D(me) returns Boolean
    	---Purpose: Returns True.
    is redefined;
    
    Polygon3D(me) returns any Polygon3D from Poly
    	---C++: return const&
    is redefined;
    
    Polygon3D(me: mutable; P: Polygon3D from Poly)
    raises
    	DomainError from Standard
    is redefined;

    Copy(me) returns CurveRepresentation from BRep;
	---Purpose: Return a copy of this representation.


fields

myPolygon3D: Polygon3D from Poly;


end Polygon3D;
