-- Created on: 1992-10-28
-- Created by: Christian CAILLET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class TransferIterator  from Transfer

    ---Purpose : Defines an Iterator on the result of a Transfer
    --           Available for Normal Results or not (Erroneous Transfer)
    --           It gives several kinds of Informations, and allows to consider
    --           various criteria (criteria are cumulative)

uses Integer, Boolean, Transient, Type,
     HSequenceOfInteger,
     Check, Binder, StatusExec, HSequenceOfBinder

raises NoSuchObject

is

    	-- --    Building the Iterator    -- --

    Create returns TransferIterator;
    ---Purpose : Creates an empty Iterator

    AddItem (me : in out; atr : Binder)  is static;
    ---Purpose : Adds a Binder to the iteration list (construction)

    SelectBinder (me : in out; atype : Type; keep : Boolean)  is static;
    ---Purpose : Selects Items on the Type of Binder : keep only
    --           Binders which are of a given Type (if keep is True) or
    --           reject only them (if keep is False)

    SelectResult (me : in out; atype : Type; keep : Boolean)  is static;
    ---Purpose : Selects Items on the Type of Result. Considers only Unique
    --           Results. Considers Dynamic Type for Transient Result,
    --           Static Type (the one given to define the Binder) else.
    --         
    --           Results which are of a given Type (if keep is True) or reject
    --           only them (if keep is False)

    SelectUnique (me : in out; keep : Boolean)  is static;
    ---Purpose : Select Items according Unicity : keep only Unique Results (if
    --           keep is True) or keep only Multiple Results (if keep is False)

    SelectItem   (me : in out; num : Integer; keep : Boolean);
    ---Purpose : Selects/Unselect (according to <keep> an item designated by
    --           its rank <num> in the list
    --           Used by sub-classes which have specific criteria

    	-- --    Queries (Iteration, etc...)    -- --

    Number (me) returns Integer is static;
    ---Purpose : Returns count of Binders to be iterated

    Start (me : in out)  is static;
    ---Purpose : Clears Iteration in progress, to allow it to be restarted

    More (me : in out) returns Boolean  is static;
    ---Purpose : Returns True if there are other Items to iterate

    Next (me : in out)  is static;
    ---Purpose : Sets Iteration to the next Item

    Value (me) returns Binder
    ---Purpose : Returns the current Binder
    	raises NoSuchObject  is static;
    --           Error if Iteration has ended
    --           Some remarkable data can be accessed by following methods :
    ---C++ : return const &


    HasResult (me) returns  Boolean  raises NoSuchObject  is static;
    ---Purpose : Returns True if current Item brings a Result, Transient
    --           (Handle) or not or Multiple. That is to say, if it corresponds
    --           to a normally acheived Transfer, Transient Result is read by
    --           specific TransientResult below.
    --           Other kind of Result must be read specifically from its Binder

    HasUniqueResult (me) returns  Boolean  raises NoSuchObject  is static;
    ---Purpose : Returns True if Current Item has a Unique Result

    ResultType (me) returns Type  raises NoSuchObject  is static;
    ---Purpose : Returns the Type of the Result of the current Item, if Unique.
    --           If No Unique Result (Error Transfert or Multiple Result),
    --           returns a Null Handle
    --           The Type is : the Dynamic Type for a Transient Result,
    --           the Type defined by the Binder Class else

    HasTransientResult  (me) returns Boolean  raises NoSuchObject  is static;
    ---Purpose : Returns True if the current Item has a Transient Unique
    --           Result (if yes, use TransientResult to get it)

    TransientResult (me) returns any Transient
    	raises NoSuchObject  is static;
    ---Purpose : Returns the Transient Result of the current Item if there is
    --           (else, returns a null Handle)
    --           Supposes that Binding is done by a SimpleBinderOfTransient
    ---C++ : return const &


    Status (me) returns StatusExec  is static;
    ---Purpose : Returns Execution Status of current Binder
    --           Normal transfer corresponds to StatusDone

    HasFails (me) returns Boolean  is static;
    ---Purpose : Returns True if Fail Messages are recorded with the current
    --           Binder. They can then be read through Check (see below)

    HasWarnings (me) returns Boolean  is static;
    ---Purpose : Returns True if Warning Messages are recorded with the current
    --           Binder. They can then be read through Check (see below)

    Check  (me) returns Check  is static;
    ---Purpose : Returns Check associated to current Binder
    --           (in case of error, it brings Fail messages)
    --           (in case of warnings, it brings Warning messages)
    ---C++ : return const

fields

    theitems  : HSequenceOfBinder;
    theselect : HSequenceOfInteger;
    themaxi   : Integer;
    thecurr   : Integer  is protected;   -- for read by sub-classes

end TransferIterator;
