-- Created on: 1995-12-06
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package BRepCheck 

	---Purpose: This package  provides tools to check the validity
	--          of the BRep.

uses MMgt,
     StdFail,
     TCollection,
     TopAbs,
     Adaptor3d,
     TopoDS,
     BRep,
     TopTools

is

    deferred class Result;   -- inherits TShared from MMgt
    
    class Vertex;            -- inherits Shape
    
    class Edge;              -- inherits Shape
    
    class Wire;              -- inherits Shape
    
    class Face;              -- inherits Shape
    
    class Shell;             -- inherits Shape
    
--    class Solid;             -- inherits Shape

    class Analyzer;


    enumeration Status is
      NoError,
      
      -- for vertices
      InvalidPointOnCurve,
      InvalidPointOnCurveOnSurface,
      InvalidPointOnSurface,
            
      -- for edges
      No3DCurve,
      Multiple3DCurve,
      Invalid3DCurve,
      NoCurveOnSurface,
      InvalidCurveOnSurface,
      InvalidCurveOnClosedSurface,
      InvalidSameRangeFlag,
      InvalidSameParameterFlag,
      InvalidDegeneratedFlag,
      
      FreeEdge,
      InvalidMultiConnexity,
      InvalidRange,
      
      
      -- for wires
      EmptyWire,
      RedundantEdge,
      SelfIntersectingWire, -- on a face

      -- for faces
      NoSurface,
      InvalidWire,
      RedundantWire,
      IntersectingWires,
      InvalidImbricationOfWires,

      -- for shells
      EmptyShell,
      RedundantFace,


      -- for shapes
      UnorientableShape,
      NotClosed,
      NotConnected,
      
      SubshapeNotInShape,
      
      BadOrientation,
      BadOrientationOfSubshape,
      
      InvalidPolygonOnTriangulation,

      InvalidToleranceValue,

      -- for exception
      CheckFail
    
    end Status;


    class ListOfStatus instantiates List from TCollection
        (Status from BRepCheck);
       
    class DataMapOfShapeListOfStatus instantiates DataMap from TCollection 
        (Shape          from TopoDS,
       	 ListOfStatus   from BRepCheck,
         ShapeMapHasher from TopTools);
	
	
    class DataMapOfShapeResult instantiates DataMap from TCollection
    	(Shape          from TopoDS,
       	 Result         from BRepCheck,
         OrientedShapeMapHasher from TopTools);
	 
	 
    -- Package method

    Add(List: in out ListOfStatus from BRepCheck; 
        Stat: Status from BRepCheck);



    Print(Stat: Status from BRepCheck;
          OS: in out OStream from Standard);

    SelfIntersection(W      : Wire from TopoDS;
    	    	   F      : Face from TopoDS;
                   E1 : out Edge from TopoDS;
                   E2 : out Edge from TopoDS)
      returns Boolean from Standard;
      
end BRepCheck;
