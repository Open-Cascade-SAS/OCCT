-- Created on: 2002-03-04
-- Created by: Michael KLOKOV
-- Copyright (c) 2002-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class SectionAttribute from BOPAlgo
    ---Purpose: Class is a container of three flags used
    ---         by intersection algorithm
    ---

is

    Create(Aproximation : Boolean from Standard = Standard_True;
           PCurveOnS1   : Boolean from Standard = Standard_True;
           PCurveOnS2   : Boolean from Standard = Standard_True)
    returns SectionAttribute from BOPAlgo;
    ---Purpose:
    --- Initializes me by flags
    
    Approximation(me: in out; theFlag: Boolean from Standard);
    ---Purpose:
    --- Modifier
    ---
    
    PCurveOnS1(me: in out; theFlag: Boolean from Standard);
    ---Purpose:
    --- Modifier
    ---
    
    PCurveOnS2(me: in out; theFlag: Boolean from Standard);
    ---Purpose:
    --- Modifier
    ---

    Approximation(me)
    returns Boolean from Standard;
    ---C++: inline
    ---Purpose:
    --- Selector
    ---
    
    PCurveOnS1(me)
    returns Boolean from Standard;
    ---C++: inline
    ---Purpose:
    --- Selector
    ---
    
    PCurveOnS2(me)
    returns Boolean from Standard;
    ---C++: inline
    ---Purpose:
    --- Selector
    ---

fields
    myApproximation : Boolean from Standard;
    myPCurve1       : Boolean from Standard;
    myPCurve2       : Boolean from Standard;

end SectionAttribute from BOPAlgo;
