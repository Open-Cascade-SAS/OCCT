-- Created on: 2009-03-20
-- Created by: ABD
-- Copyright (c) 2009-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class LayerItem from Visual3d inherits TShared from MMgt

    ---Version:

    ---Purpose: This class is drawable unit of 2d scene
    ---Keywords:
    ---Warning:
    ---References:

uses
    Boolean from Standard
is
    -------------------------
    -- Category: Constructors
    -------------------------

    Create returns LayerItem;
    ---Level: Public
    ---Purpose: Creates a layer item
    ---Category: Constructors

    ---------------------------------------------------
    -- Category: Methods to modify the class definition
    ---------------------------------------------------
    
    ComputeLayerPrs( me : mutable )
            is virtual; 
    ---Level: Public
    ---Purpose: virtual function for recompute 2D
    --        presentation (empty by default)

    RedrawLayerPrs( me : mutable )
        is virtual;
    ---Level: Public
    ---Purpose: virtual function for recompute 2D
    --        presentation (empty by default)

        IsNeedToRecompute(me)
        returns Boolean from Standard;
    ---Level: Public
        
        SetNeedToRecompute( me                 : mutable;
                            NeedToRecompute    : Boolean from Standard = Standard_True );
    ---Level: Public

fields

    MyIsNeedToRecompute : Boolean from Standard;
    
end Layer from Visual3d;
