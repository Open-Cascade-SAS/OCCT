-- File:	MeshAlgo.cdl
-- Created:	Tue May 11 16:03:43 1993
-- Author:	Didier PIFFAULT
--		<dpf@nonox>
---Copyright:	 Matra Datavision 1993, 1994


package MeshAlgo 

	---Purpose: Manages different algorithms for triangulation.
	--          (like Delaunay)


        ---Level : Advanced.  
        --  All methods of all  classes will be advanced.


uses    Standard,
	gp,
	TCollection,
	SortTools,
	TColStd,
	Bnd,
    	MeshDS


is	
        imported CellFilter from MeshAlgo;
	
        imported CircleInspector from MeshAlgo;

        deferred class Vertex from MeshAlgo;     -- signature

      	deferred class Edge from MeshAlgo;       -- signature

      	deferred class Triangle from MeshAlgo;   -- signature
	
	class Circ from MeshAlgo;
	
      	class CircleTool from MeshAlgo;


      	generic class PntComparator from MeshAlgo;


      	generic class IndexedPntComparator from MeshAlgo;


	generic class Delaunay from MeshAlgo, DataStructure,
    	    	    	ComparatorOfVertex, ComparatorOfIndexedVertex,
    	    	    	Array1OfVertex, HArray1OfVertex, 
    	    	    	HeapSortVertex, HeapSortIndexedVertex;

end MeshAlgo;
