-- File:	StepData_ECDescr.cdl
-- Created:	Fri May  9 15:46:04 1997
-- Author:	Christian CAILLET
--		<cky@heliox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1997


class ECDescr  from StepData    inherits EDescr  from StepData

    ---Purpose : Describes a Complex Entity (Plex) as a list of Simple ones

uses HSequenceOfAsciiString from TColStd, SequenceOfTransient from TColStd,
     ESDescr from StepData, Described from StepData

is

    Create returns mutable ECDescr;
    ---Purpose : Creates an ECDescr, empty

    Add (me : mutable; member : ESDescr);
    ---Purpose : Adds a member
    --  Warning : members are added in alphabetic order

    NbMembers (me) returns Integer;
    ---Purpose : Returns the count of members

    Member (me; num : Integer) returns ESDescr;
    ---Purpose : Returns a Member from its rank

    TypeList (me) returns HSequenceOfAsciiString;
    ---Purpose : Returns the ordered list of types


    	--  inherited

    Matches    (me; steptype : CString) returns Boolean;
    ---Purpose : Tells if a ESDescr matches a step type : exact or super type

    IsComplex  (me) returns Boolean;
    ---Purpose : Returns True

    NewEntity  (me) returns mutable Described;
    ---Purpose : Creates a described entity (i.e. a complex one, made of one
    --           simple entity per member)

fields

    thelist : SequenceOfTransient;

end ECDescr;
