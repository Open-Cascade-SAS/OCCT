-- Created on: 1999-10-11
-- Created by: Atelier CAS2000
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package  BRepOffsetAPI 

uses   
    Standard, 
    StdFail,
    gp, 
    GeomAbs,
    Geom,
    GeomFill,
    Approx,
    TopoDS,
    TopTools, 
    BRepAlgo,
    BRepBuilderAPI, 
    BRepSweep, 
    BRepPrimAPI,  	     
    BRepFill, 
    Law, 
    Draft, 
    BRepOffset, 
     
    TColStd,
    TCollection

is 


    --
    -- Sweeping
    -- 

    class MakePipe;        ---  inherits MakeSweep from BRepPrimAPI    

    class MakePipeShell;  ---  inherits MakeSweep from BRepPrimAPI

    class  MakeDraft; ---  inherits MakeShape from BRepBuilderAPI
    
    class DraftAngle; ---  inherits MakeShape from BRepBuilderAPI




    class FindContigousEdges;

    alias Sewing  is  Sewing from BRepBuilderAPI;
      ---Purpose: sew the shapes along their common edges
   


    --
    -- Evolved and Offseting
    -- 
    
    class MakeOffset;     ---  inherits MakeShape from BRepBuilderAPI

    class MakeOffsetShape; ---  inherits MakeShape from BRepBuilderAPI
    	--Purpose: Offset shape to shells or solids.

    class MakeThickSolid;    ---   inherits MakeOffsetShape from BRepOffsetAPI

    class MakeEvolved;    ---  inherits MakeShape from BRepBuilderAPI

 
    --
    -- Construction of Shape through sections.
    -- 

    class ThruSections;	      ---  inherits  MakeShape  from  BRepBuilderAPI

    class NormalProjection ;  ---  inherits  MakeShape  from  BRepBuilderAPI

    class MiddlePath;	      ---  inherits  MakeShape  from  BRepBuilderAPI
    
    -- 
    --   Plate
    --     
    class MakeFilling;  ---  inherits MakeShape from BRepBuilderAPI

    class SequenceOfSequenceOfReal instantiates 
    	Sequence from TCollection (SequenceOfReal from TColStd);

    class SequenceOfSequenceOfShape instantiates 
    	Sequence from TCollection (SequenceOfShape from TopTools);

end;
