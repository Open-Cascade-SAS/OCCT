-- Created on: 2001-12-13
-- Created by: Sergey KUUl
-- Copyright (c) 2001-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class TimerSentry from MoniTool

    ---Purpose: A tool to facilitate using MoniTool_Timer functionality
    --          by automatically ensuring consistency of start/stop actions
    --
    --          When instance of TimerSentry is created, a timer 
    --          with corresponding name is started
    --          When instance is deleted, timer stops

uses
    Timer from MoniTool
    
is

    Create (cname: CString from Standard) 
    returns TimerSentry from MoniTool;
        ---C++: inline
        ---Purpose: Constructor creates an instance and runs the corresponding timer
    
    Create (timer: Timer from MoniTool) 
    returns TimerSentry from MoniTool;
        ---C++: inline
        ---Purpose: Constructor creates an instance and runs the corresponding timer
    
    Destroy(me: in out);
        ---C++: inline
    	---Purpose: Destructor stops the associated timer
        ---C++: alias "Standard_EXPORT ~MoniTool_TimerSentry () { Destroy(); }"

    Timer (me) returns Timer from MoniTool;
        ---C++: inline

    Stop (me: in out);
        ---C++: inline
    	---Purpose: Manually stops the timer

fields

    myTimer: Timer from MoniTool;

end TimerSentry;
