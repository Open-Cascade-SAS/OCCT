-- Created on: 1992-09-22
-- Created by: Christian CAILLET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Graph from Interface

    	---Purpose : Gives basic data structure for operating and storing
    	--           graph results (usage is normally internal)
    	--           Entities are Mapped according their Number in the Model
    	--           
    	--           Each Entity from the Model can be known as "Present" or
    	--           not; if it is, it is Mapped with a Status : an Integer
    	--           which can be used according to needs of each algorithm
    	--           In addition, the Graph brings a BitMap which can be used
    	--           by any caller
    	--           
    	--           Also, it is bound with two lists : a list of Shared
    	--           Entities (in fact, their Numbers in the Model) which is
    	--           filled by a ShareTool, and a list of Sharing Entities,
    	--           computed by deduction from the Shared Lists
    	--           
    	--           Moreover, it is possible to redefine the list of Entities
    	--           Shared by an Entity (instead of standard answer by general
    	--           service Shareds) : this new list can be empty; it can
    	--           be changed or reset (i.e. to come back to standard answer)

uses  Transient, Type,
      HArray1OfInteger from TColStd,
      HArray1OfTransient from TColStd,
      HSequenceOfTransient from TColStd,
      HArray1OfListOfInteger  from TColStd,
      AsciiString from TCollection, HAsciiString from TCollection,
      Protocol from Interface,  GeneralLib,      InterfaceModel,   GTool,
      EntityIterator, BitMap

raises DomainError

is

    Create (amodel : InterfaceModel; lib : GeneralLib; theModeStats : Boolean = Standard_True ) returns Graph;
    ---Purpose : Creates an empty graph, ready to receive Entities from amodel
    --           Note that this way of Creation allows <me> to verify that
    --           Entities to work with are contained in <amodel>
    --           Basic Shared and Sharing lists are obtained from a General
    --           Services Library, given directly as an argument

    Create (amodel : InterfaceModel; protocol : Protocol from Interface;
    theModeStats : Boolean = Standard_True)
    	returns Graph;
    ---Purpose : Same as above, but the Library is defined through a Protocol

    Create (amodel : InterfaceModel; gtool    : GTool from Interface;
		theModeStats : Boolean = Standard_True)
    	returns Graph;
    ---Purpose : Same as above, but the Library is defined through a Protocol

    Create (amodel : InterfaceModel;theModeStats : Boolean = Standard_True) returns Graph;
    ---Purpose : Same a above but works with the Protocol recorded in the Model
    
     Create (agraph : Graph; copied : Boolean = Standard_False) returns Graph;
    ---Purpose : Creates a Graph from another one, getting all its data
    --           Remark that status are copied from <agraph>, but the other
    --           lists (sharing/shared) are copied only if <copied> = True

    
    Evaluate (me : in out )  is static private;
    ---Purpose : Performs the Evaluation of the Graph, from an initial Library,
    --           either defined through a Protocol, or given dierctly
    --           Called by the non-empty Constructors
    --           
    --           Normally, gtool suffices. But if a Graph is created from a
    --           GeneralLib directly, it cannot be used
    --           If <gtool> is defined, it has priority


    Reset (me : in out)  is static;
    ---Purpose : Erases data, making graph ready to rebegin from void
    --           (also resets Shared lists redefinitions)

    ResetStatus (me : in out)  is static;
    ---Purpose : Erases Status (Values and Flags of Presence), making graph
    --           ready to rebegin from void. Does not concerns Shared lists

    Size (me) returns Integer  is static;
    ---Purpose : Returns size (max nb of entities, i.e. Model's nb of entities)

    	-- --    Fine Actions    -- --
    	
	NbStatuses(me) returns Integer;
	 ---Purpose : Returns size of array of statuses

    EntityNumber (me; ent : Transient) returns Integer  is static;
    ---Purpose : Returns the Number of the entity in the Map, computed at
    --           creation time (Entities loaded from the Model)
    --           Returns 0 if <ent> not contained by Model used to create <me>
    --           (that is, <ent> is unknown from <me>)

    IsPresent (me; num : Integer) returns Boolean  is static;
    ---Purpose : Returns True if an Entity is noted as present in the graph
    --           (See methods Get... which determine this status)
    --           Returns False if <num> is out of range too

    IsPresent (me; ent : Transient) returns Boolean;
    ---Purpose : Same as above but directly on an Entity <ent> : if it is not
    --           contained in the Model, returns False. Else calls
    --            IsPresent(num)  with <num> given by EntityNumber

    Entity (me; num : Integer) returns any Transient  is static;
    ---Purpose : Returns mapped Entity given its no (if it is present)
    ---C++ : return const &

    Status (me; num : Integer) returns Integer  is static;
    ---Purpose : Returns Status associated to a numero (only to read it)

    SetStatus (me : in out; num : Integer; stat : Integer)  is static;
    ---Purpose : Modifies Status associated to a numero

    RemoveItem (me : in out; num : Integer)  is static;
    ---Purpose : Clears Entity and sets Status to 0, for a numero

    ChangeStatus (me : in out; oldstat, newstat : Integer)  is static;
    ---Purpose : Changes all status which value is oldstat to new value newstat

    RemoveStatus (me : in out; stat : Integer)  is static;
    ---Purpose : Removes all items of which status has a given value stat

    BitMap (me) returns BitMap;
    ---Purpose : Returns the Bit Map in order to read or edit flag values
    ---C++ : return const &

    CBitMap (me : in out) returns BitMap;
    ---Purpose : Returns the Bit Map in order to edit it (add new flags)
    ---C++ : return &

    	-- --    General Actions    -- --

    Model (me) returns InterfaceModel  is static;
    ---Purpose : Returns the Model with which this Graph was created
    ---C++ : return const &

    GetFromModel (me : in out)  is static;
    ---Purpose : Loads Graph with all Entities contained in the Model

    GetFromEntity (me : in out; ent : Transient; shared : Boolean;
    	       newstat : Integer = 0)  is static;
    ---Purpose : Gets an Entity, plus its shared ones (at every level) if
    --           "shared" is True. New items are set to status "newstat"
    --           Items already present in graph remain unchanged
    --           Of course, redefinitions of Shared lists are taken into
    --           account if there are some

    GetFromEntity (me : in out; ent : Transient; shared : Boolean;
	     newstat, overlapstat : Integer; cumul : Boolean)
	 is static;
    ---Purpose : Gets an Entity, plus its shared ones (at every level) if
    --           "shared" is True. New items are set to status "newstat".
    --           Items already present in graph are processed as follows :
    --           - if they already have status "newstat", they remain unchanged
    --           - if they have another status, this one is modified :
    --             if cumul is True,  to former status + overlapstat (cumul)
    --             if cumul is False, to overlapstat (enforce)

    GetFromIter (me : in out; iter : EntityIterator; newstat : Integer)
    	is static;
    ---Purpose : Gets Entities given by an EntityIterator. Entities which were
    --           not yet present in the graph are mapped with status "newstat"
    --           Entities already present remain unchanged

    GetFromIter (me : in out; iter : EntityIterator;
	     newstat, overlapstat : Integer; cumul : Boolean)
	 is static;
    ---Purpose : Gets Entities given by an EntityIterator and distinguishes
    --           those already present in the Graph :
    --           - new entities added to the Graph with status "newstst"
    --           - entities already present with status = "newstat" remain
    --             unchanged
    --           - entities already present with status different form
    --             "newstat" have their status modified :
    --             if cumul is True,  to former status + overlapstat (cumul)
    --             if cumul is False, to overlapstat (enforce)
    --             (Note : works as GetEntity, shared = False, for each entity)

    GetFromGraph (me : in out; agraph : Graph)
    ---Purpose : Gets all present items from another graph
    	raises DomainError  is static;
    --           Error if the other graph has not been created with same Model

    GetFromGraph (me : in out; agraph : Graph; stat : Integer)
    ---Purpose : Gets items from another graph which have a specific Status
    	raises DomainError  is static;
    --           Error if the other graph has not been created with same Model

    	-- --    Shared Lists    -- --

    HasShareErrors (me; ent : Transient) returns Boolean  is static;
    ---Purpose : Returns True if <ent> or the list of entities shared by <ent>
    --           (not redefined) contains items unknown from this Graph
    --           Remark : apart from the status HasShareError, these items
    --           are ignored

    GetShareds(me; ent : Transient) returns HSequenceOfTransient;
	---Purpose : Returns the sequence of Entities Shared by an Entity
	
    Shareds (me; ent : Transient) returns EntityIterator
    ---Purpose : Returns the list of Entities Shared by an Entity, as recorded
    --           by the Graph. That is, by default Basic Shared List, else it
    --           can be redefined by methods SetShare, SetNoShare ... see below
    	raises DomainError  is static;
    --           Error if <ent> is not contained by the model used for Creation
  

    Sharings (me; ent : Transient) returns EntityIterator
    ---Purpose : Returns the list of Entities which Share an Entity, computed
    --           from the Basic or Redefined Shared Lists
    	raises DomainError  is static;
    --           Error if <ent> is not contained by the model used for Creation

   
	GetSharings(me; ent : Transient) returns HSequenceOfTransient;
	---Purpose : Returns the sequence of Entities Sharings by an Entity
	
	TypedSharings (me; ent : Transient; type : Type) returns EntityIterator;
    ---Purpose : Returns the list of sharings entities, AT ANY LEVEL, which are
    --           kind of a given type. A sharing entity kind of this type
    --           ends the exploration of its branch
	
    RootEntities (me) returns EntityIterator  is static;
    ---Purpose : Returns the Entities which are not Shared (their Sharing List
    --           is empty) in the Model

    	-- --    Redefinitions of Shared-Sharing Lists    -- --


    Name (me; ent : Transient) returns HAsciiString;
    ---Purpose : Determines the name attached to an entity, by using the
    --           general service Name in GeneralModule
    --           Returns a null handle if no name could be computed or if
    --           the entity is not in the model
    
       
    SharingTable (me) returns  HArray1OfListOfInteger  from TColStd; --HArray1OfTransient from TColStd ;
    ---C++ : return const &
    ---Purpose : Returns the Table of Sharing lists. Used to Create
    --           another Graph from <me>
    
    InitStats(me : in out) is protected;
    ---Purpose : Initialize statuses and flags
    
    ModeStat(me) returns Boolean;
    ---Purpose : Returns mode resposible for computation of statuses;
   	
fields

    themodel    : InterfaceModel is protected ;   -- Model which contains the Entities
    thepresents : AsciiString from TCollection is protected ; -- flags present/or not
    thestats    : HArray1OfInteger from TColStd is protected; -- numeric status
    theflags    : BitMap;                       -- logical flags status
    thesharings : HArray1OfListOfInteger  from TColStd is protected;       --HArray1OfTransient from TColStd is protected;
        
end Graph;
