-- Created on: 1993-07-21
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MakeCone from BRepPrimAPI  inherits MakeOneAxis from BRepPrimAPI

	---Purpose: Describes functions to build cones or portions of cones.
    	-- A MakeCone object provides a framework for:
    	-- -   defining the construction of a cone,
    	-- -   implementing the construction algorithm, and
    	-- -   consulting the result.

uses
    Ax2      from gp,
    Cone     from BRepPrim,
    OneAxis  from BRepPrim

raises
    DomainError from Standard

is
    Create(R1, R2, H : Real)
    returns MakeCone from BRepPrimAPI
	---Purpose: Make a cone of height H radius R1 in the plane z =
	--          0, R2 in the plane Z = H. R1 and R2 may be null.
	---Level: Public
    raises
    	DomainError from Standard; -- if H <= Precision::Confusion()

    Create(R1, R2, H, angle : Real)
    returns MakeCone from BRepPrimAPI
	---Purpose: Make a cone of height H radius R1 in the plane z =
	--          0, R2 in the plane Z = H. R1 and R2 may be null.
	--          Take a section of <angle>
	---Level: Public
    raises
    	DomainError from Standard; -- if H <= Precision::Confusion()

    Create(Axes : Ax2 from gp; R1, R2, H : Real)
    returns MakeCone from BRepPrimAPI
	---Purpose: Make a cone of height H radius R1 in the plane z =
	--          0, R2 in the plane Z = H. R1 and R2 may be null.
	---Level: Public
    raises
    	DomainError from Standard; -- if H <= Precision::Confusion()

    Create(Axes : Ax2 from gp; R1, R2, H, angle : Real)
    returns MakeCone from BRepPrimAPI
	---Purpose: Make a cone of height H radius R1 in the plane z =
	--          0, R2 in the plane Z = H. R1 and R2 may be null.
	--          Take a section of <angle>
	---Level: Public
    raises
    	DomainError from Standard; -- if H <= Precision::Confusion()

    	---Purpose: Constructs a cone, or a portion of a cone, of height H,
    	-- and radius R1 in the plane z = 0 and R2 in the plane
    	-- z = H. The result is a sharp cone if R1 or R2 is equal to 0.
    	-- The cone is constructed about the "Z Axis" of either:
    	-- -   the global coordinate system, or
    	-- -   the local coordinate system Axes.
    	-- It is limited in these coordinate systems as follows:
    	-- -   in the v parametric direction (the Z coordinate), by
    	--   the two parameter values 0 and H,
    	-- -   and in the u parametric direction (defined by the
    	--   angle of rotation around the Z axis), in the case of a
    	--   portion of a cone, by the two parameter values 0 and
    	--   angle. Angle is given in radians.
    	-- The resulting shape is composed of:
    	-- -   a lateral conical face
    	-- -   two planar faces in the planes z = 0 and z = H,
    	--   or only one planar face in one of these two planes if a
    	--   radius value is null (in the case of a complete cone,
    	--   these faces are circles), and
    	-- -   and in the case of a portion of a cone, two planar
    	--   faces to close the shape. (either two parallelograms or
    	--   two triangles, in the planes u = 0 and u = angle).    
    	-- Exceptions
    	-- Standard_DomainError if:
    	-- -   H is less than or equal to Precision::Confusion(), or
    	-- -   the half-angle at the apex of the cone, defined by
    	--   R1, R2 and H, is less than Precision::Confusion()/H, or greater than
    	--   (Pi/2)-Precision::Confusion()/H.f
        
    OneAxis(me : in out) returns Address;
	---Purpose: Returns the algorithm.
	---Level: Public

    Cone(me : in out) returns Cone from BRepPrim
	---Purpose: Returns the algorithm.
	--          
	---C++: return &
	---Level: Public
    is static;

fields 

    myCone : Cone from BRepPrim;

end MakeCone;
