-- Created on: 1993-07-06
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class CurveOn2Surfaces from BRep inherits CurveRepresentation from BRep

	---Purpose: Defines a continuity between two surfaces.

uses
    Pnt      from gp,
    Surface  from Geom,
    Location from TopLoc,
    Shape    from GeomAbs,
    CurveRepresentation from BRep
    
raises
    NullObject from Standard
    
is

    Create(S1 , S2  : Surface  from Geom;
	   L1 , L2  : Location from TopLoc;
	   C        : Shape    from GeomAbs)
    returns mutable CurveOn2Surfaces from BRep;

    IsRegularity(me) returns Boolean
	---Purpose: Returns True.
    is redefined;
    
    IsRegularity(me; S1,S2 : Surface from Geom; 
                     L1,L2 : Location from TopLoc)  
    returns Boolean
	---Purpose: A curve on two surfaces (continuity). 
    is redefined;

    D0(me; U : Real; P : out Pnt from gp);
	---Purpose: Raises an error.
    
    Surface(me) returns any Surface from Geom
	---C++: return const &
    is redefined;

    Surface2(me) returns any Surface from Geom
	---C++: return const &
    is redefined;

    Location2(me) returns Location from TopLoc
	---C++: return const &
    is redefined;

    Continuity(me) returns Shape from GeomAbs
	---C++: return const &
    is redefined;
    
    Continuity(me : mutable; C : Shape from GeomAbs)
    is redefined;
    
    Copy(me) returns mutable CurveRepresentation from BRep;
	---Purpose: Return a copy of this representation.

fields
    mySurface    : Surface from Geom;
    mySurface2   : Surface from Geom;
    myLocation2  : Location from TopLoc;
    myContinuity : Shape from GeomAbs;

end CurveOn2Surfaces;
