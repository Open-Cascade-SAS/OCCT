-- Created on: 1997-02-10
-- Created by: Alexander BRIVIN
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class FontStyle from Vrml 

	---Purpose: defines a FontStyle node of VRML of properties of geometry
	--  and its appearance. 
	--  The  size  field  specifies  the  height  (in  object  space  units) 
    	--  of  glyphs  rendered  and  determines  the  vertical  spacing  of 
	--  adjacent  lines  of  text.

uses
 
    FontStyleFamily from Vrml, 
    FontStyleStyle  from Vrml
  
is
 
    Create  (  aSize    :  Real            from Standard  =  10;
    	       aFamily  :  FontStyleFamily from Vrml      =  Vrml_SERIF;
    	       aStyle   :  FontStyleStyle  from Vrml      =  Vrml_NONE  ) 
	returns  FontStyle from Vrml;

    SetSize ( me : in out; aSize    :  Real from Standard  );
    Size ( me )  returns Real  from  Standard;

    SetFamily ( me : in out;  aFamily  :  FontStyleFamily from Vrml  ); 
    Family ( me )  returns FontStyleFamily from Vrml; 
     
    SetStyle ( me : in out;  aStyle   :  FontStyleStyle from Vrml ); 
    Style ( me )  returns  FontStyleStyle from Vrml; 
    
    Print  ( me;  anOStream: in out OStream from Standard) returns OStream from Standard;
    ---C++:  return  & 


fields
 
    mySize    :  Real            from Standard;  -- Font size
    myFamily  :  FontStyleFamily from Vrml;      -- Font family
    myStyle   :  FontStyleStyle  from Vrml;      -- Font style modifications to family

end FontStyle;
