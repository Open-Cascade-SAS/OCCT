-- Created on: 1994-11-04
-- Created by: Christian CAILLET
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class TransientElem from MoniTool inherits Element

    ---Purpose : an TransientElem defines an Element for a specific input class
    --           its definition includes the value of the Key to be mapped,
    --           and the HashCoder associated to the class of the Key
    --           
    --           Transient from Standard defines the class to be keyed
    --           MapTransientHasher from TColStd is the associated Hasher
    --           DataInfo from MoniTool   is an additionnal class which helps to provide
    --             informations on the value (template : see DataInfo)

uses CString,
     Transient          from Standard,
     MapTransientHasher from TColStd,
     DataInfo           from MoniTool

is

    Create (akey : any Transient from Standard) returns mutable TransientElem;
    ---Purpose : Creates a TransientElem with a Value. This Value can then not be
    --           changed. It is used by the Hasher to compute the HashCode,
    --           which will then be stored for an immediate reading.

    Value (me) returns any Transient from Standard  is static;
    ---Purpose : Returns the contained value
    ---C++ : return const &

    Equates (me; other : Element) returns Boolean;
    ---Purpose : Specific testof equallity : defined as False if <other> has
    --           not the same true Type, else contents are compared (by
    --           C++ operator ==)

    ValueType    (me) returns Type  is redefined;
    ---Purpose : Returns the Type of the Value. By default, returns the
    --           DynamicType of <me>, but can be redefined

    ValueTypeName (me) returns CString  is redefined;
    ---Purpose : Returns the name of the Type of the Value. Default is name
    --           of ValueType, unless it is for a non-handled object

fields

    theval  : Transient from Standard;

end TransientElem;
