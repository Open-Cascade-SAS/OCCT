-- Created on: 1992-08-21
-- Created by: Christophe MARION
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ShapeData from HLRTest inherits TShared from MMgt

    	---Purpose: Contains the colors of a shape.

uses
    Color from Draw
    
is
    Create(CVis,COVis,CIVis,CHid,COHid,CIHid : Color from Draw)
    returns mutable ShapeData from HLRTest; 
    
    VisibleColor(me: mutable; CVis : Color from Draw)
    	---C++: inline
    is static;

    VisibleOutLineColor(me: mutable; COVis : Color from Draw)
    	---C++: inline
    is static;

    VisibleIsoColor(me: mutable; CIVis : Color from Draw)
    	---C++: inline
    is static;

    HiddenColor(me: mutable; CHid : Color from Draw)
    	---C++: inline
    is static;

    HiddenOutLineColor(me: mutable; COHid : Color from Draw)
    	---C++: inline
    is static;

    HiddenIsoColor(me: mutable; CIHid : Color from Draw)
    	---C++: inline
    is static;

    VisibleColor(me) returns Color from Draw
    	---C++: inline
    is static;

    VisibleOutLineColor(me) returns Color from Draw
    	---C++: inline
    is static;

    VisibleIsoColor(me) returns Color from Draw
    	---C++: inline
    is static;

    HiddenColor(me)  returns Color from Draw
    	---C++: inline
    is static;

    HiddenOutLineColor(me)  returns Color from Draw
    	---C++: inline
    is static;

    HiddenIsoColor(me)  returns Color from Draw
    	---C++: inline
    is static;

fields
    myVColor  : Color from Draw;
    myVOColor : Color from Draw;
    myVIColor : Color from Draw;
    myHColor  : Color from Draw;
    myHOColor : Color from Draw;
    myHIColor : Color from Draw;

end ShapeData;
