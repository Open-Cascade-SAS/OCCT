-- Created on: 1997-05-13
-- Created by: Alexander BRIVIN
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class IsoAspect from VrmlConverter inherits LineAspect from VrmlConverter

 	---Purpose: qualifies the aspect properties for  
	--          the VRML conversation of iso curves . 

uses 

    Material    from   Vrml

is

    Create
    returns mutable IsoAspect from VrmlConverter;

    ---Purpose: create a default IsoAspect. 
    --  Default value: myNumber  - 10.

    Create  (aMaterial: Material from Vrml; 
    	    	 OnOff: Boolean from Standard;
               aNumber: Integer from Standard)
    returns mutable IsoAspect from VrmlConverter;
	    

    SetNumber (me: mutable; aNumber: Integer from Standard) 
    --Purpose: defines the number of U or V isoparametric curves 
    --         to be drawn for a single face.
    is static;

    Number (me) returns Integer from Standard 
    ---Purpose: returns the number of U or V isoparametric curves drawn for a
    --          single face.
    is static;

    
fields

    myNumber: Integer from Standard;

end IsoAspect;
