-- Created on: 1996-12-24
-- Created by: Alexander BRIVIN
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Cone from Vrml 

	---Purpose: defines a Cone node of VRML specifying geometry shapes.
    	-- This  node  represents  a  simple  cone,  whose  central  axis  is  aligned 
	-- with  the  y-axis.  By  default ,  the  cone  is  centred  at  (0,0,0) 
	-- and  has  size  of  -1  to  +1  in  the  all  three  directions. 
	-- the  cone  has  a  radius  of  1  at  the  bottom  and  height  of  2, 
	-- with  its  apex  at  1  and  its  bottom  at  -1.  The  cone  has  two  parts: 
	-- the  sides  and  the  bottom
uses
     
    ConeParts from Vrml
is

    Create ( aParts        : ConeParts from Vrml = Vrml_ConeALL; 
    	     aBottomRadius : Real      from Standard = 1; 
             aHeight       : Real      from Standard = 2 )  
        returns Cone from Vrml;
    
    SetParts ( me : in out; aParts : ConeParts from Vrml );
    Parts ( me )  returns  ConeParts from Vrml;

    SetBottomRadius ( me : in out; aBottomRadius : Real from Standard );
    BottomRadius ( me )  returns Real  from  Standard;

    SetHeight ( me : in out; aHeight : Real from Standard );
    Height ( me )  returns Real  from  Standard;

    Print  ( me;  anOStream: in out OStream from Standard) returns OStream from Standard;
    ---C++:  return  & 

fields

    myParts        : ConeParts from Vrml;      -- Visible parts of cone
    myBottomRadius : Real      from Standard;  -- Radius of bottom circular face
    myHeight       : Real      from Standard;  -- Size in y dimension
   
end Cone;
