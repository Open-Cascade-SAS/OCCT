-- Created on: 1991-04-04
-- Created by: Remi GILET
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


package GccGeo


    ---Purpose :
    -- This package provides an implementation of analytic algorithms
    -- (using only non-persistant entities) used to create 2d lines or
    -- circles with geometric constraints.

uses GccEnt,
     GccInt,
     IntCurve,
     GeomAbs,
     TColStd,
     Standard,
     StdFail,
     TColgp,
     gp

is

generic class CurvePGTool;

generic class ParGenCurve;

generic class Circ2dTanCen;
    -- Create a 2d circle TANgent to a 2d entity and CENtered on a 2d point.

generic class Circ2d2TanRad;
    -- Create a 2d circle TANgent to 2 2d entities with the given RADius.

generic class Circ2dTanOnRad;
    -- Create a 2d circle TANgent to a 2d entity and centered ON a 2d 
    -- entity (not a point) with the given radius.

generic class Circ2d2TanOn;
    -- Create a 2d circle TANgent to 2 2d entities (circle, line or point) 
    -- and centered ON a 2d curve.

end GccGeo;
