-- Created on: 1992-05-27
-- Created by: Remi LEQUETTE
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.





class TFace from BRep inherits TFace from TopoDS

	---Purpose: The Tface from BRep  is  based  on the TFace  from
	--          TopoDS. The TFace contains :
	--          
	--          * A suface, a tolerance and a Location.
	--          
	--          * A NaturalRestriction flag,   when this  flag  is
	--          True the  boundary of the  face is known to be the
	--          parametric space (Umin, UMax, VMin, VMax).
	--          
	--          *  An    optional Triangulation.   If  there  is a
	--          triangulation the surface can be absent.
	--          
	--          The  Location is  used   for the Surface.
	--          
	--          The triangulation  is in the same reference system
	--          than the TFace.     A point on mySurface must   be
	--          transformed with myLocation,  but  not a point  on
	--          the triangulation.
	--          
	--          The Surface may  be shared by different TFaces but
	--          not the  Triangulation, because the  Triangulation
	--          may be modified by  the edges. 
	--          
uses
    Surface       from Geom,
    Location      from TopLoc,
    TShape        from TopoDS,
    Triangulation from Poly
    
is

    Create returns mutable TFace from BRep;
	---Purpose: Creates an empty TFace.
	
    Surface(me) returns any Surface from Geom;
	---C++: inline
	---C++: return const &
    
    Triangulation(me) returns any Triangulation from Poly;
	---C++: inline
	---C++: return const &
    	
    Location(me) returns Location from TopLoc;
	---C++: inline
	---C++: return const &
    	
    Tolerance(me) returns Real;
	---C++: inline

    Surface(me : mutable; S : Surface from Geom);
	---C++: inline
    	
    Triangulation(me : mutable; T : Triangulation from Poly);
	---C++: inline
    	
    Location(me : mutable; L : Location from TopLoc);
	---C++: inline

    Tolerance(me : mutable; T : Real);
	---C++: inline

    NaturalRestriction(me) returns Boolean;
	---C++: inline
    
    NaturalRestriction(me : mutable; N : Boolean);
	---C++: inline
    
    EmptyCopy(me) returns mutable TShape from TopoDS
	---Purpose: Returns a copy  of the  TShape  with no sub-shapes.
	--          The new Face has no triangulation.
    is redefined;
    
fields

    mySurface            : Surface       from Geom;
    myTriangulation      : Triangulation from Poly;
    myLocation           : Location      from TopLoc;
    myTolerance          : Real;
    myNaturalRestriction : Boolean;

end TFace;

