-- Created on: 2009-05-05
-- Created by: Sergey ZARITCHNY <sergey.zaritchny@opencascade.com> 
-- Copyright (c) 2009-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class BooleanOperationDriver from DNaming inherits Driver from TFunction

	---Purpose: Driver  for Fuse,  Cut,  Common
uses
     Label            from TDF, 
     Logbook          from TFunction,
     Function         from TFunction,
     ExtendedString   from TCollection,
     BooleanOperation from BRepAlgoAPI

is
    Create returns mutable BooleanOperationDriver from DNaming;
    ---Purpose: Constructor

    ---Purpose: validation
    --          ==========

    Validate(me; theLog : in out Logbook from TFunction)
    is redefined;
    ---Purpose: Validates labels of a function in <log>.
    --          In regeneration mode this method must be called (by the
    --          solver) even if the function is not executed, to build
    --          the valid label scope.

    ---Purpose: execution of function
    --          ======================

    MustExecute (me; theLog : Logbook from TFunction)
    ---Purpose: Analyse in <log> if the loaded function must be executed
    --          (i.e.arguments are modified) or not.
    --          If the Function label itself is modified, the function must
    --          be executed.
    returns Boolean from Standard
    is redefined;

    Execute (me; theLog : in out Logbook from TFunction)
    ---Purpose: Execute the function and push in <log> the impacted
    --          labels (see method SetImpacted).
    returns Integer from Standard
    is redefined;
 
    LoadNamingDS(me; theResultLabel : Label from TDF; MS : in out BooleanOperation from BRepAlgoAPI)  
    is private; 

    LoadSectionNDS(me; theResultLabel : Label from TDF; MS : in out BooleanOperation from BRepAlgoAPI)  
    is private; 

    CheckAndLoad(me; theMkOpe : in out BooleanOperation from BRepAlgoAPI; 
    	    	     theFunction : Function from TFunction)   
    returns Boolean from Standard is private; 
    
end BooleanOperationDriver;


