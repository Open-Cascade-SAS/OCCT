-- File:	MeshDS.cdl
-- Created:	Mon Mar 15 17:47:36 1993
-- Author:	Didier PIFFAULT
--		<dpf@phylox>
---Copyright:	 Matra Datavision 1993


package MeshDS 

	---Purpose: This package  describes the common  data  structure for
	--          the differents MESH algorithms. 
        --  Level : Advanced.  
        --  All methods of all  classes will be advanced.

uses    Standard,
    	MMgt,
    	TCollection,
	gp,
	Bnd


is      enumeration DegreeOfFreedom is 
    	    Free,
	    InVolume,
    	    OnSurface,
    	    OnCurve,
    	    Fixed,
    	    Frontier,
    	    Deleted;
	    
        imported DataMapOfInteger from MeshDS;
	imported MapOfIntegerInteger from MeshDS;
	imported MapOfInteger from MeshDS;
	imported ListOfInteger from MeshDS;
	imported BaseAllocator from MeshDS;
	imported PairOfIndex from MeshDS;

	deferred generic class Node;       -- Signature

	deferred generic class Link;       -- Signature

	deferred generic class Element2d;  -- Signature
	
	generic class Mesh2d,   NodeHasher,
	       	    	    	LinkHasher, 
    	    	    	    	ElemHasher,
    	    	    	    	IDMapOfNode,
	       	    	    	IDMapOfLink, 
    	    	    	    	IMapOfElement,
    	    	    	    	Selector;


end MeshDS;
