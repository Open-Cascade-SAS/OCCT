-- Created on: 1999-09-13
-- Created by: data exchange team
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class FixSmallFace from ShapeFix inherits Root from ShapeFix

	---Purpose: Fixing face with small size

uses
    Shape from TopoDS,
    Face from TopoDS,
    Edge from TopoDS,
    Compound from TopoDS,
    CheckSmallFace from ShapeAnalysis
    
is
    Create returns FixSmallFace;
    ---Purpose :
    Init(me: mutable; S : Shape from TopoDS); 
    ---Purpose :
    
    Perform(me:mutable);	
    ---Purpose :
    -- Fixing case of spot face
    FixSpotFace (me: mutable) returns Shape from TopoDS;
    ---Purpose : Fixing case of spot face, if tol = -1 used local tolerance.
    ReplaceVerticesInCaseOfSpot(me; F : in out Face from TopoDS; tol : Real) returns Boolean;
    ---Purpose : Compute average vertex and replacing vertices by new one.

     RemoveFacesInCaseOfSpot(me; F :  Face from TopoDS) returns Boolean;
    ---Purpose : Remove spot face from compound
    --
    
     -- Fixing case of strip face   
     FixStripFace(me: mutable; wasdone: Boolean = Standard_False) returns Shape from TopoDS;
    ---Purpose : Fixing case of strip face, if tol = -1 used local tolerance

    ReplaceInCaseOfStrip(me;F : in out Face from TopoDS; E1 : in out  Edge from TopoDS; E2 : in out  Edge from TopoDS;tol : Real) returns Boolean;
    ---Purpose : Replace veretces and edges.
    --
    RemoveFacesInCaseOfStrip(me; F :  Face from TopoDS) returns Boolean;
    ---Purpose : Remove strip face from compound.
    
    ComputeSharedEdgeForStripFace(me; F :  Face from TopoDS; E1 : Edge from TopoDS; E2 : Edge from TopoDS; 
    F1 :  Face from TopoDS;     tol : Real ) 
    returns Edge from TopoDS;
    ---Purpose : Compute average edge for strip face

     -- Fixing case split
    
    FixSplitFace(me: mutable; S: Shape from TopoDS) returns Shape from TopoDS;
    ---Purpose : 
    --
    
    SplitFaces(me: mutable) returns Shape from TopoDS;
    ---Purpose : Split faces by splitting vertices
    --
    
    SplitOneFace(me: mutable; F : in out Face from TopoDS;theSplittedFaces: in out Compound from TopoDS) returns Boolean;
    ---Purpose : Compute data for face splitting.
    --
    
    RemoveSmallFaces(me:mutable) returns Shape from TopoDS;
    ---Purpose : Remove small faces from compound.
  
    --Fixes after removing
    FixFace(me: mutable; F: Face from TopoDS) returns Face from TopoDS;
    FixShape(me: mutable) returns Shape from TopoDS;

    Shape(me : mutable) returns Shape from TopoDS;
    
    FixPinFace (me: mutable;F : in out Face from TopoDS) returns Boolean;

fields

    myShape    : Shape from TopoDS;
    myResult   : Shape from TopoDS;
    myStatus   : Integer; -- error status
    myAnalyzer : CheckSmallFace from ShapeAnalysis;




end FixSmallFace;
