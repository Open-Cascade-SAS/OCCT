-- Created on: 1993-02-25
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class BlockIterator from BOP 

    ---Purpose:  
     
    --  Auxiliary class to provide 
    --  simple iteration on indexes that 
    --  belongs to the integer range  [Lower,Upper]  
    --  with increment =1 

raises

    NoMoreObject from Standard

is

    Create  
    	returns BlockIterator from BOP;
    	---Purpose:  
    	--- Empty  Constructor 
    	---
    Create(Lower,Upper : Integer from Standard) 
    	returns BlockIterator from BOP;
    	---Purpose:  
    	--- Creates an object with initial range 
    	--- of  [Lower,Upper]  	     
    	---
    
    Initialize(me : in out)  
    	is static;
    	---Purpose:  
    	--- Initialize an object with initial range 
    	--- of  [Lower,Upper]  	     
    	---
    More(me)  
    	returns Boolean from Standard  
    	is static;
    	---Purpose:  
    	--- Support of Iteration 
    	---
    Next(me : in out)  
    	raises NoMoreObject  
    	is static;
    	---Purpose:  
    	--- Support of Iteration 
    	---
    Value(me)  
    	returns Integer from Standard  
    	is static;
    	---Purpose:  
    	--- Support of Iteration 
    	---
    Extent(me)  
    	returns Integer from Standard  
    	is static;
    	---Purpose:  
    	--- Returns the extension=myUpper - myLower + 1;   
    	---
    
fields

    myLower : Integer from Standard;
    myUpper : Integer from Standard;
    myValue : Integer from Standard;

end BlockIterator;
