-- Created on: 1993-05-05
-- Created by: Christian CAILLET
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Protocol  from IGESSolid  inherits  Protocol from IGESData

    ---Purpose : Description of Protocol for IGESSolid

uses Type, Protocol from Interface

is

    Create returns mutable Protocol from IGESSolid;

    NbResources (me) returns Integer  is redefined;
    ---Purpose : Gives the count of Resource Protocol. Here, one
    --           (Protocol from IGESGeom)

    Resource (me; num : Integer) returns Protocol from Interface  is redefined;
    ---Purpose : Returns a Resource, given a rank.

    TypeNumber (me; atype : any Type) returns Integer  is redefined;
    ---Purpose : Returns a Case Number, specific of each recognized Type
    --           This Case Number is then used in Libraries : the various
    --           Modules attached to this class of Protocol must use them
    --           in accordance (for a given value of TypeNumber, they must
    --           consider the same Type as the Protocol defines)

end Protocol;
