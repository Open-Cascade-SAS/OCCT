-- Created by: Peter KURNEV
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

class PaveBlock from BOPDS 
    inherits TShared from MMgt  
    
---Purpose:  
-- The class BOPDS_PaveBlock is to store  
-- the information about pave block on an edge. 
-- Two adjacent paves on edge make up pave block.    

uses   
    Box from Bnd, 
    BaseAllocator from BOPCol, 
    MapOfInteger from BOPCol,
    Pave from BOPDS,
    ListOfPave from BOPDS, 
    ListOfPaveBlock from BOPDS,
    CommonBlock from BOPDS 
    
--raises

is 
    Create 
    returns mutable PaveBlock from BOPDS; 
    ---Purpose:  
    --- Empty contructor  
    --- 
    Create (theAllocator: BaseAllocator from BOPCol) 
    returns mutable PaveBlock from BOPDS; 
    ---Purpose:  
    ---  Contructor    
    ---  <theAllocator> - the allocator to manage the memory     
    --- 
     
    SetPave1(me:mutable; 
        thePave:Pave from BOPDS); 
    ---Purpose: 
    --- Modifier   
    --- Sets the first pave <thePave> 
     
    Pave1(me) 
    returns Pave from BOPDS; 
    ---C++: return const &     
    ---Purpose: 
    --- Selector 
    --- Returns the first pave        	 
     
    SetPave2(me:mutable; 
        thePave:Pave from BOPDS); 
    ---Purpose: 
    --- Modifier   
    --- Sets the second pave <thePave>     
     
    Pave2(me) 
    returns Pave from BOPDS; 
    ---C++: return const &  
    ---Purpose:  
    --- Selector 
    --- Returns the second pave 

    SetEdge(me:mutable; 
        theEdge:Integer from Standard); 
    ---Purpose: 
    --- Modifier   
    --- Sets the index of edge of pave block <theEdge>      
    Edge(me) 
        returns Integer from Standard;  
    ---Purpose:  
    --- Selector 
    --- Returns the index of edge of pave block
 
    HasEdge(me) 
    returns Boolean from Standard; 
    ---Purpose: 
    --- Query
    --- Returns true if the pave block has edge 
	 
    HasEdge(me; 
        theEdge:out Integer from Standard) 
    returns Boolean from Standard; 
    ---Purpose: 
    --- Query
    --- Returns true if the pave block has edge 
    --- Returns the index of edge <theEdge> 
	
    SetOriginalEdge  (me:mutable;   
        theEdge:Integer from Standard);  
    ---Purpose: 
    --- Modifier   
    --- Sets the index of original edge  
    --- of the pave block <theEdge>   
	 
    OriginalEdge(me) 
    returns Integer from Standard; 
    ---Purpose:  
    --- Selector 
    --- Returns the index of original edge of pave block 
	
    IsSplitEdge(me) 
    returns Boolean from Standard; 
    ---Purpose: 
    --- Query
    --- Returns true if the edge is equal to the original edge   
    --- of the pave block    
     
    Range(me; 
        theT1:out Real from Standard; 
        theT2:out Real from Standard);
    ---Purpose:  
    --- Selector 
    --- Returns the parametric range <theT1,theT2>  
    --- of the pave block  
     
    HasSameBounds(me; 
        theOther: PaveBlock from BOPDS) 
    returns Boolean from Standard; 
    ---Purpose: 
    --- Query
    --- Returns true if the pave block has pave indices   
    --- that equal to the  pave indices of the pave block   
    --- <theOther> 
	 
    Indices(me; 
        theIndex1:out Integer from Standard; 
        theIndex2:out Integer from Standard); 
    ---Purpose: 
    --- Selector 
    --- Returns the pave indices  <theIndex1,theIndex2>  
    --- of the pave block   
	
    -- 
    -- extras
    --  
    IsToUpdate(me) 
    returns Boolean from Standard; 
    ---Purpose:  
    --- Query
    --- Returns true if the pave block contains extra paves 
	 
    AppendExtPave(me:mutable; 
        theLP:Pave from BOPDS);  
    ---Purpose: 
    --- Modifier 
    --- Appends extra paves <theLP> 
	 
    AppendExtPave1(me:mutable; 
        thePave:Pave from BOPDS);  
    ---Purpose: 
    --- Modifier 
    --- Appends extra pave <thePave>     
      
    ExtPaves(me) 
    returns ListOfPave from BOPDS; 
    ---C++: return const &  
    ---Purpose: 
    --- Selector 
    --- Returns the  extra paves 
    
    ChangeExtPaves(me:mutable) 
    returns ListOfPave from BOPDS; 
    ---C++: return &  
    ---Purpose: 
    --- Selector / Modifier
    --- Returns the extra paves 
 
    Update(me:mutable; 
        theLPB  : out ListOfPaveBlock from BOPDS; 
        theFlag : Boolean from Standard=Standard_True);
    ---Purpose: 
    --- Modifier  
    --- Updates the pave block. The extra paves are used 
    --- to create new pave blocks <theLPB>. 
    --- <theFlag> - if true, the first pave and the second  
    --- pave are used to produce new pave blocks. 
	 
    ContainsParameter(me; 
        thePrm:Real from Standard; 
        theTol:Real from Standard) 
    returns Boolean from Standard; 
    ---Purpose: 
    --- Query 
    --- Returns true if the extra paves contain the pave 
    --- with given value of the parameter <thePrm> 
    ---  <theTol>  - the value of the tolerance to compare 
	 
    -- 
    -- common block   
    -- 
    SetCommonBlock(me:mutable; 
        theCB:CommonBlock from BOPDS); 
    ---Purpose: 
    --- Modifier  
    --- Sets the common block <theCB> 
	 
    CommonBlock(me) 
    returns CommonBlock from BOPDS;     
    ---C++: return const & 
    ---Purpose: 
    --- Selector  
    --- Returns the common block 
	 
    IsCommonBlock(me) 
    returns Boolean from Standard; 
    ---Purpose: 
    --- Query 
    --- Returns true if the pave block is common block    
     
    IsCommonBlockOnEdge(me)  
    returns Boolean from Standard; 	 
    ---Purpose: 
    --- Query 
    --- Returns true if the pave block is common block 
    --- that contains at least one pave block  
	 
    RealPaveBlock(me) 
    returns PaveBlock from BOPDS;  
    ---Purpose: 
    --- Selector  
    --- Returns the real common block  
    -- 
    -- shrunk data   
    -- 
    SetShrunkData(me:mutable;  
        theTS1:Real from Standard;
        theTS2:Real from Standard;
        theBox:Box from Bnd);  
    ---Purpose: 
    --- Modifier  
    --- Sets the shrunk data for the pave block 
    --- <theTS1>,  <theTS2> - shrunk range 
    --- <theBox> - the bounding box 
	 
    ShrunkData(me; 
        theTS1:out Real from Standard;
        theTS2:out Real from Standard;  
        theBox:out Box from Bnd);
    ---Purpose: 
    --- Selector
    --- Returns  the shrunk data for the pave block 
    --- <theTS1>,  <theTS2> - shrunk range 
    --- <theBox> - the bounding box  
	
    HasShrunkData(me) 
    returns Boolean from Standard; 
    ---Purpose: 
    --- Query 
    --- Returns true if the pave block contains 
    --- the shrunk data 
     
    Dump(me);


fields 
    --general 
    myAllocator : BaseAllocator from BOPCol is protected; 
    myEdge         :  Integer from Standard is protected; 
    myOriginalEdge :  Integer from Standard is protected;
    myPave1        :  Pave from BOPDS is protected;
    myPave2        :  Pave from BOPDS is protected;
    --extras 
    myExtPaves     :  ListOfPave from BOPDS is protected; 
    --common block 
    myCommonBlock  :  CommonBlock from BOPDS is protected; 
    --shrunk data  
    myTS1          :  Real from Standard is protected;     
    myTS2          :  Real from Standard is protected;   
    myShrunkBox    :  Box   from Bnd is protected;  
    --dummies
    myMFence       :  MapOfInteger from BOPCol is protected;   
 
end PaveBlock;

