-- Created by: DAUTRY Philippe
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

--      	----------------------------

---Version:	0.0
--Version	Date		Purpose
--		0.0	Aug 27 1997	Creation


class XLinkIterator from TDocStd 

	---Purpose: Iterates on Reference attributes.
  --          This is an iterator giving all the external references
  --          of a Document.

uses Document from TDocStd,
     XLink     from TDocStd,
     XLinkPtr  from TDocStd

raises

    NoMoreObject from Standard

is

    Create
    returns XLinkIterator from TDocStd;
	---Purpose: Returns an empty iterator;

    Create (D : Document from TDocStd)
    returns XLinkIterator from TDocStd;
    	---Purpose: Creates an iterator on Reference of <D>.
    
    Initialize (me  : in out; D : Document from TDocStd);
    	---Purpose: Restarts an iteration with <D>.
    
    More (me) returns Boolean;
	---Purpose: Returns True if there is a current Item in the
	--          iteration.
	--          
	---C++: inline
    
    Next (me : in out)
    	raises NoMoreObject from Standard;
    	---Purpose: Move to the next item; raises if there is no more item.
    
    Value (me) returns XLinkPtr from TDocStd;
	---Purpose: Returns the current item; a null handle if there is none.
	--          
	---C++: inline

    Init (me : in out; D : Document from TDocStd) is private;


fields

    myValue : XLinkPtr from TDocStd;

end XLinkIterator;
