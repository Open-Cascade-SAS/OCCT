-- Created on: 1993-07-06
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class CurveOnSurface from PBRep inherits GCurve from PBRep

	---Purpose: Representation  of a  curve   by a   curve  in the
	--          parametric space of a surface.

uses
    Curve    from PGeom2d,
    Surface  from PGeom,
    Pnt2d    from gp,
    Location from PTopLoc

is

    Create(PC : Curve    from PGeom2d;
    	   CF : Real     from Standard;
	   CL : Real     from Standard;
    	   S  : Surface  from PGeom; 
    	   L  : Location from PTopLoc)
    returns mutable CurveOnSurface from PBRep;
    	---Purpose: CF is curve first parameter
    	--          CL is curve last parameter
    	--          As far as they can't be computed from a Persistent Curve
    	--          they are given in the CurveOnSurface constructor

    Surface(me) returns  Surface from PGeom
    is static;
    	---Level: Internal 

    PCurve(me) returns  Curve from PGeom2d
    is static;
    	---Level: Internal 

    IsCurveOnSurface(me) returns Boolean
	---Purpose: Returns True.
    is redefined;
    
    SetUVPoints(me : mutable; Pnt1, Pnt2 : Pnt2d from gp);
    
    FirstUV(me) returns Pnt2d from gp;

    LastUV(me) returns Pnt2d from gp;
    
fields
    
    myPCurve      : Curve   from PGeom2d;
    mySurface     : Surface from PGeom;
    myUV1         : Pnt2d   from gp;
    myUV2         : Pnt2d   from gp;
    
end CurveOnSurface;
