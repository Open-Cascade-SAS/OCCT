-- File:	IGESAppli_ToolLineWidening.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolLineWidening  from IGESAppli

    ---Purpose : Tool to work on a LineWidening. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses LineWidening from IGESAppli,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolLineWidening;
    ---Purpose : Returns a ToolLineWidening, ready to work


    ReadOwnParams (me; ent : mutable LineWidening;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : LineWidening;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : LineWidening;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a LineWidening <ent>, from
    --           its specific (own) parameters

    OwnCorrect (me; ent : mutable LineWidening) returns Boolean  is static;
    ---Purpose : Sets automatic unambiguous Correction on a LineWidening
    --           (NbPropertyValues forced to 5, Level cleared if Subordinate != 0)

    DirChecker (me; ent : LineWidening) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : LineWidening;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : LineWidening; entto : mutable LineWidening;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : LineWidening;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolLineWidening;
