-- Created on: 2000-05-24
-- Created by: data exchange team
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class EdgeDivide from ShapeUpgrade inherits Tool from ShapeUpgrade

	---Purpose: 

uses

    Edge from TopoDS,
    Face from TopoDS,
    HSequenceOfReal from TColStd,
    SplitCurve3d from ShapeUpgrade,
    SplitCurve2d from ShapeUpgrade

is

    Create returns EdgeDivide from ShapeUpgrade;
    	---Purpose: Empty constructor
    
    Clear (me: mutable);
    
    SetFace(me: mutable; F: Face from TopoDS);
    	---C++: inline
    	---Purpose: Sets supporting surface by face
    
    Compute(me: mutable; E: Edge from TopoDS) 
    returns Boolean is virtual;
    
    HasCurve2d(me) returns Boolean;
    	---C++: inline
    
    HasCurve3d(me) returns Boolean;
    	---C++: inline
    
    Knots2d(me) returns HSequenceOfReal from TColStd;
    	---C++: inline
    
    Knots3d(me) returns HSequenceOfReal from TColStd;
    	---C++: inline
    
    SetSplitCurve2dTool(me: mutable; splitCurve2dTool: SplitCurve2d from ShapeUpgrade);
    	---Purpose: Sets the tool for splitting pcurves.
    
    SetSplitCurve3dTool(me: mutable; splitCurve3dTool: SplitCurve3d from ShapeUpgrade);
    	---Purpose: Sets the tool for splitting 3D curves.
    
    GetSplitCurve2dTool(me) returns SplitCurve2d from ShapeUpgrade
    is virtual;
    	---Purpose: Returns the tool for splitting pcurves.
    
    GetSplitCurve3dTool(me) returns SplitCurve3d from ShapeUpgrade
    is virtual;
    	---Purpose: Returns the tool for splitting 3D curves.
	---Remark: here TopoDS_Edge can be used to transfer some specific information (tolerance, etc)
    
fields

    myFace      : Face from TopoDS is protected;
    myHasCurve2d: Boolean is protected;
    myHasCurve3d: Boolean is protected;
    myKnots2d   : HSequenceOfReal from TColStd is protected;
    myKnots3d   : HSequenceOfReal from TColStd is protected;
    
    mySplitCurve3dTool: SplitCurve3d from ShapeUpgrade;
    mySplitCurve2dTool: SplitCurve2d from ShapeUpgrade;

end EdgeDivide;
