-- Created on: 1998-07-28
-- Created by: LECLERE Florence
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class FuseFace from TopOpeBRepBuild

	---Purpose: 

uses Shape                     from TopoDS,
     Face                      from TopoDS,
     Edge                      from TopoDS,
     Vertex                    from TopoDS,
     DataMapOfShapeListOfShape from TopTools,
     ListOfShape               from TopTools


is


    Create
    	returns FuseFace from TopOpeBRepBuild;
    	---C++: inline
    	--   
	
	
    Create(LIF : ListOfShape from TopTools;
   	   LRF : ListOfShape from TopTools;     
	   CXM : Integer from Standard)
	   
    	---C++: inline
    	--      
    	returns FuseFace from TopOpeBRepBuild;


    Init(me: in out; LIF : ListOfShape from TopTools;
	       	     LRF : ListOfShape from TopTools;
	    	     CXM : Integer from Standard)    
    	is static;


    PerformFace(me: in out)
  
    	is static;


    PerformEdge(me: in out)
  
    	is static;

    ClearEdge(me: in out)
    
    	is static;
	
    ClearVertex(me: in out)
    
    	is static;
	
    IsDone(me)
    
    	returns Boolean from Standard
	---C++: inline
	is static;	
	
    IsModified(me)
    
    	returns Boolean from Standard
	---C++: inline
	is static;	
	    
    LFuseFace(me)
    
        returns ListOfShape from TopTools
	---C++: return const&
    	is static;

    LInternEdge(me)
    
        returns ListOfShape from TopTools
	---C++: return const&
    	is static;
	
    LExternEdge(me)
    
        returns ListOfShape from TopTools
	---C++: return const&
    	is static;
	
    LModifEdge(me)
    
        returns ListOfShape from TopTools
	---C++: return const&
    	is static;
	
    LInternVertex(me)
    
        returns ListOfShape from TopTools
	---C++: return const&
    	is static;
	
    LExternVertex(me)
    
        returns ListOfShape from TopTools
	---C++: return const&
    	is static;
	
    LModifVertex(me)
    
        returns ListOfShape from TopTools
	---C++: return const&
    	is static;
	
		
fields

    myLIF      : ListOfShape               from TopTools;
    myLRF      : ListOfShape               from TopTools;
    myLFF      : ListOfShape               from TopTools;
    
    myLIE      : ListOfShape               from TopTools is protected;
    myLEE      : ListOfShape               from TopTools is protected;
    myLME      : ListOfShape               from TopTools is protected;
        
    myLIV      : ListOfShape               from TopTools is protected;
    myLEV      : ListOfShape               from TopTools is protected;
    myLMV      : ListOfShape               from TopTools is protected;

    myInternal : Boolean                   from Standard; 
    myModified : Boolean                   from Standard;
    myDone     : Boolean                   from Standard;
    
end FuseFace;    
