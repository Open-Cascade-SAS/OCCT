-- File:	RWStepRepr_RWMeasureRepresentationItem.cdl
-- Created:	Wed Sep  8 11:41:18 1999
-- Author:	Andrey BETENEV
--		<abv@doomox.nnov.matra-dtv.fr>
---Copyright:	 Matra Datavision 1999


class RWMeasureRepresentationItem from RWStepRepr 

	---Purpose : Read & Write Module for MeasureRepresentationItem

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     MeasureRepresentationItem from StepRepr,
     EntityIterator from Interface

is

    Create returns RWMeasureRepresentationItem;

    ReadStep (me; data : StepReaderData; num : Integer;
	          ach : in out Check; ent : mutable MeasureRepresentationItem from StepRepr);

    WriteStep (me; SW : in out StepWriter; ent : MeasureRepresentationItem from StepRepr);

    Share(me; ent : MeasureRepresentationItem from StepRepr; iter : in out EntityIterator from Interface);

end RWMeasureRepresentationItem;
