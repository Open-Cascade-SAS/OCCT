-- Created on: 2005-01-21
-- Created by: Alexander SOLOVYOV
-- Copyright (c) 2005-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class DataSource3D from MeshVS inherits DataSource from MeshVS

uses
  Integer                             from Standard,
  Array1OfPnt                         from TColgp,

  HArray1OfSequenceOfInteger          from MeshVS,
  DataMapOfHArray1OfSequenceOfInteger from MeshVS

is

  GetPrismTopology  ( me; BasePoints : Integer ) returns HArray1OfSequenceOfInteger from MeshVS;
  GetPyramidTopology( me; BasePoints : Integer ) returns HArray1OfSequenceOfInteger from MeshVS;

  CreatePrismTopology  ( myclass; BasePoints : Integer ) returns HArray1OfSequenceOfInteger from MeshVS;
  CreatePyramidTopology( myclass; BasePoints : Integer ) returns HArray1OfSequenceOfInteger from MeshVS;

fields
  myPrismTopos, myPyramidTopos : DataMapOfHArray1OfSequenceOfInteger from MeshVS;

end DataSource3D from MeshVS;
