-- Created on: 1994-04-01
-- Created by: Yves FRICAUD
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class PolyBis from Bisector 

	---Purpose: Polygon of PointOnBis

uses
    PointOnBis from Bisector,
    Trsf2d     from gp

is
    Create returns PolyBis from Bisector;
    
    Append ( me : in out; Point : PointOnBis from Bisector) 
    is static ;
						    		
    Length (me) returns Integer
    is static ;
    
    IsEmpty (me) returns Boolean
    is static;

    Value (me ; Index : Integer) returns PointOnBis from Bisector
       ---C++: return const&
    is static;
    
    First (me) returns PointOnBis from Bisector
       ---C++: return const&
    is static;
    
    Last (me) returns PointOnBis from Bisector
       ---C++: return const&
    is static;
    
    Interval (me ; U :Real) returns Integer from Standard
    is static;
    
    Transform (me : in out ; T :Trsf2d)
    is static;
    
fields

    thePoints       : PointOnBis from Bisector [30];
    nbPoints        : Integer    from Standard;
    
end PolyBis;

