-- Created on: 2004-06-15
-- Created by: Sergey ZARITCHNY <szy@opencascade.com>
-- Copyright (c) 2004-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class LocationSet from BinTools 

	---Purpose: The class LocationSet stores a set of location in
	--          a relocatable state.
	--          
	--          It can be created from Locations.
	--          
	--          It can create Locations.


uses
    Location             from TopLoc,
    IndexedMapOfLocation from TopLoc

raises
    OutOfRange           from Standard

is
    Create returns LocationSet from BinTools;
	---Purpose: Returns an empty set of locations.
	
    Clear(me : in out)
	---Purpose: Clears the content of the set.
    is static;
	
    Add(me : in out; L : Location from TopLoc) returns Integer
	---Purpose: Incorporate a new Location in the  set and returns
	--          its index.
    is static;
    
    Location(me; I : Integer) returns Location from TopLoc
	---Purpose: Returns the location of index <I>.
	--          
	---C++: return const &
    raises
    	OutOfRange from Standard
    is static;

    Index(me; L : Location from TopLoc) returns Integer
	---Purpose: Returns the index of <L>.
    is static; 
     
    NbLocations(me) returns Integer
	---Purpose: Returns number of locations.
    is static; 
    	
    Write(me; OS : in out OStream)
	---Purpose: Writes the content of  me  on the stream <OS> in a
	--          format that can be read back by Read.
    is static;
	
    Read(me : in out; IS : in out IStream)
	---Purpose: Reads the content of me from the  stream  <IS>. me
	--          is first cleared.
	--          
    is static;
	
fields
 
    myMap : IndexedMapOfLocation from TopLoc;

end LocationSet;

