-- Created on: 1995-03-08
-- Created by: Bruno DUMORTIER
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MakeHalfSpace from BRepPrimAPI  inherits MakeShape from BRepBuilderAPI

	---Purpose: Describes functions to build half-spaces.
    	-- A half-space is an infinite solid, limited by a surface. It
    	-- is built from a face or a shell, which bounds it, and with
    	-- a reference point, which specifies the side of the
    	-- surface where the matter of the half-space is located.
    	-- A half-space is a tool commonly used in topological
    	-- operations to cut another shape.
    	-- A MakeHalfSpace object provides a framework for:
    	-- -   defining and implementing the construction of a half-space, and
    	-- -   consulting the result.

uses
    Shape      from TopoDS,
    Vertex     from TopoDS,
    Face       from TopoDS,
    Shell      from TopoDS,
    Solid      from TopoDS,
    Pnt        from gp, 
    MakeShape from BRepBuilderAPI

raises
    NotDone from StdFail
is

    Create(Face   : Face from TopoDS;
    	   RefPnt : Pnt  from gp)
    returns MakeHalfSpace from BRepPrimAPI;
	---Purpose: Make a HalfSpace defined with a Face and a Point.
	---Level: Public

    Create(Shell  : Shell from TopoDS;
    	   RefPnt : Pnt   from gp)
    returns MakeHalfSpace from BRepPrimAPI;
	---Purpose: Make a HalfSpace defined with a Shell and a Point.
	---Level: Public


    ----------------------------------------------
    -- Results
    ----------------------------------------------

    Solid(me) returns Solid from TopoDS
	---Purpose: Returns the constructed half-space as a solid.
    	---C++: return const &
	---C++: alias "Standard_EXPORT operator TopoDS_Solid() const;" 
    raises
    	NotDone from StdFail
    is static; 

fields

    mySolid : Solid from TopoDS;

end MakeHalfSpace;
