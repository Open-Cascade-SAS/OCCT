-- Created on: 1993-01-04
-- Created by: J.P. BOUDIER - J.P. TIRAULT
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Date from Quantity 

inherits Storable from Standard 

    	---Purpose: This class provides services to manage date information.
    	--          A date represents the following time intervals:
    	-- year, month, day, hour, minute, second,
    	-- millisecond and microsecond.
    	-- Current time is expressed in elapsed seconds
    	-- and microseconds beginning from 00:00 GMT,
    	-- January 1, 1979 (zero hour). The valid date can
    	-- only be later than this one.
    	-- Note: a Period object gives the interval between two dates.


uses Period


raises DateDefinitionError from Quantity , OutOfRange from Standard

is
   
  Create returns Date;
    	---Purpose:  Constructs a default date
    	-- (00:00 GMT, January 1, 1979 (zero hour)); use the function
    	--   SetValues to define the required date; or

  Create ( mm, dd, yyyy, hh, mn, ss : Integer ; mis , mics : Integer = 0)
          returns Date
    	---Purpose:   Constructs a date from the year yyyy, the
    	-- month mm, the day dd, the hour hh, the minute
    	-- mn, the second ss, the millisecond mis
    	-- (defaulted to 0) and the microsecond mics (defaulted to 0)..
    	--          With:      1 <= mm <= 12
    	--                     1 <= dd <= max number of days of <mm>
    	--                     1979 <= yyyy
    	--                     0 <= hh <= 23
    	--                     0 <= mn <= 59
    	--                     0 <= ss <= 59
    	--                     0 <= mis <= 999
    	--                     0 <= mics <= 999 
    	-- Exceptions
    	-- Quantity_DateDefinitionError if mm, dd, hh,
    	-- mn, ss, mis and mics are not the components of the valid date.
    raises DateDefinitionError;

  Values (me ; mm, dd, yy, hh, mn, ss, mis, mics : out Integer)  is static;
    	---Purpose: Gets a complete Date.
    	-- -   in mm - the month,
    	-- -   in dd - the day,
    	-- -   in yyyy - the year,
    	-- -   in hh - the hour,
    	-- -   in mn - the minute,
    	-- -   in ss - the second,
    	-- -   in mis - the millisecond, and
    	-- -   in mics - the microsecond
  SetValues (me : out; mm, dd, yy, hh, mn, ss : Integer; 
             mis, mics : Integer = 0)
    	---Purpose: Assigns to this date the year yyyy, the month
    	-- mm, the day dd, the hour hh, the minute mn, the
    	-- second ss, the millisecond mis (defaulted to 0)
    	-- and the microsecond mics (defaulted to 0).
    	-- Exceptions
    	-- Quantity_DateDefinitionError if mm, dd, hh,
    	-- mn, ss, mis and mics are not components of a valid date.
    raises DateDefinitionError is static;

  Difference (me  : out; anOther : Date) returns Period is static;
    	---Purpose: Subtracts one Date from another one to find the period
    	--          between and returns the value.
    	--          The result is the absolute value between the difference
    	--          of two dates.

  Subtract (me  : out; aPeriod : Period) returns Date 
    	---Purpose: Subtracts a period from a Date and returns the new Date.
    	--          Raises an exception if the result date is anterior to
    	--          Jan 1, 1979.
    	---C++: alias operator -
  raises OutOfRange is static;

  Add(me  : out; aPeriod : Period) returns Date is static;
    	---Purpose: Adds a Period to a Date and returns the new Date.
    	---C++: alias operator +

  Year (me : out) returns Integer is static;
    	---Purpose: Returns year of a Date.

  Month (me : out) returns Integer is static;
    	---Purpose: Returns month of a Date.

  Day (me : out) returns Integer is static;
    	---Purpose: Returns Day of a Date.

  Hour (me : out) returns Integer is static;
    	---Purpose: Returns Hour of a Date.

  Minute (me : out) returns Integer is static;
    	---Purpose: Returns minute of a Date.

  Second (me : out) returns Integer is static;
    	---Purpose: Returns seconde of a Date.

  MilliSecond (me : out) returns Integer is static;
    	---Purpose: Returns millisecond of a Date.

  MicroSecond (me : out) returns Integer is static;
    	---Purpose: Returns microsecond of a Date.

  IsEqual (me ; anOther : Date) returns Boolean is static;
      	---Purpose: Returns TRUE if both <me> and <other> are equal.
      	-- This method is an alias of operator ==.
      	---C++: alias operator ==
  

  IsEarlier (me ; anOther : Date) returns Boolean is static;
     	---Purpose: Returns TRUE if <me> is earlier than <other>.
     	---C++: alias operator <

  IsLater (me ; anOther : Date) returns Boolean is static;
     	---Purpose: Returns TRUE if <me> is later then <other>.
     	---C++: alias operator >
  
  IsValid (myclass ; mm, dd, yy, hh, mn, ss : Integer; 
             mis, mics : Integer = 0) returns Boolean;
	---Purpose: Checks the validity of a date - returns true if a
    	-- date defined from the year yyyy, the month mm,
    	-- the day dd, the hour hh, the minute mn, the
    	-- second ss, the millisecond mis (defaulted to 0)
    	-- and the microsecond mics (defaulted to 0) is valid.
    	-- A date must satisfy the conditions above:
    	-- -   yyyy is greater than or equal to 1979,
    	-- -   mm lies within the range [1, 12] (with 1
    	--   corresponding to January and 12 to December),
    	-- -   dd lies within a valid range for the month mm
    	--   (from 1 to 28, 29, 30 or 31 depending on
    	--   mm and whether yyyy is a leap year or not),
    	-- -   hh lies within the range [0, 23],
    	-- -   mn lies within the range [0, 59],
    	-- -   ss lies within the range [0, 59],
    	-- -   mis lies within the range [0, 999],
    	-- -   mics lies within the range [0, 999].C
    
  IsLeap (myclass  ; yy : Integer ) returns Boolean;
    	---Purpose: Returns true if a year is a leap year.
    	--          The leap years are divisable by 4 and not by 100 except 
    	--          the years divisable by 400.
    	---C++: inline

 fields
  mySec  : Integer;
  myUSec : Integer;
end Date from Quantity;

