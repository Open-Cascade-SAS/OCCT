-- Created on: 1998-02-02
-- Created by: Philippe MANGIN
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



private  class LocFunction from GeomFill 

	---Purpose: 

uses 
 LocationLaw from GeomFill,
 Array1OfVec   from TColgp, 
 Mat  from  gp

is 
    Create( Law  :  LocationLaw  from  GeomFill) 
    returns  LocFunction  from  GeomFill; 
     
    
   D0(me : in  out; 
      Param: Real;
      First, Last : Real)
      ---Purpose: compute the section for v = param           
   returns Boolean; 
	
   D1(me : in  out;
      Param: Real;
      First, Last : Real)
      ---Purpose: compute the first  derivative in v direction  of the
      --           section for v =  param 
   returns Boolean;
   
    D2(me : in  out;
      Param: Real;
      First, Last : Real)      
      ---Purpose: compute the second derivative  in v direction of the
      --          section  for v = param  
   returns Boolean; 
    
   DN(me  :  in  out;
      Param       : Real;
      First, Last : Real; 
      Order       :  Integer; 
      Result      :  in  out  Real; 
      Ier         :  out  Integer); 

fields 
  myLaw  :  LocationLaw  from  GeomFill;
  V,  DV,  D2V  :  Array1OfVec  from  TColgp; 
  M,  DM,  D2M  :  Mat  from  gp;
end LocFunction;
