-- Created on: 1991-01-08
-- Created by: Didier Piffault
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

--- Modified by  hl1 (juillet 96) : ajout de SeqOfBox




--------------------------------------------------------
---              I n f o r m a t i o n               ---
---                                                  ---
---  The Bnd_Tool class is now in the package Intf.  ---
--------------------------------------------------------





package Bnd 

        ---Purpose: Supports the Boundings Volumes.  A Bounding Volume
        --          is used to bound a shape to optimising algorithms.
        --          If  a point is  outside the Bounding   Volume of a
        --          shape it is also  outside the shape.  The contrary
        --          is not necessarily true.
        --          
        --          Various classes are  then implemented to  describe
        --          the usual  Bounding volumes. Not  all  classes are
        --          implemented.
        --          
        --          in 3D :
        --          Box                -- Implemented
        --          BoundSortBox       -- Implemented
        --          
        --          in 2D :
        --          Box2d              -- Implemented
        --          BoundSortBox2d     -- Implemented
        --          
        --          

        ---Level : Public. 
        --  All methods of all  classes will be public.

        
uses    Standard,
        TCollection,
        TColStd,
        gp,
	MMgt


is  class Box;
    class Array1OfBox instantiates Array1 from TCollection
                                   (Box from Bnd);
    class HArray1OfBox instantiates HArray1 from TCollection
                                   (Box from Bnd,
                                    Array1OfBox from Bnd);

   class Sphere;
   class Array1OfSphere instantiates Array1 from TCollection
   	 			     (Sphere from Bnd);
   class HArray1OfSphere instantiates HArray1 from TCollection
   	 		 	      (Sphere from Bnd,
				      Array1OfSphere from Bnd);


    class Box2d;
    class Array1OfBox2d instantiates Array1 from TCollection
                                   (Box2d from Bnd);
    class HArray1OfBox2d instantiates HArray1 from TCollection
                                   (Box2d from Bnd,
                                    Array1OfBox2d from Bnd);


    class BoundSortBox2d;
    class BoundSortBox;
    class SeqOfBox instantiates Sequence from TCollection (Box from Bnd);
        ---Purpose: This sequence used to store the bounding boxes of sub-Shapes.
    
    --- Optimized boxes (no Gap, no infinity supported)
    generic class B2x;
    generic class B3x;

    class B2d instantiates B2x from Bnd (Real from Standard);
    -- 2D box with double-precision coordinates

    class B2f instantiates B2x from Bnd (ShortReal from Standard);
    -- 2D box with single-precision coordinates

    class B3d instantiates B3x from Bnd (Real from Standard);
    -- 3D box with double-precision coordinates

    class B3f instantiates B3x from Bnd (ShortReal from Standard);
    -- 3D box with single-precision coordinates

end Bnd;
