-- File:	TCompSolid.cdl
-- Created:	Mon Dec 17 11:18:44 1990
-- Author:	Remi Lequette
--		<rle@topsn3>
---Copyright:	 Matra Datavision 1990, 1992



class TCompSolid from PTopoDS inherits TShape from PTopoDS

	---Purpose: A  topological Composite  Solid shape.

uses
    ShapeEnum from TopAbs

is
    Create returns mutable TCompSolid from PTopoDS;
	---Purpose: The new  TCompSolid is empty.
    ---Level: Internal 
    	
    ShapeType(me) returns ShapeEnum from TopAbs;
    ---Level: Internal 

end TCompSolid;
