-- File:	IGESAppli_ToolElementResults.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolElementResults  from IGESAppli

    ---Purpose : Tool to work on a ElementResults. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses ElementResults from IGESAppli,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolElementResults;
    ---Purpose : Returns a ToolElementResults, ready to work


    ReadOwnParams (me; ent : mutable ElementResults;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : ElementResults;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : ElementResults;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a ElementResults <ent>, from
    --           its specific (own) parameters

    DirChecker (me; ent : ElementResults) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : ElementResults;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : ElementResults; entto : mutable ElementResults;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : ElementResults;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolElementResults;
