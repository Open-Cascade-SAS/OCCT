-- Created on: 1993-07-21
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.





deferred class Command from BRepLib 

	---Purpose: Root class for all commands in BRepLib.  
	--          
	--          Provides :
	--          
	--          * Managements of the notDone flag.
	--          
	--          * Catching of exceptions (not implemented).
	--          
	--          * Logging (not implemented).

raises
    NotDone from StdFail
    
is
    Delete(me:out) is virtual;
    ---C++: alias "Standard_EXPORT virtual ~BRepLib_Command(){Delete() ; }"
    
    Initialize;
	---Purpose: Set done to False.
    
    IsDone(me) returns Boolean
	---Level: Public
    is static;
    
    Done(me : in out)
	---Purpose: Set done to true.
	---Level: Public
    is static protected;
    
    NotDone(me : in out)
	---Purpose: Set done to false.
	---Level: Public
    is static protected;
    
    
    
    Check(me)
	---Purpose: Raises NotDone if done is false.
	---Level: Public
    raises NotDone from StdFail
    is static;

fields 
    myDone : Boolean;

end Command;
