-- Created on: 1994-05-26
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SolidSurfaceInterference from TopOpeBRepDS 
    inherits Interference from TopOpeBRepDS

	---Purpose: 

uses

    Transition  from TopOpeBRepDS,
    Kind        from TopOpeBRepDS,
    OStream     from Standard    
    
is

    Create(Transition   : Transition from TopOpeBRepDS;
	   SupportType  : Kind from TopOpeBRepDS;
	   Support      : Integer;
	   GeometryType : Kind from TopOpeBRepDS;
	   Geometry     : Integer)
    returns SolidSurfaceInterference from TopOpeBRepDS;

    Dump(me; OS : in out OStream from Standard) returns OStream
    is redefined;
    ---C++: return &

end SolidSurfaceInterference from TopOpeBRepDS;
