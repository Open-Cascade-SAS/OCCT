-- Created on: 1993-07-27
-- Created by: Jean Louis FRENKEL
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class PixelInterpolation from Image

	---Purpose: The class PixelInterpolation is used to compute a Pixel 
	--            value on non-integer Image coordinate. This Pixel type
	--	      is called SubPixel .
	--          PixelInterpolation is the default and is the simplest one,
	--	      SubPixel value on non-integer Image coordinate is the 
	--	      value of the nearest Pixel at integer coordinate.
	--	    The user can create a new kind of PixelInterpolation with a
	--	      new algorithm by creating a new derived PixelInterpolation
	--	      class and redefined Interpolate() method.
	--	    If V1  is the value of the nearest Image Pixel
	--		V = V1 is the Image SubPixel value on non-integer 
	--	      coordinate (FX,FY)

uses

    Pixel       	from Aspect,
    Image	    	from Image,
    ColorPixel       	from Aspect,
    IndexPixel       	from Aspect,
    DColorImage 	from Image,
    DIndexedImage 	from Image

is

    	Create returns PixelInterpolation from Image ;
	---Level: Public
    	---Purpose: Create a PixelInterpolation  object.

	Interpolate( me ; aImage   : Image from Image ;
		          X,Y      : Real  from Standard ;
			  LowerX,LowerY,UpperX,UpperY : Integer from Standard ;
		          RetPixel : in out Pixel from Aspect ) 
		returns Boolean from Standard
		is virtual ;
	---Level: Public
    	---Purpose: Compute SubPixel's value on non-integer Image coordinate.
	--	    LowerX,LowerY,UpperX,UpperY is the Image Min Max, it's used
	--	    to check if the SubPixel coordinate X,Y is outside of image.
	--          Return True  if Interpolation Succes.
	--	    Retrun False if the SubPixel is out from Image.

	Interpolate( me ; aImage   : DColorImage from Image ;
		          FX,FY      : Real  from Standard ;
			  LowerX,LowerY,UpperX,UpperY : Integer from Standard ;
		          RetPixel : in out ColorPixel from Aspect ) 
		returns Boolean from Standard
		is virtual ;
	---Level: Public
    	---Purpose: Compute SubPixel's value on non-integer Image coordinate for
	--	      DColorImage and ColorPixel.
	--	    LowerX,LowerY,UpperX,UpperY is the Image Min Max, it's used
	--	      to check if the SubPixel coordinate FX,FY is outside of 
	--	      image.
	--          Return True  if Interpolation Succes.
	--	    Return False if the SubPixel is out from Image.


	Interpolate( me ; aImage   : DIndexedImage from Image ;
		          FX,FY      : Real  from Standard ;
			  LowerX,LowerY,UpperX,UpperY : Integer from Standard ;
		          RetPixel : in out IndexPixel from Aspect ) 
		returns Boolean from Standard
		is virtual ;
	---Level: Public
    	---Purpose: Compute SubPixel's value on non-integer Image coordinate for
	--	      DIndexedImage and IndexPixel.
	--	    LowerX,LowerY,UpperX,UpperY is the Image Min Max, it's use
	--	    check if the SubPixel coordinate X,Y is outside of image.
	--          Return True  if Interpolation Succes.
	--	    Return False if the SubPixel is out from Image.

	DoInterpolate( me ; aImage   : Image from Image ;
		            X,Y      : Real  from Standard ;
			    LowerX,LowerY,UpperX,UpperY: Integer from Standard ;
		            RetPixel : in out Pixel from Aspect ) 
		returns Boolean from Standard is static private ;

end PixelInterpolation from Image;
