-- Created on: 1997-04-14
-- Created by: Christian CAILLET
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class SelectBasicGeom  from IGESSelect  inherits SelectExplore

    ---Purpose : This selection returns the basic geometric elements
    --           contained in an IGES Entity
    --           Intended to run a "quick" transfer. I.E. :
    --           - for a Group, considers its Elements
    --           - for a Trimmed or Bounded Surface or a Face (BREP),
    --             considers the 3D curves of each of its loops
    --           - for a Plane (108), considers its Bounding Curve
    --           - for a Curve itself, takes it
    --           
    --           Also, FREE surfaces are taken, because curve 3d is known for
    --           them. (the ideal should be to have their natural bounds)
    --           
    --           If <curvesonly> is set, ONLY curves-3d are returned

uses AsciiString from TCollection, Transient, EntityIterator, Graph,
     IGESEntity from IGESData

is

    Create (mode : Integer) returns mutable SelectBasicGeom;
    ---Purpose : Creates a SelectBasicGeom, which allways works recursively
    --           mode = -1 : Returns Surfaces (without trimming)
    --           mode = +1 : Returns Curves 3D (free or bound of surface)
    --           mode = +2 : Returns Basic Curves 3D : as 1 but CompositeCurves
    --                        are returned in detail
    --           mode = 0  : both

    CurvesOnly (me) returns Boolean;

    Explore (me; level : Integer; ent : Transient; G : Graph;
    	     explored : in out EntityIterator)
    	returns Boolean;
    ---Purpose : Explores an entity, to take its contained Curves 3d
    --           Works recursively


    ExploreLabel (me) returns AsciiString from TCollection;
    ---Purpose : Returns a text defining the criterium : "Curves 3d" or
    --           "Basic Geometry"

    SubCurves (myclass; ent : IGESEntity; explored : in out EntityIterator)
    	returns Boolean;
    ---Purpose : This method can be called from everywhere to get the curves
    --           as sub-elements of a given curve :
    --           CompositeCurve : explored lists its subs + returns True
    --           Any Curve : explored is not filled but returned is True
    --           Other : returned is False

fields

    thegeom : Integer;  -- -1 : Surfaces only  1 : Curves 3D only  0 : both

end SelectBasicGeom;
