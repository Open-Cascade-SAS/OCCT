-- Created on: 1992-08-28
-- Created by: Remi LEQUETTE
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



package GeomTools 

	---Purpose: The GeomTools package provides  utilities for Geometry.
	--          
	--          *  SurfaceSet,  CurveSet, Curve2dSet  : Tools used
	--          for dumping, writing and reading.
	--          
	--          * Methods to dump, write, read curves and surfaces.

uses
    Geom,
    Geom2d,
    TColStd,
    Message

is

    class UndefinedTypeHandler;
    --
    --  Dump, Write, Read tools
    
    class SurfaceSet;
	---Purpose: A set of Surfaces from Geom.
    	
    class CurveSet;
	---Purpose: A set of Curves from Geom.
    	
    class Curve2dSet;
	---Purpose: A set of Curves from Geom2d.
    	
    --
    --     Methods
    --     
    
    Dump(S : Surface from Geom; OS : in out OStream);
	  ---Purpose: Dumps the surface on the stream.

    Write(S : Surface from Geom; OS : in out OStream);
	  ---Purpose: Writes the surface on the stream.

    Read(S : in out Surface from Geom; IS : in out IStream); 
	  ---Purpose: Reads the surface from the stream.


    Dump(C : Curve from Geom; OS : in out OStream);
	  ---Purpose: Dumps the Curve on the stream.

    Write(C : Curve from Geom; OS : in out OStream);
	  ---Purpose: Writes the Curve on the stream.

    Read(C : in out Curve from Geom; IS : in out IStream); 
	  ---Purpose: Reads the Curve from the stream.


    Dump(C : Curve from Geom2d; OS : in out OStream);
	  ---Purpose: Dumps the Curve on the stream.

    Write(C : Curve from Geom2d; OS : in out OStream);
	  ---Purpose: Writes the Curve on the stream.

    Read(C : in out Curve from Geom2d; IS : in out IStream); 
	  ---Purpose: Reads the Curve from the stream.
	  
    SetUndefinedTypeHandler(aHandler: UndefinedTypeHandler from GeomTools);
    
    GetUndefinedTypeHandler returns UndefinedTypeHandler from GeomTools;

end GeomTools;


