-- Created on: 1997-12-10
-- Created by: Denis PASCAL
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class Relation from TDataStd inherits Attribute from TDF
    
    ---Purpose: Relation attribute. 
    --          ==================
    --
    --            *  Data Structure of  the  Expression is stored in a
    --           string and references to variables used by the string
    --
    --  Warning:  To be consistent,  each  Variable  referenced by  the
    --          relation must have its equivalent in the string


uses Attribute       from TDF,
     Label           from TDF,
     GUID            from Standard,
     Real            from Standard,
     DataSet         from TDF,
     RelocationTable from TDF,
     ExtendedString  from TCollection,
     AttributeList   from TDF
     

is

    ---Purpose: class methods
    --          =============

    GetID (myclass)    
    	---C++: return const & 
    returns GUID from Standard;
    

    Set (myclass ; label : Label from TDF)
    ---Purpose: Find, or create, an Relation attribute.
    returns Relation from TDataStd;
    
    ---Purpose: Real methods
    --          ============

    Create
    returns mutable Relation from TDataStd;
    
    Name (me)
    ---Purpose: build and return the relation name
    returns ExtendedString from TCollection;
    
    SetRelation (me : mutable; E : ExtendedString from TCollection);
    
    GetRelation (me)
    returns ExtendedString from TCollection; 
    ---C++: return const &
    
    GetVariables (me : mutable)
    ---C++: return &
    returns AttributeList from TDF;    
    
    ---Category: TDF_Attribute methods
    --           =====================
    
    ID (me) 
    ---C++: return const &  
    returns GUID from Standard;

    Restore (me: mutable; With : Attribute from TDF);

    NewEmpty(me)
    returns mutable Attribute from TDF;

    Paste (me; Into : mutable Attribute from TDF;
	       RT   : mutable RelocationTable from TDF);    

    Dump(me; anOS : in out OStream from Standard)
    returns OStream from Standard
    is redefined;
    ---C++: return &

fields

    myRelation   : ExtendedString from TCollection;
    myVariables  : AttributeList from TDF;  

end Relation;
