-- Created on: 1992-09-30
-- Created by: Christian CAILLET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class AllShared  from IFGraph  inherits GraphContent

    	---Purpose : this class determines all Entities shared by some specific
    	--           ones, at any level (those which will be lead in a Transfer
    	--           for instance)

uses Transient, EntityIterator, Graph

is

    Create (agraph : Graph) returns AllShared;
    ---Purpose : creates an AllShared from a graph, empty ready to be filled

    Create (agraph : Graph; ent : any Transient)
    	returns AllShared;
    ---Purpose : creates an AllShared which memrizes Entities shared by a given
    --           one, at any level, including itself

    GetFromEntity (me : in out; ent : any Transient);
    ---Purpose : adds an entity and its shared ones to the list (allows to
    --           cumulate all Entities shared by some ones)

    GetFromIter (me : in out; iter : EntityIterator);
    ---Purpose : Adds Entities from an EntityIterator and all their shared
    --           ones at any level

    ResetData (me : in out);
    ---Purpose : Allows to restart on a new data set

    	-- --   Results   -- --
    	--   More-Next-Value give all entities noted as shared,
    	--   including the entities given for construction or to GetFromEntity

    Evaluate (me : in out) is redefined;
    ---Purpose : does the specific evaluation (shared entities atall levels)

fields

    thegraph : Graph;

end AllShared;
