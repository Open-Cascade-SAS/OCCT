-- Created on: 1993-02-19
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package BRepAdaptor 

	---Purpose: The BRepAdaptor package provides classes to access 
	--          the geometry of the BRep models.
	--          
	--          OverView of classes
	--          
	--          * Surface :  Provides the methods  of Surface from
	--          Adpator on a Face.
	--          
	--          *  Curve  : Provides  the  methods of  Curve  from
	--          Adaptor3d on an Edge.
	--          
	--          * Curve2d : Provides  the methods of  Curve2d from
	--          Adaptor2d on an Edge on a Face.
	--          

uses
    gp, 
    TCollection,
    TColgp,
    TColStd,
    GeomAbs,
    Adaptor3d,
    Adaptor2d,
    Geom,
    Geom2d,
    GeomAdaptor,
    Geom2dAdaptor,
    TopoDS,
    BRep

is

    class Surface;
	---Purpose: Transforms a Face in a Surface from Adaptor3d.
	
    class Curve;
	---Purpose: Transforms an Edge in a Curve from Adaptor3d.

    class Curve2d;
	---Purpose: Transforms an Edge   on a Face  in  a Curve2d from
	--          Adaptor2d. 

    class  CompCurve; 
    	---Purpose: Transforms a Wire in a Curve from Adaptor3d.
    	
    class HSurface instantiates GenHSurface from Adaptor3d
    	(Surface from BRepAdaptor);

    class HCurve instantiates GenHCurve from Adaptor3d
    	(Curve from BRepAdaptor);

    class HCurve2d instantiates GenHCurve2d from Adaptor2d
    	(Curve2d from BRepAdaptor); 
	 
    class HCompCurve instantiates GenHCurve from Adaptor3d
    	(CompCurve from BRepAdaptor); 
	 
    class Array1OfCurve 
    	instantiates Array1 from TCollection (Curve from BRepAdaptor); 
	 
    class HArray1OfCurve
    	instantiates HArray1 from TCollection (Curve from BRepAdaptor,
    	    	    	    	Array1OfCurve from BRepAdaptor);

end BRepAdaptor;
