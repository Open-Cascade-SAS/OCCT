-- Created on: 1995-03-27
-- Created by: Christophe MARION
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class FaceData from HLRTopoBRep

	---Purpose: Contains the  3 ListOfShape of  a Face  ( Internal
	--          OutLines, OutLines on restriction and IsoLines ).

uses
    Shape       from TopoDS,
    ListOfShape from TopTools

is
    Create returns FaceData from HLRTopoBRep;

    FaceIntL(me) 
    returns ListOfShape from TopTools
	---C++: inline
	---C++: return const &
    is static;

    FaceOutL(me) 
    returns ListOfShape from TopTools
	---C++: inline
	---C++: return const &
    is static;

    FaceIsoL(me) 
    returns ListOfShape from TopTools
	---C++: inline
	---C++: return const &
    is static;

    AddIntL(me : in out) 
    returns ListOfShape from TopTools
	---C++: inline
	---C++: return &
    is static;

    AddOutL(me : in out) 
    returns ListOfShape from TopTools
	---C++: inline
	---C++: return &
    is static;

    AddIsoL(me : in out) 
    returns ListOfShape from TopTools
	---C++: inline
	---C++: return &
    is static;

fields

    myIntL : ListOfShape from TopTools;
    -- For a face the list of internal OutLines.

    myOutL : ListOfShape from TopTools;
    -- For a face the list of not OutLines on restriction.

    myIsoL : ListOfShape from TopTools;
    -- For a face the list of IsoLines.

end FaceData;
