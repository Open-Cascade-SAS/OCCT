-- Created on: 1998-01-15
-- Created by: Denis PASCAL
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Comment from TDataStd inherits Attribute from TDF

	---Purpose: Comment attribute. may be  associated to any label
	--          to store user comment.

uses Attribute         from TDF,
     Label             from TDF,
     GUID              from Standard,
     ExtendedString    from TCollection,
     DataSet           from TDF,
     RelocationTable   from TDF,
     AttributeSequence from TDF,
     Data              from TDF


is    


    ---Purpose: class methods
    --          =============

    GetID (myclass)   
  	---C++: return const & 
    	---Purpose: Returns the GUID for comments.  
    returns GUID from Standard;    

    Set (myclass; label : Label from TDF)
    ---Purpose:  Find, or create  a   Comment attribute.  the  Comment
    --          attribute is returned.
    returns Comment from TDataStd;    

    Set (myclass; label : Label from TDF; string  : ExtendedString from TCollection)
    ---Purpose: Finds, or creates a Comment attribute and sets the string.
    --          the Comment attribute is returned.
    returns Comment from TDataStd;
    
    ---Purpose: Comment methods
    --          ============
    
    Create 
    returns mutable Comment from TDataStd;
        
    Set (me : mutable; S : ExtendedString from TCollection);

    
    Get (me)
    returns ExtendedString from TCollection;    
    ---Purpose:
    --    Returns the comment attribute.
    ---C++: return const & 

    ---Category: TDF_Attribute methods
    --           =====================
    
    ID (me)
     	---C++: return const & 
    returns GUID from Standard;

    Restore (me: mutable; with : Attribute from TDF);

    NewEmpty (me)
    returns mutable Attribute from TDF;

    Paste (me; into : mutable Attribute from TDF;
	       RT   : mutable RelocationTable from TDF);    

    Dump(me; anOS : in out OStream from Standard)
    	returns OStream from Standard
    	is redefined;
	---C++: return &

    AfterRetrieval(me: mutable;
    	    	   forceIt : Boolean from Standard = Standard_False)
    	returns Boolean from Standard
    	is redefined static;


fields

    myString : ExtendedString from TCollection;

end Comment;
