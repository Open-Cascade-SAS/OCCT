-- Created on: 1993-03-22
-- Created by: Philippe DAUTRY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package PColgp  

        ---Purpose :   This package  provides   some instantiations of
        --         generic classes  from PCollection with objects from gp. 
	 
uses PCollection, gp

is



    -- HArray1 of 2D objects.

  class HArray1OfCirc2d
    instantiates HArray1 from PCollection (Circ2d from gp);
  class HArray1OfDir2d
    	instantiates HArray1 from PCollection (Dir2d from gp);
  class HArray1OfLin2d
    	instantiates HArray1 from PCollection (Lin2d from gp);
  class HArray1OfPnt2d
    	instantiates HArray1 from PCollection (Pnt2d from gp);
  class HArray1OfVec2d
    	instantiates HArray1 from PCollection (Vec2d from gp);
  class HArray1OfXY
    	instantiates HArray1 from PCollection (XY from gp);


    -- HArray1 of 3D objects.

  class HArray1OfDir
    	instantiates HArray1 from PCollection (Dir from gp);
  class HArray1OfPnt
    	instantiates HArray1 from PCollection (Pnt from gp);
  class HArray1OfVec
    	instantiates HArray1 from PCollection (Vec from gp);
  class HArray1OfXYZ
    	instantiates HArray1 from PCollection (XYZ from gp);


    -- HArray2 of 2D objects.

  class HArray2OfCirc2d
    	instantiates HArray2 from PCollection (Circ2d from gp);
  class HArray2OfDir2d
    	instantiates HArray2 from PCollection (Dir2d from gp);
  class HArray2OfLin2d
    	instantiates HArray2 from PCollection (Lin2d from gp);
  class HArray2OfPnt2d
    	instantiates HArray2 from PCollection (Pnt2d from gp);
  class HArray2OfVec2d
    	instantiates HArray2 from PCollection (Vec2d from gp);
  class HArray2OfXY
    	instantiates HArray2 from PCollection (XY from gp);


    -- HArray2 of 3D objects.

  class HArray2OfDir
    	instantiates HArray2 from PCollection (Dir from gp);
  class HArray2OfPnt
    	instantiates HArray2 from PCollection (Pnt from gp);
  class HArray2OfVec
    	instantiates HArray2 from PCollection (Vec from gp);
  class HArray2OfXYZ
    	instantiates HArray2 from PCollection (XYZ from gp);


    -- HSequences of 2D objects.

  class HSequenceOfDir
    	instantiates HSequence  from PCollection (Dir from gp);
  class HSequenceOfPnt
    	instantiates HSequence  from PCollection (Pnt from gp);
  class HSequenceOfVec
    	instantiates HSequence  from PCollection (Vec from gp);
  class HSequenceOfXYZ
    	instantiates HSequence  from PCollection (XYZ from gp);


    -- HSequences of 2D objects.

--  class HSequenceOfDir2d
--    	instantiates HSequence  from PCollection (Dir2d from gp);
--  class HSequenceOfPnt2d
--    	instantiates HSequence  from PCollection (Pnt2d from gp);
--  class HSequenceOfVec2d
--    	instantiates HSequence  from PCollection (Vec2d from gp);
--  class HSequenceOfXY
--    	instantiates HSequence  from PCollection (XY from gp);


end PColgp;
