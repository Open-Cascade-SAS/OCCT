-- File:        Vector.cdl
-- Created:     Fri Dec  1 11:11:31 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class Vector from StepGeom 

inherits GeometricRepresentationItem from StepGeom 

uses

	Direction from StepGeom, 
	Real from Standard, 
	HAsciiString from TCollection
is

	Create returns mutable Vector;
	---Purpose: Returns a Vector


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aOrientation : mutable Direction from StepGeom;
	      aMagnitude : Real from Standard) is virtual;

	-- Specific Methods for Field Data Access --

	SetOrientation(me : mutable; aOrientation : mutable Direction);
	Orientation (me) returns mutable Direction;
	SetMagnitude(me : mutable; aMagnitude : Real);
	Magnitude (me) returns Real;

fields

	orientation : Direction from StepGeom;
	magnitude : Real from Standard;

end Vector;
