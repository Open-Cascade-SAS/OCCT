-- Created on: 1998-07-22
-- Created by: Christian CAILLET
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Vars  from XSDRAW    inherits    Vars  from XSControl

    ---Purpose : Vars for DRAW session (i.e. DBRep and DrawTrSurf)

uses CString, Transient,
     Pnt from gp, Pnt2d from gp,
     Geometry from Geom, Curve from Geom, Curve from Geom2d, Surface from Geom,
     Shape from TopoDS

is

    Create returns mutable Vars from XSDRAW;

    Set (me : mutable; name : CString; val : Transient)  is redefined;

--    Get (me; name : CString) returns Transient  is redefined; unused here


    GetGeom (me; name : in out CString) returns Geometry  is redefined;

    GetCurve2d (me; name : in out CString) returns Curve from Geom2d  is redefined;

    GetCurve   (me; name : in out CString) returns Curve from Geom  is redefined;

    GetSurface (me; name : in out CString) returns Surface from Geom  is redefined;

    SetPoint   (me : mutable; name : CString; val : Pnt   from gp)  is redefined;

    SetPoint2d (me : mutable; name : CString; val : Pnt2d from gp)  is redefined;

    GetPoint   (me; name : in out CString; pnt : out Pnt   from gp) returns Boolean  is redefined;

    GetPoint2d (me; name : in out CString; pnt : out Pnt2d from gp) returns Boolean  is redefined;


    SetShape   (me : mutable; name : CString; val : Shape from TopoDS)  is redefined;

    GetShape   (me; name : in out CString) returns Shape from TopoDS  is redefined;

end Vars;
