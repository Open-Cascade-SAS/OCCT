-- Created on: 1995-07-18
-- Created by: Modelistation
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class CurveTool from Extrema

uses Pnt          from gp,
     Vec          from gp,
     Circ         from gp,
     Elips        from gp,
     Hypr         from gp,
     Parab        from gp,
     Lin          from gp,
     Array1OfReal from TColStd,
     BezierCurve  from Geom,
     BSplineCurve from Geom,
     CurveType    from GeomAbs,
     Shape        from GeomAbs,
     Curve        from Adaptor3d
     
is


    FirstParameter(myclass; C : Curve from Adaptor3d)
    returns Real from Standard;
    	---C++: inline

    LastParameter(myclass; C : Curve from Adaptor3d)
    returns Real from Standard;
    	---C++: inline
    
    Continuity(myclass; C: Curve from Adaptor3d) returns Shape from GeomAbs;
    	---C++: inline

    NbIntervals(myclass; C: in out Curve from Adaptor3d; S : Shape from GeomAbs) returns Integer;
	---Purpose: Returns  the number  of  intervals for  continuity
	--          <S>. May be one if Continuity(me) >= <S>
    	---C++: inline


    Intervals(myclass; C: in out Curve from Adaptor3d; T : in out Array1OfReal from TColStd; 
    	          S : Shape from GeomAbs);
	---Purpose: Stores in <T> the  parameters bounding the intervals
	--          of continuity <S>.
	--          
	--          The array must provide  enough room to  accomodate
	--          for the parameters. i.e. T.Length() > NbIntervals()
    	---C++: inline
    
    IsPeriodic(myclass;C: Curve from Adaptor3d) returns Boolean;
 
    Period(myclass; C: Curve from Adaptor3d) returns Real;
    	---C++: inline


    Resolution(myclass; C: Curve from Adaptor3d; R3d: Real) returns Real;
    	---C++: inline


    GetType(myclass;C: Curve from Adaptor3d) returns CurveType from GeomAbs;
    	---C++: inline


    Value(myclass; C : Curve from Adaptor3d;
                   U : Real    from Standard)
    returns Pnt from gp;
    	---C++: inline
    
    D1 (myclass; C :     Curve from Adaptor3d;
                 U :     Real    from Standard;
                 P : out Pnt from gp;
                 V : out Vec from gp);
    	---C++: inline
    
    D2 (myclass; C      :     Curve from Adaptor3d;
                 U      :     Real    from Standard;
                 P      : out Pnt from gp;
                 V1, V2 : out Vec from gp);
     	---C++: inline

   Line(myclass; C : Curve from Adaptor3d) returns Lin from gp;
     	---C++: inline
   
   Circle(myclass; C : Curve from Adaptor3d) returns Circ from gp;
     	---C++: inline

   Ellipse(myclass; C : Curve from Adaptor3d) returns Elips from gp;
     	---C++: inline

   Hyperbola(myclass; C : Curve from Adaptor3d) returns  Hypr from gp;
     	---C++: inline

   Parabola(myclass; C : Curve from Adaptor3d) returns Parab from gp;
     	---C++: inline

   Degree(myclass; C : Curve from Adaptor3d) returns Integer;
     	---C++: inline
     
   IsRational(myclass; C : Curve from Adaptor3d) returns Boolean;
     	---C++: inline
     
   NbPoles(myclass; C : Curve from Adaptor3d) returns Integer;
     	---C++: inline
     
   NbKnots(myclass; C : Curve from Adaptor3d) returns Integer;
     	---C++: inline
     
   Bezier(myclass; C : Curve from Adaptor3d) returns BezierCurve from Geom;
     	---C++: inline

   BSpline(myclass; C : Curve from Adaptor3d) returns BSplineCurve from Geom;
     	---C++: inline
     

end CurveTool;
