-- Created on: 1995-01-26
-- Created by: CAL
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


-- Modified: TCL G002A, 28-11-00, new section "inquire methods"
-- SAV 04/07/02 : DrawVertex() redefined.


class Marker from Graphic2d inherits Line from Graphic2d

	---Version:

	---Purpose: The primitive Marker

	---Keywords: Primitive, Marker
	---Warning:
	---References:

uses
	Drawer		from Graphic2d,
	GraphicObject	from Graphic2d,
	Length		from Quantity,
	PlaneAngle	from Quantity, 
	FStream         from Aspect,
	IFStream	from Aspect


raises
	MarkerDefinitionError	from Graphic2d

is
	-------------------------
	-- Category: Constructors
	-------------------------

	Create (aGraphicObject: GraphicObject from Graphic2d;
		X, Y: Length from Quantity)
	returns mutable Marker from Graphic2d;
	---Level: Public
	---Purpose: Creates a pixel point marker at position <X>,<Y>
	---Category: Constructors

	Create (aGraphicObject: GraphicObject from Graphic2d;
		anIndex: Integer from Standard;
		X, Y: Length from Quantity;
		aWidth: Length from Quantity;
		anHeight: Length from Quantity;
		anAngle: PlaneAngle from Quantity = 0.0)
	returns mutable Marker from Graphic2d
	---Level: Public
	---Purpose: Creates the predefined marker index <anIndex> 
	--	    at position <X>,<Y> and size <aWidth>,<aHeight>.
	--	    Angle is measured counterclockwise with 0 radian
	--	    at 3 o'clock.
	---Category: Constructors
	---Trigger: Raises MarkerDefinitionError if the
	--	    marker index is <= 0 or undefined in the MarkMap,
	--          or the marker size <aWidth,anHeight> is null.
	raises MarkerDefinitionError from Graphic2d;

	--------------------------
	-- Category: Draw and Pick
	--------------------------

	Draw (me : mutable; aDrawer: Drawer from Graphic2d)
	is static protected;
	---Level: Internal
	---Purpose: Draws the marker <me>.

	Pick (me : mutable; X, Y: ShortReal from Standard;
		aPrecision: ShortReal from Standard;
		aDrawer: Drawer from Graphic2d)
	returns Boolean from Standard
	is static protected;
	---Level: Internal
	---Purpose: Returns Standard_True if the marker <me> is picked,
	--	    Standard_False if not.
	--  Warning: Checks only if the point <X>, <Y> is in the
	--	    boundary rectangle of <me>

	DrawVertex( me : mutable; aDrawer: Drawer from Graphic2d;
                    anIndex: Integer from Standard)
        is redefined protected;

     --------------------------------------
	-- Category: Inquire methods
	--------------------------------------

    Position( me; X, Y: out Length from Quantity );  
	---Level: Public
	---Purpose: returns the coordinates of the position of the marker
	
    Size( me; aW, aH: out Length from Quantity );  
	---Level: Public
	---Purpose: returns the width and height of the marker
	
	Index( me ) returns Integer from Standard;
	---Level: Public
	---Purpose: returns the index of marker in the map of markers
	
    Angle( me ) returns PlaneAngle from Quantity;
	---Level: Public
	---Purpose: returns the angle of the marker

	----------------------------------------------------------------------

	Save( me; aFStream: in out FStream from Aspect ) is virtual;
--	Retrieve( me; aIFStream: in out IFStream from AIS2D ) is virtual;

fields

	myMarkIndex: Integer from Standard;
	myX:		 ShortReal from Standard;
	myY:		 ShortReal from Standard;
	myWidth:	 ShortReal from Standard;
	myHeight:	 ShortReal from Standard;
	myAngle:	 ShortReal from Standard;

end Marker from Graphic2d;
