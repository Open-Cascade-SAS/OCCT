-- File:	RWStepBasic_RWIdentificationRole.cdl
-- Created:	Wed May 10 15:09:08 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class RWIdentificationRole from RWStepBasic

    ---Purpose: Read & Write tool for IdentificationRole

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    IdentificationRole from StepBasic

is
    Create returns RWIdentificationRole from RWStepBasic;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : IdentificationRole from StepBasic);
	---Purpose: Reads IdentificationRole

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: IdentificationRole from StepBasic);
	---Purpose: Writes IdentificationRole

    Share (me; ent : IdentificationRole from StepBasic;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWIdentificationRole;
