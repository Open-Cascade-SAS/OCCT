-- Created on: 1993-01-09
-- Created by: CKY / Contract Toubro-Larsen ( TCD )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class DrawingSize from IGESGraph  inherits IGESEntity

        ---Purpose: defines IGESDrawingSize, Type <406> Form <16>
        --          in package IGESGraph
        --
        --          Specifies the drawing size in drawing units. The
        --          origin of the drawing is defined to be (0,0) in
        --          drawing space

uses  Integer, Real  -- no one specific type


is

        Create returns mutable DrawingSize;

        -- Specific Methods pertaining to the class

        Init (me      : mutable;
              nbProps : Integer;
              aXSize  : Real;
              aYSize  : Real);
        ---Purpose : This method is used to set the fields of the class
        --           DrawingSize
        --      - nbProps : Number of property values (NP = 2)
        --      - aXSize  : Extent of Drawing along positive XD axis
        --      - aYSize  : Extent of Drawing along positive YD axis

        -- Specific Access Methods : According to each type of Entity

        NbPropertyValues (me) returns Integer;
        ---Purpose : returns the number of property values in <me> (NP = 2)

        XSize (me) returns Real;
        ---Purpose : returns the extent of Drawing along positive XD axis

        YSize (me) returns Real;
        ---Purpose : returns the extent of Drawing along positive YD axis

fields

--
-- Class    : IGESGraph_DrawingSize
--
-- Purpose  : Declaration of the variables specific to a Drawing Size.
--
-- Reminder : A Drawing Size is defined by :
--                  - Number of property values
--                  - X Size
--                  - Y Size
--

        theNbPropertyValues : Integer;

        theXSize            : Real;

        theYSize            : Real;

end DrawingSize;
