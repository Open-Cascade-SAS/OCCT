-- Created on: 2000-01-19
-- Created by: data exchange team
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class AlgoContainer from XSAlgo inherits TShared from MMgt

    ---Purpose: 

uses

    Curve             from Geom2d,
    Surface           from Geom,
    Edge              from TopoDS,
    Face              from TopoDS,
    Shape             from TopoDS,
    Caller            from XSAlgo,
    ToolContainer     from XSAlgo,
    WireData          from ShapeExtend,
    Wire              from ShapeAnalysis,
    Wire              from ShapeFix,
    TransientProcess  from Transfer,
    FinderProcess     from Transfer,
    ProgressIndicator from Message
    
is

    Create returns mutable AlgoContainer from XSAlgo;
    	---Purpose: Empty constructor
	
    SetToolContainer (me: mutable; TC: ToolContainer from XSAlgo);
    	---C++    : inline
    	---Purpose: Sets ToolContainer
	
    ToolContainer (me) returns ToolContainer from XSAlgo;
    	---C++    : inline
    	---Purpose: Returns ToolContainer
	

    PrepareForTransfer (me) is virtual;
    	---Purpose: Performs actions necessary for preparing environment
    	--          for transfer. Empty in Open version.
	
    ProcessShape (me; shape:
                  Shape from TopoDS; 
                  Prec, MaxTol: Real;
                  rscfile: CString;
                  seq: CString;
                  info: out Transient;
                  progress: ProgressIndicator from Message = 0)
    returns Shape from TopoDS is virtual;
    	---Purpose: Does shape processing with specified tolerances
    	--          and returns resulting shape and associated information 
      --          in the form of Transient.
      --          This information should be later transmitted to 
      --          MergeTransferInfo in order to be recorded in the
      --          translation map
      --
      ---Default behaviour:
      --          Applies sequence with name identified by parameter named 
      --          <seq> (see Interface_Static), defined in resource file
      --          identified by parameter with name <rscfile>, to shape,
      --          and keeps info of substitutions made during the process.
      --          The Prec and MaxTol define run-time parameters 
      --          Runtime.Tolerance and Runtime.MaxTolerance which can be 
      --          referred from the resource file
      --          ("param : &Runtime.Tolerance")
      --          In the info returns ShapeProcess_ShapeContext with recorded
      --          modifications. If info has already this type on input, uses it.
      --
      --          If resource file is not found, or sequence is not defined 
      --          there, performs default fixes:
      --        - if <seq> is write.iges.sequence or write.step.sequence, does DirectFaces
      --        - if <seq> is read.iges.sequence or read.step.sequence, performs FixShape

    CheckPCurve (me; edge  : Edge from TopoDS;
                 face  : Face from TopoDS;
                 preci : Real;
                 isSeam: Boolean)
    returns Boolean is virtual;
    	---Purpose: Checks quality of pcurve of the edge on the given face, 
      --          and corrects it if necessary.
      ---Remark : In Open CASCADE does nothing.

    MergeTransferInfo (me; TP : TransientProcess from Transfer;
                       info: Transient;
                       startTPitem: Integer = 1) is virtual;
    MergeTransferInfo (me; FP : FinderProcess from Transfer;
                       info: Transient) is virtual;
    	---Purpose: Updates translation map (TP or FP) with information
    	--          resulting from ShapeProcessing
    	--          Parameter startTPitem can be used for optimisation, to
    	--          restrict modifications to entities stored in TP starting
    	--          from item startTPitem

fields

    myTC : ToolContainer from XSAlgo;
    
end AlgoContainer;
