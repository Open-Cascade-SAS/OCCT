-- Created on: 1997-05-06
-- Created by: Jean-Louis Frenkel, Remi Lequette
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package CDM


uses TCollection,TColStd,Resource

is

    enumeration CanCloseStatus is CCS_OK, CCS_NotOpen, CCS_UnstoredReferenced,CCS_ModifiedReferenced,CCS_ReferenceRejection
    end CanCloseStatus from CDM;


    class MetaData;

    deferred class MessageDriver;

    deferred class Document;

    class ReferenceIterator;

    class NullMessageDriver; 

    class COutMessageDriver;


---Category: classes to manager automatic naming of documents.

    private alias NamesDirectory is DataMapOfStringInteger from TColStd;
    ---Purpose: this map will allows to get a directory object from a name.

    imported PresentationDirectory;

    imported DataMapIteratorOfPresentationDirectory;
    ---Purpose: this map will allows to get a directory object from a name.
         
    private pointer DocumentPointer to Document from CDM;
    private class Reference;    

    imported ListOfReferences;

    imported ListIteratorOfListOfReferences;
    deferred class Application;
    
    imported MetaDataLookUpTable;
    
    imported DataMapIteratorOfMetaDataLookUpTable;
         
         
---Category: reusable classes

    imported DocumentHasher;
    imported MapOfDocument;
    imported MapIteratorOfMapOfDocument;
    imported ListOfDocument;
    imported ListIteratorOfListOfDocument;

end CDM;
