-- Created on: 2000-05-24
-- Created by: data exchange team
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Application from XCAFApp inherits Application from TDocStd

    ---Purpose: Implements an Application for the DECAF documents

uses
    SequenceOfExtendedString from TColStd,
    Document from TDocStd

is

    Create returns Application from XCAFApp is protected;


    ---Purpose: methods from CDF_Application
    --          ============================


    Formats(me: mutable; Formats: out SequenceOfExtendedString from TColStd) 
    is redefined;    


    ResourcesName (me: mutable) returns CString from Standard is redefined;

    ---Purpose: methods from TDocStd_Application
    --          ================================

    InitDocument (me; aDoc : Document from TDocStd) is redefined;
    ---Purpose: Set XCAFDoc_DocumentTool attribute
    
    ---API: method for initialisation

    GetApplication (myclass) returns Application from XCAFApp;
    ---Purpose: Initializes (for the first time) and returns the 
    --          static object (XCAFApp_Application)
    --          This is the only valid method to get XCAFApp_Application
    --          object, and it should be called at least once before
    --          any actions with documents in order to init application

end Application;
