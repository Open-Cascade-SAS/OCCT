-- Created on: 1993-01-09
-- Created by: CKY / Contract Toubro-Larsen ( SIVA )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SolidOfLinearExtrusion from IGESSolid  inherits IGESEntity

        ---Purpose: defines SolidOfLinearExtrusion, Type <164> Form Number <0>
        --          in package IGESSolid
        --          Solid of linear extrusion is defined by translatin an
        --          area determined by a planar curve

uses

        Dir             from gp,
        XYZ             from gp

is

        Create returns SolidOfLinearExtrusion;

        -- Specific Methods pertaining to the class

        Init (me         : mutable;
              aCurve     : IGESEntity;
              aLength    : Real;
              aDirection : XYZ);
        ---Purpose : This method is used to set the fields of the class
        --           SolidOfLinearExtrusion
        --       - aCurve     : the planar curve that is to be translated
        --       - aLength    : the length of extrusion
        --       - aDirection : the vector specifying the direction of extrusion
        --                      default (0,0,1)

        Curve (me) returns IGESEntity;
        ---Purpose : returns the planar curve that is to be translated

        ExtrusionLength (me) returns Real;
        ---Purpose : returns the Extrusion Length

        ExtrusionDirection (me) returns Dir;
        ---Purpose : returns the Extrusion direction

        TransformedExtrusionDirection (me) returns Dir;
        ---Purpose : returns ExtrusionDirection after applying TransformationMatrix

fields

--
-- Class    : IGESSolid_SolidOfLinearExtrusion
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class SolidOfLinearExtrusion.
--
-- Reminder : A SolidOfLinearExtrusion instance is defined by :
--            a planar curve(Curve) that is translated by a distance(Length)
--            in the direction specified by a vector(I1,J1,K1).
--

        theCurve     : IGESEntity;
            --  the planar curve

        theLength    : Real;
            -- the length of the extrusion

        theDirection : XYZ;
            -- the vector defining the direction of the extrusion

end SolidOfLinearExtrusion;
