-- Created on: 1993-05-12
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



deferred generic class SurfaceTool from Contap
    (TheSurface as any)
                                   

	---Purpose: Template class for a tool on a surface.
	--          It is possible to implement this class with an 
	--          instantiation of the Surface2Tool from Adaptor3d.


uses SurfaceType from GeomAbs,
     Pln         from gp,
     Sphere      from gp,
     Cylinder    from gp,
     Cone        from gp,
     Pnt         from gp,
     Vec         from gp

 is


    GetType(myclass; S: TheSurface)
    
    	returns SurfaceType from GeomAbs;


    Plane(myclass; S: TheSurface)
    
	---Purpose: Returns the plane from gp when GetType returns
	--          GeomAbs_Plane.
    
    	returns Pln from gp;


    Cylinder(myclass; S: TheSurface)
    
	---Purpose: Returns the cylinder from gp when GetType returns
	--          GeomAbs_Cylinder.
    
    	returns Cylinder from gp;


    Sphere(myclass; S: TheSurface)
    
	---Purpose: Returns the sphere from gp when GetType returns
	--          GeomAbs_Sphere.
    
    	returns Sphere from gp;


    Cone(myclass; S: TheSurface)
    
	---Purpose: Returns the cone from gp when GetType returns
	--          GeomAbs_Cone.
    
    	returns Cone from gp;



    UIntervalFirst(myclass ; S: TheSurface)
	   
	---Purpose: Returns the first U parameter of the surface.

    	returns Real from Standard;
    
    
    VIntervalFirst(myclass ; S: TheSurface)
	   
	---Purpose: Returns the first V parameter of the surface.

    	returns Real from Standard;
    
    
    UIntervalLast(myclass ; S: TheSurface)
	   
	---Purpose: Returns the last U parameter of the surface.

    	returns Real from Standard;
    
    
    VIntervalLast(myclass ; S: TheSurface)
	   
	---Purpose: Returns the last V parameter of the surface.

    	returns Real from Standard;
    
    
    Value (myclass ; S: TheSurface;
           U,V : Real from Standard)
	   
	---Purpose: Returns the point of parameter (U,V) on the surface.

    	 returns Pnt from gp;


    D1(myclass; S: TheSurface; U,V: Real from Standard; 
                P: out Pnt from gp; D1U,D1V: out Vec from gp);
		
	---Purpose: Returns the point of parameter (U,V) on the surface,
	--          and the first derivatives in the directions u and v.

    
    D2(myclass; S: TheSurface; U,V: Real from Standard; P: out Pnt from gp;
                       D1U,D1V,D2U,D2V,D2UV: out Vec from gp);
		       
	---Purpose: Returns the point of parameter (U,V) on the surface,
	--          and the first and the second derivatives in the
	--          directions u and v.

    
    UResolution(myclass; S : TheSurface; Tol3d: Real from Standard)
    
	---Purpose: Returns the numerical resolution in the U direction,
	--          for a given resolution in 3d space.

    	returns Real from Standard;


    VResolution(myclass; S : TheSurface; Tol3d: Real from Standard)
    
	---Purpose: Returns the numerical resolution in the V direction,
	--          for a given resolution in 3d space.

    	returns Real from Standard;


end SurfaceTool;
