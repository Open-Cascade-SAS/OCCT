-- Created on: 1995-03-10
-- Created by: Mister rmi
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Modified by rob (18/10/96) : add methods to store a constant sensitivity



deferred class SensitiveEntity from Select2D inherits SensitiveEntity from SelectBasics

	---Purpose: A framework to define what all sensitive 2D entities have in common.
    	-- This framework can be used to create new 2D sensitive entities.

uses 
    EntityOwner  from SelectBasics, 
    Array1OfPnt2d from TColgp, 
    Box2d from Bnd,
    Projector from Select2D 
    
raises 
    NotImplemented from Standard

is

    Initialize(anOwnerId: EntityOwner from SelectBasics);

    NeedsConversion (me) returns Boolean is virtual;
    	---Purpose: returns Standard_False unless if redefined...
    	---Level: Public 
    	---C++: inline

    Convert(me:mutable;aProjector: Projector from Select2D) is virtual;
    	---Purpose: Processes the projection of the sensitive primitives in
    	-- the active view.   This must be performed before the selection action.
    	-- This function must be implemented in daughter classes.
    
    MaxBoxes(me) returns Integer is virtual;
    	---Purpose: Returns the maximum number of boxes.


    SetOwnTolerance(me:mutable; aValue : Real from Standard) ;
    	---Purpose: Sets and stores a tolerance value in the argument
    	-- aTol of the function Matches inherited from SelectBasics_SensitiveEntity.

    UnsetOwnTolerance(me:mutable);
    	---Purpose: Removes the in the argument aTol of the function
    	-- Matches inherited from SelectBasics_SensitiveEntity.
    
    HasOwnTolerance(me) returns Boolean from Standard;
    	---Purpose: Returns true if the entity has a setting for the
    	-- argument aTol   of the function Matches inherited
    	-- from SelectBasics_SensitiveEntity.


    OwnTolerance(me) returns Real from Standard;
    	---Purpose: Returns the tolerance value in the argument aTol of
    	-- the function Matches inherited from SelectBasics_SensitiveEntity.
    
    Is3D(me) returns Boolean from Standard is redefined static;
    	--- Purpose: Returns true if this object can provide 3D information.

        Matches (me  :mutable; 
             Polyline:Array1OfPnt2d from TColgp;
	     aBox:Box2d from Bnd;
             aTol: Real from Standard)
    returns Boolean from Standard is redefined virtual;
    	---Purpose: Free contur selection for 2d is not defined


fields

    myOwnTolerance : Real from Standard is protected;

end SensitiveEntity;
