-- File:	Dynamic_RealParameter.cdl
-- Created:	Wed Feb  3 15:49:43 1993
-- Author:	Gilles DEBARBOUILLE
--		<gde@bravox>
---Copyright:	 Matra Datavision 1993



class RealParameter from Dynamic

inherits

    Parameter from Dynamic
	---Purpose: This  inherited class from Parameter describes all
	--          the parameters, which  are characterized by a real
	--          value.

uses

    OStream from Standard,
    CString from Standard,
    Real    from Standard


is

    Create(aparameter : CString from Standard )
    
    ---Level: Public 
    
    ---Purpose: Creates a RealParameter with <aparameter> as name.
    
    returns mutable RealParameter from Dynamic;

    Create(aparameter : CString from Standard ; avalue : Real from Standard) 
    
    ---Level: Public 
    
    ---Purpose: With  the name  of the Parameter  <aparameter> and the
    --          real <avalue>, creates an instance of RealParameter.
    
    returns mutable RealParameter from Dynamic;
    
    Value(me) returns Real from Standard
    
    ---Level: Public 
    
    ---Purpose: Returns the value of the parameter which is a real.
    
    is static;

    Value (me : mutable ; avalue : Real from Standard)
    
    ---Level: Public 
    
    --- Purpose: Sets the real <avalue> in <me>.

    is static;
    
    Dump(me ; astream : in out OStream from Standard)
    
    ---Level: Internal 
    
    ---Purpose: Useful for debugging.

    is redefined;
    
fields

    thevalue : Real from Standard;

end RealParameter;
