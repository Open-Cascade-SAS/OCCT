-- Created on: 1993-09-30
-- Created by: Denis PASCAL
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class SC from GraphTools inherits TShared from MMgt

    ---Purpose: This  class is used  to  identify a  Strong Component.
    --          The user has not to used its methods.

uses SCList            from GraphTools,
     SequenceOfInteger from TColStd

raises OutOfRange   from Standard,
       NoSuchObject from Standard
    
is

    Create returns mutable SC;
	
    Reset (me : mutable);
    ---Level: Public

    AddVertex (me : mutable; V : Integer from Standard); 
    ---Level: Public

    NbVertices (me) returns Integer from Standard;
    ---Level: Public

    GetVertex (me; index: Integer from Standard) 
    ---Level: Public
    returns Integer from Standard;
	
    AddFrontSC (me : mutable; SC : SC from GraphTools);
    ---Level: Public
 
    GetFrontSC (me) returns SCList from GraphTools;
    ---Level: Public
    ---C++: return const & 	
	
    AddBackSC (me : mutable; SC : SC from GraphTools);
    ---Level: Public

    GetBackSC (me) returns SCList from GraphTools;
    ---Level: Public
    ---C++: return const & 	

fields
	
    myBackSC   : SCList            from GraphTools;
    myVertices : SequenceOfInteger from TColStd;
    myFrontSC  : SCList            from GraphTools;

end SC;


