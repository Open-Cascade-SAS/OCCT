-- File:	StepFEA_SymmetricTensor23d.cdl
-- Created:	Tue Dec 10 18:13:00 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V2.0
-- Copyright:	Open CASCADE 2002

class SymmetricTensor23d from StepFEA
inherits SelectType from StepData

    ---Purpose: Representation of STEP SELECT type SymmetricTensor23d

uses
    SelectMember from StepData,
    HArray1OfReal from TColStd,
    HArray1OfReal from TColStd

is
    Create returns SymmetricTensor23d from StepFEA;
	---Purpose: Empty constructor

    CaseNum (me; ent: Transient) returns Integer;
	---Purpose: Recognizes a kind of SymmetricTensor23d select type
	--          return 0 

    CaseMem (me; ent: SelectMember from StepData) returns Integer is redefined;
	---Purpose: Recognizes a items of select member SymmetricTensor23dMember
	--          1 -> IsotropicSymmetricTensor23d
	--          2 -> OrthotropicSymmetricTensor23d
	--          3 -> AnisotropicSymmetricTensor23d
	--          0 else


     NewMember(me) returns SelectMember from StepData is redefined;
	---Purpose: Returns a new select member the type SymmetricTensor23dMember

    SetIsotropicSymmetricTensor23d(me: in out; aVal :Real);
	---Purpose: Set Value for IsotropicSymmetricTensor23d

    IsotropicSymmetricTensor23d (me) returns Real;
	---Purpose: Returns Value as IsotropicSymmetricTensor23d (or Null if another type)

    SetOrthotropicSymmetricTensor23d(me: in out; aVal :HArray1OfReal from TColStd);
	---Purpose: Set Value for OrthotropicSymmetricTensor23d

    OrthotropicSymmetricTensor23d (me) returns HArray1OfReal from TColStd;
	---Purpose: Returns Value as OrthotropicSymmetricTensor23d (or Null if another type)

    SetAnisotropicSymmetricTensor23d(me: in out; aVal :HArray1OfReal from TColStd);
	---Purpose: Set Value for AnisotropicSymmetricTensor23d

    AnisotropicSymmetricTensor23d (me) returns HArray1OfReal from TColStd;
	---Purpose: Returns Value as AnisotropicSymmetricTensor23d (or Null if another type)

end SymmetricTensor23d;
