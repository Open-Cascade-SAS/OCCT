-- Created on: 1998-06-11
-- Created by: data exchange team
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Vertex from ShapeBuild 

    ---Purpose: Provides low-level functions used for constructing vertices

uses
    Pnt from gp,
    Vertex from TopoDS

is

    CombineVertex ( me; V1, V2: Vertex from TopoDS; tolFactor: Real = 1.0001 ) 
    returns Vertex from TopoDS;
    	---Purpose: Combines new vertex from two others. This new one is the 
    	--          smallest vertex which comprises both of the source vertices. 
    	--          The function takes into account the positions and tolerances 
        --          of the source vertices.
    	--          The tolerance of the new vertex will be equal to the minimal
        --          tolerance that is required to comprise source vertices 
    	--          multiplied by tolFactor (in order to avoid errors because
	--          of discreteness of calculations).

    CombineVertex ( me; pnt1, pnt2: Pnt from gp; tol1, tol2: Real;
    	    	    tolFactor: Real = 1.0001 ) 
    returns Vertex from TopoDS;
    	---Purpose: The same function as above, except that it accepts two points
	--          and two tolerances instead of vertices

end Vertex;
