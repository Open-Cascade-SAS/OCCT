-- Created on: 1995-03-24
-- Created by: Robert COUBLANC
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class SensitiveFace from Select3D 
inherits SensitivePoly from Select3D

    ---Purpose: Sensitive Entity to make a face selectable.
    -- In some cases this class can raise Standard_ConstructionError and 
    -- Standard_OutOfRange exceptions. For more details see Select3D_SensitivePoly.

uses
    EntityOwner       from SelectBasics,
    Projector         from Select3D,
    Lin               from gp,
    ListOfBox2d       from SelectBasics,
    PickArgs          from SelectBasics,
    Array1OfPnt       from TColgp,
    HArray1OfPnt      from TColgp,
    Array1OfPnt2d     from TColgp,
    Box2d             from Bnd,
    TypeOfSensitivity from Select3D,
    Location          from TopLoc, 
    SensitiveEntity   from Select3D

raises
    ConstructionError from Standard,
    OutOfRange from Standard

is

    Create (OwnerId      : EntityOwner from SelectBasics;
            ThePoints    : Array1OfPnt from TColgp;
            Sensitivity  : TypeOfSensitivity = Select3D_TOS_INTERIOR)
     returns mutable SensitiveFace;
        ---Level: Public 
        ---Purpose: Constructs a sensitive face object defined by the
        -- owner OwnerId, the array of points ThePoints, and
        -- the sensitivity type Sensitivity.
        -- The array of points is the outer polygon of the geometric face.

    Create (OwnerId      : EntityOwner from SelectBasics;
            ThePoints    : HArray1OfPnt from TColgp;
            Sensitivity  : TypeOfSensitivity = Select3D_TOS_INTERIOR)
     returns mutable SensitiveFace;
        ---Level: Public 
        ---Purpose: Constructs a sensitive face object defined by the
        -- owner OwnerId, the array of points ThePoints, and
        -- the sensitivity type Sensitivity.
        -- The array of points is the outer polygon of the geometric face.
   
    Matches (me : mutable;
             thePickArgs : PickArgs from SelectBasics;
             theMatchDMin, theMatchDepth : out Real from Standard)
    returns Boolean is redefined virtual;
    ---Level: Public
    ---Purpose: Checks whether the sensitive entity matches the picking
    -- detection area (close to the picking line).
    -- For details please refer to base class declaration.

    Matches (me  :mutable; 
             XMin,YMin,XMax,YMax : Real from Standard;
             aTol: Real from Standard) 
    returns Boolean
    is redefined virtual;
    ---Level: Public 
     
    Matches (me  :mutable; 
             Polyline:Array1OfPnt2d from TColgp;
             aBox:Box2d from Bnd;
             aTol: Real from Standard) 
    returns Boolean
    is redefined virtual;
    ---Level: Public 
    

    ComputeDepth (me;
                  thePickLine : Lin from gp;
                  theDepthMin, theDepthMax : Real from Standard)
    returns Real from Standard
    is virtual;
    ---Level: Public
    ---Purpose: Computes the depth values for all 3D points defining this face and returns
    -- the minimal value among them.
    -- If the "minimal depth" approach is not suitable and gives wrong detection results
    -- in some particular case, a custom sensitive face class can redefine this method.

    ComputeDepth(me;EyeLine: Lin from gp)
    is private;
    ---Level: Public
    ---Purpose: Warning: Obsolete.
    -- Use newer version of the method with min, max limits passed as arguments.

    Dump(me; S: in out OStream;FullDump : Boolean from Standard = Standard_True) is redefined virtual; 

    GetConnected(me: mutable; theLocation : Location from TopLoc) 
    returns SensitiveEntity from Select3D 
    is redefined virtual; 
        ---Level: Public 
        ---Purpose: Returns the copy of this


fields

    mytype          : TypeOfSensitivity;
end SensitiveFace;
