-- Created on: 1993-07-23
-- Created by: Jean Louis FRENKEL
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class IndexPixel from Aspect inherits Pixel from Aspect

is
	Create
	returns IndexPixel from Aspect;

	Create (anIndex: Integer from Standard)
	returns IndexPixel from Aspect;

	Value(me)
	returns Integer from Standard
	is static ;

	SetValue(me: in out; anIndex: Integer from Standard) is static ;

	HashCode (me; Upper : Integer )
	returns Integer
	is redefined static ;
	---Level: Public
	---Purpose: Returns a hashed value denoting <me>. This value is in
	--         the range 1..<Upper>.
	---C++:  function call

	Print( me ; s : in out OStream )
	is redefined static ;
	---Level: Public
	---Purpose : Prints the contents of <me> on the stream <s>

    	IsEqual(me; Other : IndexPixel from Aspect) returns Boolean;
	    ---C++: alias operator==

    	IsNotEqual(me; Other : IndexPixel from Aspect) returns Boolean;
           ---C++: alias operator!=

fields
	myIndex: Integer from Standard;

end IndexPixel from Aspect;
