-- Created on: 1995-04-13
-- Created by: Robert COUBLANC
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class SensitiveBox   from Select3D 
inherits SensitiveEntity from Select3D

	---Purpose: A framework to define selection by a sensitive box.         

uses
    Pnt              from gp,
    Pnt2d            from gp,
    Box              from Bnd,
    Box2d            from Bnd,
    Projector        from Select3D,
    Lin              from gp,
    EntityOwner      from SelectBasics,
    ListOfBox2d      from SelectBasics,
    PickArgs         from SelectBasics,
    Array1OfPnt2d    from TColgp,
    Location         from TopLoc

is


    Create (OwnerId      : EntityOwner from SelectBasics;
    	    BoundingBox  : Box from Bnd)
    returns mutable SensitiveBox;
	---Purpose: Constructs a sensitive box object defined by the
    	-- owner OwnerId, and the bounding box BoundingBox.
    Create (OwnerId         : EntityOwner from SelectBasics;
    	    XMin,YMin,ZMin,
    	    XMax,YMax,ZMax  : Real)
    returns mutable SensitiveBox;
	---	Purpose: Constructs a sensitive box object defined by the
    	-- owner OwnerId, and the coordinates Xmin, YMin, ZMin, XMax, YMax, ZMax.
    	-- Xmin, YMin and ZMin define the minimum point in
    	-- the front lower left hand corner of the box,
    	-- and   XMax, YMax   and ZMax define the maximum
    	-- point in the back upper right hand corner of the box.     
	    
    Project (me:mutable;aProjector : Projector from Select3D) 
    is redefined static;
    	---Level: Public 
    	---Purpose: projection of the sensitive primitive in order to
    	--          get 2D boxes for the Sort Algorithm
    
    Areas   (me:mutable ; boxes : in out ListOfBox2d from SelectBasics) 
    is redefined static;
    	---Level: Public 
    	---Purpose: gives the 2D boxes which represent the Box in the 
    	--          selection process...

    GetConnected(me:mutable;aLocation: Location from TopLoc)
    returns SensitiveEntity from Select3D is redefined static;

    Matches (me : mutable;
             thePickArgs : PickArgs from SelectBasics;
             theMatchDMin, theMatchDepth : out Real from Standard)
    returns Boolean is redefined static;
    ---Level: Public
    ---Purpose: Checks whether the sensitive entity matches the picking
    -- detection area (close to the picking line).
    -- For details please refer to base class declaration.

    Matches (me  :mutable; 
             XMin,YMin,XMax,YMax : Real from Standard;
             aTol: Real from Standard)
    returns Boolean is redefined static;
     
    Matches (me  :mutable; 
             Polyline:Array1OfPnt2d from TColgp;
	     aBox:Box2d from Bnd;
             aTol: Real from Standard) 
    returns Boolean
    is redefined virtual;
    	---Level: Public 
    
   
    ComputeDepth(me;EyeLine: Lin from gp) 
    returns Real from Standard;

    Dump(me; S: in out OStream;FullDump : Boolean from Standard = Standard_True) is redefined virtual;

    Box(me) returns Box from Bnd;
    ---Purpose: Returns the sensitive 3D box used at the time of construction.
    ---C++: inline
    ---C++: return const &


    ProjectBox(me:mutable;aPrj: Projector from Select3D;aBox:Box from Bnd)
    is static private;

fields

    mybox3d   : Box   from Bnd;
    mybox2d   : Box2d from Bnd;

end SensitiveBox;










