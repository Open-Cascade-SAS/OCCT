-- File:	RWStepFEA_RWDummyNode.cdl
-- Created:	Thu Dec 12 17:51:04 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWDummyNode from RWStepFEA

    ---Purpose: Read & Write tool for DummyNode

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    DummyNode from StepFEA

is
    Create returns RWDummyNode from RWStepFEA;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : DummyNode from StepFEA);
	---Purpose: Reads DummyNode

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: DummyNode from StepFEA);
	---Purpose: Writes DummyNode

    Share (me; ent : DummyNode from StepFEA;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWDummyNode;
