-- Created on: 1993-06-17
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package TopOpeBRepTool 

	---Purpose: This package provides services used by the TopOpeBRep
	--          package performing topological operations on the BRep
	--          data structure.
	--          

uses

    Standard,
    TColStd,
    TCollection,
    TColgp,
    TopAbs,
    TopoDS,
    TopTools,
    TopExp,
    GeomAbs,
    Geom,
    GeomAdaptor,
    Geom2d,
    Geom2dAdaptor,
    gp,
    Bnd,
    BRepClass,
    TopClass,
    BRepClass3d,
    BRep,
    BRepAdaptor,
    Geom2dInt,
    IntSurf

is

    enumeration OutCurveType is 
    BSPLINE1,APPROX,INTERPOL
    end OutCurveType; 
     
    class GeomTool;
    class AncestorsTool;

    pointer PSoClassif to SolidClassifier from BRepClass3d;

    class C2DF;
    imported ListOfC2DF;
    imported ListIteratorOfListOfC2DF;    
    imported DataMapOfOrientedShapeC2DF;
    imported DataMapIteratorOfDataMapOfOrientedShapeC2DF;
    imported DataMapOfShapeListOfC2DF;
    imported DataMapIteratorOfDataMapOfShapeListOfC2DF;
    
    imported IndexedDataMapOfSolidClassifier;
	 
    imported Plos;
    class SolidClassifier;
    
    class CurveTool;
    imported IndexedDataMapOfShapeBox2d;
    imported IndexedDataMapOfShapeBox;

    class HBoxTool;
    class BoxSort;

    class ShapeExplorer;
    class ShapeTool;
    class ShapeClassifier;
    pointer PShapeClassifier to ShapeClassifier from TopOpeBRepTool;

    class connexity;
    imported IndexedDataMapOfShapeconnexity; 

    class face;
    imported DataMapOfShapeface;
    imported DataMapIteratorOfDataMapOfShapeface; 
    class CLASSI;
    
    class TOOL;	    
    class CORRISO;	
    class REGUW;	    
    class REGUS;	    

    class makeTransition;
    class mkTondgE;
    
    class PurgeInternalEdges;

    class FuseEdges;
    ---Purpose:  Fuse  edges (in a   wire) of a  shape   where we have
    --          useless vertex.

   
    PurgeClosingEdges(F, FF   : in Face from TopoDS; 
    	    	      MWisOld : in DataMapOfShapeInteger from TopTools;
		      MshNOK  : in out IndexedMapOfOrientedShape from TopTools)
    returns Boolean from Standard;
    ---Purpose: In case face <FF> is built on UV-non-connexed  wires
    --          (with the two closing edges  FORWARD and REVERSED, in
    --          spite of one only), we find out the faulty edge, add 
    --          the faulty shapes (edge,wire,face) to <MshNOK>.
    --          <FF> is a face descendant of <F>.
    --          <MWisOld>(wire) = 1 if wire is wire of <F>
    --                            0    wire results from <F>'s wire splitted.
    --          returns false if purge fails                  
		      
    PurgeClosingEdges(F       : in Face from TopoDS; 
    	    	      LOF     : in ListOfShape from TopTools;
    	    	      MWisOld : in DataMapOfShapeInteger from TopTools;
		      MshNOK  : out IndexedMapOfOrientedShape from TopTools)
    returns Boolean from Standard;	
    --          <LOF> is the list of <F>'s descendant faces.
    --          returns false if purge fails    

    CorrectONUVISO(F       : in Face from TopoDS; 
    	    	   Fsp     : in out Face from TopoDS)
    returns Boolean from Standard;	
    --            <Fsp> is one of  <F>'s split, corrects <Fsp> to have
    --           it connexed in UV space.

    MakeFaces(F      : in Face from TopoDS; 
              LOF    : in ListOfShape from TopTools;
	      MshNOK : in IndexedMapOfOrientedShape from TopTools;
    	      LOFF   : out ListOfShape from TopTools)	
    returns Boolean from Standard;
    ---Purpose: Builds up the correct list of faces <LOFF> from <LOF>, using
    --          faulty shapes from map <MshNOK>.	
    --          <LOF> is the list of <F>'s descendant faces.
    --          returns false if building fails    
    		   
    Regularize(aFace : in Face from TopoDS;
    	       aListOfFaces : out ListOfShape from TopTools;
	       ESplits : in out DataMapOfShapeListOfShape from TopTools)
    returns Boolean from Standard;
    ---Purpose: Returns <False>  if  the  face is  valid (the UV
    --          representation  of  the  face is   a set   of  pcurves
    --          connexed by points with   connexity 2).  
    --          Else,  splits <aFace> in order to return a list of valid 
    --          faces.
    
    RegularizeWires(aFace : in Face from TopoDS;
    	            OldWiresNewWires : out DataMapOfShapeListOfShape from TopTools;		 
	       	    ESplits : in out DataMapOfShapeListOfShape from TopTools)
    returns Boolean from Standard;
    ---Purpose: Returns <False>  if  the  face is  valid (the UV
    --          representation  of  the  face is   a set   of  pcurves
    --          connexed by points with   connexity 2).  
    --          Else,  splits wires of the face, these are boundaries of the
    --          new faces to build up; <OldWiresNewWires> describes (wire,
    --          splits of wire); <ESplits> describes (edge, edge's splits) 
        
    RegularizeFace(aFace : in Face from TopoDS;
    	           OldWiresnewWires : in DataMapOfShapeListOfShape from TopTools;	 
	           aListOfFaces : out ListOfShape from TopTools)
    returns Boolean from Standard;
    ---Purpose:  Classify wire's splits of map <OldWiresnewWires> in order to 
    --           compute <aListOfFaces>, the splits of <aFace>.

    RegularizeShells(aSolid : in Solid from TopoDS;
    	    	     OldSheNewShe : out DataMapOfShapeListOfShape from TopTools;	
		     FSplits : in out DataMapOfShapeListOfShape from TopTools)
    returns Boolean from Standard; 
    ---Purpose: Returns <False> if the shell is valid (the solid is a set
    --          of faces connexed by edges with connexity 2).
    --          Else, splits faces of the shell; <OldFacesnewFaces> describes
    --          (face, splits of face).
    
    -- NYI RegularizeSolid(...)

    Print(OCT  : OutCurveType from TopOpeBRepTool; S  : in out OStream) 
    returns OStream;
    ---C++: return &
    ---Purpose: Prints <OCT> as string on stream <S>; returns <S>.

	
end TopOpeBRepTool;
