-- Created on: 1997-04-23
-- Created by: Alexander BRIVIN
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Curve from VrmlConverter 

    	---Purpose: Curve - computes the presentation of objects to be
    	--          seen  as curves  (the  computation  will  be  made
    	--          with a constant  number  of  points),  converts this one
    	--          into  VRML  objects  and  writes (adds) them  into
    	--          anOStream.   All  requested   properties  of   the
    	--          representation are specify  in aDrawer  of  Drawer
    	--          class (VrmlConverter).    
    	--          This kind of the presentation is converted into   
    	--          IndexedLineSet ( VRML ). 

    
uses
 
    Curve    from   Adaptor3d,
    Length   from   Quantity,
    Drawer   from   VrmlConverter

is

    Add(myclass; aCurve     : Curve          from Adaptor3d;
                 aDrawer    : Drawer         from VrmlConverter;
    	    	 anOStream  : in out OStream from Standard);

    ---Purpose: adds to the OStream the drawing of the curve aCurve.
    --          The aspect is defined by LineAspect in aDrawer.
    --          


    Add(myclass; aCurve     : Curve          from Adaptor3d;
                 U1,U2      : Real           from Standard;
                 aDrawer    : Drawer         from VrmlConverter;
    	    	 anOStream  : in out OStream from Standard);
		    
    ---Purpose: adds to the OStream the drawing of the curve aCurve.
    --          The aspect is defined by LineAspect in aDrawer.
    --          The drawing will be limited between the points of parameter
    --          U1 and U2.

    Add(myclass; aCurve       : Curve          from Adaptor3d;
    	    	 U1, U2       : Real           from Standard;
    	    	 anOStream    : in out OStream from Standard;
    	    	 aNbPoints    : Integer        from Standard);

    ---Purpose: adds to the OStream the drawing of the curve aCurve.
    --          The aspect is the current aspect.
    --          The drawing will be limited between the points of parameter
    --          U1 and U2. aNbPoints defines  number of points on  one interval. 

end Curve;
