-- Created on: 1994-09-02
-- Created by: Yves FRICAUD
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

generic class NumericCurInf from LProp (Curve as any;
    	    	    	    	        Vec   as any; -- as Vec or Vec2d
		     	                Pnt   as any; -- as Pnt or Pnt2d
		   	                Dir   as any; -- as Dir or Dir2d Vec  
    	    	    	    	    	Tool  as any) -- as Tool(Curve, Pnt, Vec) 
					
	---Purpose: Computes the locals extremas of curvature and the 
    	--          inflections of a bounded curve in 2d. 

uses
    CurAndInf from LProp
    
private class FCurExt instantiates FuncCurExt from LProp (Curve,Vec,Pnt,Dir,Tool); 
private class FCurNul instantiates FuncCurNul from LProp (Curve,Vec,Pnt,Dir,Tool);

is
    Create;
    
    PerformCurExt (me : in out; C : Curve; Result : in out CurAndInf) 
    	---Purpose: Computes the locals extremas of curvature.
    is static;
    
    PerformInf    (me : in out; C : Curve; Result : in out CurAndInf)
       	---Purpose: Computes the inflections.
    is static;
    
    PerformCurExt (me     : in out; 
    	           C      : Curve ; 
                   UMin   : Real;
    	    	   UMax   : Real;
    	    	   Result : in out CurAndInf) 
    	---Purpose: Computes the locals extremas of curvature.
    	--          in the interval of parmeters [UMin,UMax].
    is static;
    
    PerformInf    (me     : in out;
        	   C      : Curve ; 
                   UMin   : Real;
    	    	   UMax   : Real;
    	    	   Result : in out CurAndInf)
       	---Purpose: Computes the inflections in the interval of 
       	--          parmeters [UMin,UMax].
    is static;
    
    IsDone (me) returns Boolean
	---Purpose: True if the solutions are found.
    is static;
    
fields
    isDone : Boolean from Standard;

end NumericCurInf;
