-- File:        PresentationStyleByContext.cdl
-- Created:     Mon Dec  4 12:02:29 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWPresentationStyleByContext from RWStepVisual

	---Purpose : Read & Write Module for PresentationStyleByContext

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     PresentationStyleByContext from StepVisual,
     EntityIterator from Interface

is

	Create returns RWPresentationStyleByContext;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable PresentationStyleByContext from StepVisual);

	WriteStep (me; SW : in out StepWriter; ent : PresentationStyleByContext from StepVisual);

	Share(me; ent : PresentationStyleByContext from StepVisual; iter : in out EntityIterator);

end RWPresentationStyleByContext;
