-- Created on: 1995-01-25
-- Created by: Jean-Louis Frenkel
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Modified by Rob : 20-feb-1997
-- Modified by Rob : 16-dec-1997 : kind of presentation

deferred class Presentation from PrsMgr
inherits TShared  from MMgt

uses 

    PresentationManager from PrsMgr,
    KindOfPrs from PrsMgr

is

    Initialize(aPresentationManager: PresentationManager from PrsMgr)
    is protected;

    KindOfPresentation(me) returns KindOfPrs from PrsMgr is deferred;    
    ---Purpose: 2D or 3D
    
    Display(me: mutable) is deferred private;
    
    Erase(me: mutable) is deferred private;

    SetVisible (me: mutable; theValue: Boolean from Standard) is deferred private;

    Highlight(me: mutable) is deferred private;
    
    Unhighlight (me) is deferred private;
    
    IsHighlighted(me) returns Boolean from Standard
    is deferred private;

    IsDisplayed(me) returns Boolean from Standard
    is deferred private;

    Destroy ( me : mutable )
    is virtual; 
    ---Level: Public    
    ---Purpose: Destructor
    ---C++:     alias ~

    DisplayPriority(me) returns Integer from Standard
    is deferred private;
    
    SetDisplayPriority(me:mutable;aNewPrior:Integer from Standard)
    is deferred private;

    SetZLayer ( me : mutable;
                theLayerId : Integer from Standard )
      is deferred private;
    ---Purpose: Set Z layer ID for the presentation

    GetZLayer ( me )
      returns Integer from Standard is deferred private;
    ---Purpose: Get Z layer ID for the presentation

    Clear(me: mutable) 
    is deferred private;
    
---Category: Inquire Methods
--            
    PresentationManager(me) returns mutable PresentationManager
    ---Purpose: returns the PresentationManager in which the
    --          presentation has been created.
    is static;
    ---C++: inline
    ---C++: return const&


---Category: Internal Methods

    SetUpdateStatus(me:mutable; aStat : Boolean from Standard);
    ---C++: inline
    
    MustBeUpdated(me) returns Boolean from Standard;
    ---C++: inline


fields

    myPresentationManager: PresentationManager from PrsMgr is protected;
    myMustBeUpdated      : Boolean from Standard is protected;

friends
    class PresentationManager from PrsMgr
        
end Presentation from PrsMgr;
