-- Created on: 2000-02-14
-- Created by: Denis PASCAL
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

private class NamingTool from TNaming 

	---Purpose: 


uses Label   from TDF,
     LabelMap from TDF,
     NamedShape from TNaming,
     MapOfShape from TopTools,
     Shape      from TopoDS


is


    CurrentShape  (myclass;
    	           Valid    :        LabelMap   from TDF;
                   Forbiden :        LabelMap   from TDF;
		   NS       :        NamedShape from TNaming;
		   MS       : in out MapOfShape from TopTools);
		   
    CurrentShapeFromShape  (myclass;
                            Valid    :        LabelMap   from TDF;
                    	    Forbiden :        LabelMap   from TDF;
		    	    Acces    :        Label      from TDF;
		    	    S        :        Shape      from TopoDS;
		    	    MS       : in out MapOfShape from TopTools);
		   
    BuildDescendants (myclass;
                      NS       : NamedShape from TNaming;
    	    	      Labels   : in out LabelMap   from TDF);



end NamingTool from TNaming;



