-- Created on: 1999-10-11
-- Created by: data exchange team
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SiUnitAndAreaUnit from StepBasic inherits SiUnit from StepBasic

	---Purpose: 

uses

    AreaUnit from StepBasic,
    DimensionalExponents

is

    Create returns mutable SiUnitAndAreaUnit from StepBasic;
    	---Purpose: Returns a SiUnitAndAreaUnit
    
    SetAreaUnit(me: mutable; anAreaUnit: mutable AreaUnit from StepBasic);
    
    AreaUnit(me) returns mutable AreaUnit from StepBasic;
    
    SetDimensions(me : mutable; aDimensions : mutable DimensionalExponents) is redefined;
    
    Dimensions(me) returns mutable DimensionalExponents is redefined;
    
fields

    areaUnit: AreaUnit from StepBasic;

end SiUnitAndAreaUnit;
