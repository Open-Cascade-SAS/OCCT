-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DateTimeSelect from StepBasic inherits SelectType from StepData

	-- <DateTimeSelect> is an EXPRESS Select Type construct translation.
	-- it gathers : Date, LocalTime, DateAndTime

uses

	Date,
	LocalTime,
	DateAndTime
is

	Create returns DateTimeSelect;
	---Purpose : Returns a DateTimeSelect SelectType

	CaseNum (me; ent : Transient) returns Integer;
	---Purpose: Recognizes a DateTimeSelect Kind Entity that is :
	--        1 -> Date
	--        2 -> LocalTime
	--        3 -> DateAndTime
	--        0 else

	Date (me) returns any Date;
	---Purpose : returns Value as a Date (Null if another type)

	LocalTime (me) returns any LocalTime;
	---Purpose : returns Value as a LocalTime (Null if another type)

	DateAndTime (me) returns any DateAndTime;
	---Purpose : returns Value as a DateAndTime (Null if another type)


end DateTimeSelect;

