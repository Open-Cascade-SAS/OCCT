-- Created on: 2002-12-12
-- Created by: data exchange team
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class Surface3dElementDescriptor from StepElement
inherits ElementDescriptor from StepElement

    ---Purpose: Representation of STEP entity Surface3dElementDescriptor

uses
    ElementOrder from StepElement,
    HAsciiString from TCollection,
    HArray1OfHSequenceOfSurfaceElementPurposeMember from StepElement,
    Element2dShape from StepElement

is
    Create returns Surface3dElementDescriptor from StepElement;
	---Purpose: Empty constructor

    Init (me: mutable; aElementDescriptor_TopologyOrder: ElementOrder from StepElement;
                       aElementDescriptor_Description: HAsciiString from TCollection;
                       aPurpose: HArray1OfHSequenceOfSurfaceElementPurposeMember from StepElement;
                       aShape: Element2dShape from StepElement);
	---Purpose: Initialize all fields (own and inherited)

    Purpose (me) returns HArray1OfHSequenceOfSurfaceElementPurposeMember from StepElement;
	---Purpose: Returns field Purpose
    SetPurpose (me: mutable; Purpose: HArray1OfHSequenceOfSurfaceElementPurposeMember from StepElement);
	---Purpose: Set field Purpose

    Shape (me) returns Element2dShape from StepElement;
	---Purpose: Returns field Shape
    SetShape (me: mutable; Shape: Element2dShape from StepElement);
	---Purpose: Set field Shape

fields
    thePurpose: HArray1OfHSequenceOfSurfaceElementPurposeMember from StepElement;
    theShape: Element2dShape from StepElement;

end Surface3dElementDescriptor;
