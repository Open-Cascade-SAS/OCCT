-- Created on: 2004-03-05
-- Created by: Mikhail KUZMITCHEV
-- Copyright (c) 2004-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


package QANCollection

uses
    Draw,
    TCollection, 
    TColStd,
    gp

is
    class  ListOfPnt   instantiates  List  from  TCollection    (Pnt  from  gp);
    class  QueueOfPnt  instantiates  Queue from  TCollection    (Pnt  from  gp);
    class  StackOfPnt  instantiates  Stack from  TCollection    (Pnt  from  gp);
    class  SListOfPnt  instantiates  SList from  TCollection    (Pnt  from  gp);
    class  DataMapOfRealPnt instantiates DataMap from TCollection  
                                        (Real from Standard, 
                                         Pnt from gp, 
                                         MapRealHasher from TColStd);
    class  IndexedDataMapOfRealPnt instantiates IndexedDataMap from TCollection
                                        (Real from Standard, 
                                         Pnt from gp, 
                                         MapRealHasher from TColStd);
    class  DoubleMapOfRealInteger instantiates DoubleMap from TCollection  
                                        (Real from Standard, 
                                         Integer from Standard, 
                                         MapRealHasher from TColStd, 
                                         MapIntegerHasher from TColStd);


---    HashCode (thePnt   : Pnt from gp;
---              theUpper : Integer from Standard)
---    returns Integer from Standard;
    
---    IsEqual (thePnt1   : Pnt from gp;
---             thePnt2   : Pnt from gp)
---    returns Boolean from Standard;
    
    Commands(DI : in out Interpretor from Draw);
    Commands1(DI : in out Interpretor from Draw);
    Commands2(DI : in out Interpretor from Draw);
    Commands3(DI : in out Interpretor from Draw);

end;
