-- Created on: 1993-10-14
-- Created by: Christian CAILLET
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class ToolTransformationMatrix  from IGESGeom

    ---Purpose : Tool to work on a TransformationMatrix. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses TransformationMatrix from IGESGeom,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolTransformationMatrix;
    ---Purpose : Returns a ToolTransformationMatrix, ready to work


    ReadOwnParams (me; ent : mutable TransformationMatrix;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : TransformationMatrix;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : TransformationMatrix;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a TransformationMatrix <ent>, from
    --           its specific (own) parameters

    OwnCorrect (me; ent : mutable TransformationMatrix) returns Boolean  is static;
    ---Purpose : Sets automatic unambiguous Correction on a TransformationMatrix
    --           (FormNumber if 0 or 1, recomputed according Positive/Negative)

    DirChecker (me; ent : TransformationMatrix) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : TransformationMatrix;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : TransformationMatrix; entto : mutable TransformationMatrix;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : TransformationMatrix;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolTransformationMatrix;
