-- File:	IGESDimen_ToolRadiusDimension.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolRadiusDimension  from IGESDimen

    ---Purpose : Tool to work on a RadiusDimension. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses RadiusDimension from IGESDimen,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolRadiusDimension;
    ---Purpose : Returns a ToolRadiusDimension, ready to work


    ReadOwnParams (me; ent : mutable RadiusDimension;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : RadiusDimension;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : RadiusDimension;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a RadiusDimension <ent>, from
    --           its specific (own) parameters

    DirChecker (me; ent : RadiusDimension) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : RadiusDimension;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : RadiusDimension; entto : mutable RadiusDimension;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : RadiusDimension;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolRadiusDimension;
