-- Created on: 1994-08-26
-- Created by: Frederic MAUPAS
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class MakeAxis2Placement2d from GeomToStep inherits Root from GeomToStep

    ---Purpose: This class implements the mapping between classes 
    --          Axis2Placement from Geom and Ax2, Ax22d from gp, and the class
    --          Axis2Placement2d from StepGeom which describes an
    --          axis2_placement_2d from Prostep. 
   
uses Ax2              from gp,
     Ax22d            from gp,
     Axis2Placement   from Geom,
     Axis2Placement2d from StepGeom
     
raises NotDone from StdFail
     
is 

Create ( A : Ax2 from gp ) returns MakeAxis2Placement2d;

Create ( A : Ax22d from gp ) returns MakeAxis2Placement2d;

--Create ( A : Axis2Placement from Geom ) returns MakeAxis2Placement2d;

Value (me) returns Axis2Placement2d from StepGeom
    raises NotDone
    is static;
    ---C++: return const&

fields

    theAxis2Placement2d : Axis2Placement2d from StepGeom;
    	-- TheOP solution from StepGeom
    	
end MakeAxis2Placement2d;


