-- File:	StepBasic_MassUnit.cdl
-- Created:	Thu Dec 12 15:38:08 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class MassUnit from StepBasic
inherits NamedUnit from StepBasic

    ---Purpose: Representation of STEP entity MassUnit

uses
    DimensionalExponents from StepBasic

is
    Create returns MassUnit from StepBasic;
	---Purpose: Empty constructor

end MassUnit;
