-- Created on: 1998-10-14
-- Created by: Andre LIEUTIER
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class D3 from Plate
---Purpose : define an order 3 derivatives of a 3d valued
--          function of a 2d variable
--         

uses XYZ from gp

is
    Create(duuu,duuv,duvv,dvvv : XYZ from gp) returns D3;
    Create(ref  :  D3  from  Plate) returns D3;

fields
    
    Duuu, Duuv,Duvv,Dvvv : XYZ from gp;

friends
    class GtoCConstraint from Plate,
    class FreeGtoCConstraint from Plate
    
end;
