-- Created on: 1993-06-16
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class ShellFaceSet from TopOpeBRepBuild 
    inherits ShapeSet from TopOpeBRepBuild

---Purpose: a bound is a shell, a boundelement is a face.
-- The ShapeSet stores :
-- - a list of shell (bounds),
-- - a list of face (boundelements) to start reconstructions,
-- - a map of edge giving the list of face incident to an edge.

uses

    Shape from TopoDS,
    Solid from TopoDS,
    AsciiString from TCollection,
    ListOfShape from TopTools
    
is

    Create returns ShellFaceSet from TopOpeBRepBuild; 
    ---Purpose: Creates a ShellFaceSet to build blocks of faces 
    -- connected by edges.

    Create(S : Shape from TopoDS; Addr : Address from Standard = NULL) 
    returns ShellFaceSet from TopOpeBRepBuild; 
    ---Purpose: Creates a ShellFaceSet to build blocks of faces 
    -- connected by edges.

    Solid(me) returns Solid from TopoDS is static;
    ---C++: return const &

    AddShape(me:in out;S:Shape) is redefined;
    AddStartElement(me:in out;S:Shape) is redefined;
    AddElement(me:in out;S:Shape) is redefined;

    DumpSS(me:in out) is redefined;
    SName(me;S:Shape from TopoDS;sb:AsciiString = "";sa:AsciiString = "")
    returns AsciiString from TCollection is redefined;
    SName(me;S:ListOfShape from TopTools;sb:AsciiString = "";sa:AsciiString = "")
    returns AsciiString from TCollection is redefined;
    SNameori(me;S:Shape;sb:AsciiString = "";sa:AsciiString = "")
    returns AsciiString from TCollection is redefined;
    SNameori(me;S:ListOfShape from TopTools;sb:AsciiString = "";sa:AsciiString = "")
    returns AsciiString from TCollection is redefined;

fields

    mySolid : Solid from TopoDS;

end ShellFaceSet from TopOpeBRepBuild;
