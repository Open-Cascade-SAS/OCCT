-- Created on: 1995-10-17
-- Created by: Laurent BOURESCHE
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class BoundWithSurf from GeomFill inherits Boundary from GeomFill 

	---Purpose: Defines a 3d curve as a boundary for a
    	-- GeomFill_ConstrainedFilling algorithm.
    	-- This curve is attached to an existing surface.
    	--  Defines a  constrained boundary for  filling  
 	--          the computations are done with a CurveOnSurf and a
 	--          normals field  defined by the normalized normal to
 	--          the surface along the PCurve.

uses
    Pnt            from gp,
    Vec            from gp,
    Function       from Law,
    CurveOnSurface from Adaptor3d

is

    Create(CurveOnSurf : CurveOnSurface from Adaptor3d;
           Tol3d       : Real from Standard;
    	   Tolang      : Real from Standard)
    returns mutable BoundWithSurf from GeomFill;
    	---Purpose:
    	-- Constructs a boundary object defined by the 3d curve CurveOnSurf.
    	-- The surface to be filled along this boundary will be in the
    	-- tolerance range defined by Tol3d.
    	-- What's more, at each point of CurveOnSurf, the angle
    	-- between the normal to the surface to be filled along this
    	-- boundary, and the normal to the surface on which
    	-- CurveOnSurf lies, must not be greater than TolAng.
    	-- This object is to be used as a boundary for a
    	-- GeomFill_ConstrainedFilling framework.
    	-- Warning
    	-- CurveOnSurf is an adapted curve, that is, an object
    	-- which is an interface between:
    	-- -   the services provided by a curve lying on a surface from the package Geom
    	-- -   and those required of the curve by the computation algorithm which uses it.
    	-- The adapted curve is created in the following way:
    	-- Handle(Geom_Surface) mySurface = ... ;
    	-- Handle(Geom2d_Curve) myParamCurve = ... ;
    	-- // where myParamCurve is a 2D curve in the parametric space of the surface mySurface
    	-- Handle(GeomAdaptor_HSurface)
    	--    Surface = new
    	-- GeomAdaptor_HSurface(mySurface);
    	-- Handle(Geom2dAdaptor_HCurve)
    	--    ParamCurve = new
    	-- Geom2dAdaptor_HCurve(myParamCurve);
    	-- CurveOnSurf = Adaptor3d_CurveOnSurface(ParamCurve,Surface);
    	-- The boundary is then constructed with the CurveOnSurf object:
    	-- Standard_Real Tol = ... ;
    	-- Standard_Real TolAng = ... ;
    	-- myBoundary =  GeomFill_BoundWithSurf (
    	-- CurveOnSurf, Tol, TolAng );  
    
    
    

  Value(me; 
          U : Real from Standard) 
    returns Pnt from gp;

    D1(me; 
       U : Real from Standard; 
       P : out Pnt from gp; 
       V : out Vec from gp) ;

    HasNormals(me)
    returns Boolean from Standard
    is redefined;

    Norm(me; 
         U : Real from Standard)
    returns Vec from gp
    is redefined;
    
    D1Norm(me; 
           U  : Real from Standard;
	   N  : out Vec from gp;
	   DN : out Vec from gp)
    is redefined;
    
    Reparametrize(me           : mutable;
    	    	  First, Last  : Real from Standard;
                  HasDF, HasDL : Boolean from Standard;
                  DF, DL       : Real from Standard;
                  Rev          : Boolean from Standard);
		  
    Bounds(me; First, Last : out Real from Standard);

    IsDegenerated(me) returns Boolean from Standard;

fields

    myConS : CurveOnSurface from Adaptor3d;
    myPar  : Function       from Law;

end BoundWithSurf;

