-- File:        SurfaceStyleSilhouette.cdl
-- Created:     Mon Dec  4 12:02:32 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWSurfaceStyleSilhouette from RWStepVisual

	---Purpose : Read & Write Module for SurfaceStyleSilhouette

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     SurfaceStyleSilhouette from StepVisual,
     EntityIterator from Interface

is

	Create returns RWSurfaceStyleSilhouette;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable SurfaceStyleSilhouette from StepVisual);

	WriteStep (me; SW : in out StepWriter; ent : SurfaceStyleSilhouette from StepVisual);

	Share(me; ent : SurfaceStyleSilhouette from StepVisual; iter : in out EntityIterator);

end RWSurfaceStyleSilhouette;
