-- Created on: 1992-08-21
-- Created by: Christophe MARION
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class BiPnt2D from HLRBRep

    	---Purpose: Contains the colors of a shape.

uses
    Boolean from Standard,
    Real    from Standard,
    Pnt2d   from gp,
    Shape   from TopoDS
    
is
    Create
    returns BiPnt2D from HLRBRep; 
    
    Create(x1,y1,x2,y2         : Real    from Standard;
           S                   : Shape   from TopoDS;
           reg1,regn,outl,intl : Boolean from Standard)
    returns BiPnt2D from HLRBRep; 
    
    P1(me) returns Pnt2d from gp
    	---C++: inline
    	---C++: return const &
    is static;

    P2(me) returns Pnt2d from gp
    	---C++: inline
    	---C++: return const &
    is static;

    Shape(me) returns Shape from TopoDS
    	---C++: inline
    	---C++: return const &
    is static;

    Shape(me : in out; S : Shape from TopoDS)
    	---C++: inline
    is static;

    Rg1Line(me) returns Boolean from Standard
    	---C++: inline
    is static;

    Rg1Line(me : in out; B : Boolean from Standard)
    	---C++: inline
    is static;

    RgNLine(me) returns Boolean from Standard
    	---C++: inline
    is static;

    RgNLine(me : in out; B : Boolean from Standard)
    	---C++: inline
    is static;

    OutLine(me) returns Boolean from Standard
    	---C++: inline
    is static;

    OutLine(me : in out; B : Boolean from Standard)
    	---C++: inline
    is static;

    IntLine(me) returns Boolean from Standard
    	---C++: inline
    is static;

    IntLine(me : in out; B : Boolean from Standard)
    	---C++: inline
    is static;

fields
    myP1    : Pnt2d   from gp;
    myP2    : Pnt2d   from gp;
    myShape : Shape   from TopoDS;
    myFlags : Boolean from Standard;

end BiPnt2D;
