-- Created on: 1996-04-30
-- Created by: cle
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package Storage
    
    	---Purpose: Storage package is used to write and read persistent objects.
    	--     These objects are read and written by a retrieval or storage
    	--  algorithm (Storage_Schema object) in a container (disk, memory,
    	-- network ...). Drivers (FSD_File objects) assign a physical
    	-- container for data to be stored or retrieved.
    	-- The standard procedure for an application in
    	-- reading a container is the following:
    	-- -   open the driver in reading mode,
    	-- -   call the Read function from the schema,
    	--   setting the driver as a parameter. This   function returns 
    	-- an instance of the   Storage_Data class which contains the   data being read,
    	-- -   close the driver.
    	-- The standard procedure for an application in writing a container is the following:
    	-- -   open the driver in writing mode,
    	-- -   create an instance of the Storage_Data   class, then
    	--    add the persistent data to write   with the function AddRoot,
    	-- -   call the function Write from the schema,
    	--   setting the driver and the Storage_Data   instance as parameters,
    	-- -      close the driver. 
   
uses TCollection,
     TColStd,
     MMgt
is
    exception StreamModeError inherits Failure from Standard;
    exception StreamFormatError inherits Failure from Standard;
    exception StreamWriteError inherits Failure from Standard;
    exception StreamReadError inherits Failure from Standard;
	    exception StreamUnknownTypeError inherits StreamReadError from Storage;
    	    exception StreamTypeMismatchError inherits StreamReadError from Storage;
	    exception StreamExtCharParityError inherits StreamReadError from Storage;
	    
    enumeration Error
    is
      VSOk,                 -- no problem
      VSOpenError,          -- while opening the stream
      VSModeError,          -- the stream is opened with a wrong mode for operation 
      VSCloseError,         -- while closing the stream
      VSAlreadyOpen,        -- stream is already opened
      VSNotOpen,            -- stream not opened
      VSSectionNotFound,    -- the section is not found
      VSWriteError,         -- error during writing
      VSFormatError,        -- wrong format error occured while reading
      VSUnknownType,        -- try to read an unknown type
      VSTypeMismatch,       -- try to read a wrong primitive type (read a char while expecting a real)
      VSInternalError,      -- internal error
      VSExtCharParityError, -- problem with 16bit characters, may be a 8bit character is inserted inside 16bit string
      VSWrongFileDriver     -- we try to read a file with a wrong driver (occured while reading header section)
    end;
     	---Purpose: Error codes returned by the ErrorStatus
    	-- function on a Storage_Data set of data during a
    	-- storage or retrieval operation :
    	-- -   Storage_VSOk : no problem has been detected
    	-- -   Storage_VSOpenError : an error has
    	--  occurred when opening the driver
    	-- -   Storage_VSModeError : the driver has not
    	--  been opened in the correct mode
    	-- -   Storage_VSCloseError : an error has
    	--   occurred when closing the driver
    	-- -   Storage_VSAlreadyOpen : the driver is   already open
    	-- -   Storage_VSNotOpen : the driver is not   open
    	-- -   Storage_VSSectionNotFound : a section
    	--   has not been found in the driver
    	-- -   Storage_VSWriteError : an error occurred when writing the driver
    	-- -   Storage_VSFormatError : the file format is wrong
    	-- -   Storage_VSUnknownType : a type is not known from the schema
    	-- -   Storage_VSTypeMismatch : trying to read   a wrong type
    	-- -   Storage_VSInternalError : an internal error  has been detected
    	-- -   Storage_VSExtCharParityError : an error
    	--   has occurred while reading 16 bit characte   
 
    enumeration OpenMode
    is
        VSNone,
    	VSRead,
	VSWrite,
	VSReadWrite
    end;
    	---Purpose:
    	-- Specifies opening modes for a file:
    	-- -   Storage_VSNone : no mode is specified
    	-- -   Storage_VSRead : the file is open for  reading operations
    	-- -   Storage_VSWrite : the file is open for writing operations
    	-- -   Storage_VSReadWrite : the file is open
    	--   for both reading and writing operations.

    enumeration SolveMode
    is
    	AddSolve,
	WriteSolve,
	ReadSolve
    end;
    
    imported BucketOfPersistent;
    
    imported Position; -- typedef long
    
    deferred class BaseDriver;

    deferred class CallBack;
      class DefaultCallBack;
	  
    class HeaderData;
          class Data;
	  
    class TypeData;

    class RootData;
    class Root;
    
    class Schema;
        
    imported SeqOfRoot;
    
    imported transient class HSeqOfRoot;

    -- PRIVATE
    
    private class InternalData;
    private class stCONSTclCOM;

    private class TypedCallBack;
    
    imported PType;			

    imported MapOfPers;

    imported DataMapIteratorOfMapOfPers;
        
    imported MapOfCallBack;
        
    imported DataMapIteratorOfMapOfCallBack;
  							  
    imported ArrayOfCallBack;
    imported transient class HArrayOfCallBack;
 
    imported ArrayOfSchema;
    imported transient class HArrayOfSchema;
    
    imported PArray;  
    imported transient class HPArray;
    
    -- METHODS
    
    Version returns AsciiString from TCollection;
    ---Purpose: returns the version of Storage's read/write routines

end;
