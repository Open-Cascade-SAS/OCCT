-- Created by: Peter KURNEV
-- Copyright (c) 2010-2014 OPEN CASCADE SAS
-- Copyright (c) 2007-2010 CEA/DEN, EDF R&D, OPEN CASCADE
-- Copyright (c) 2003-2007 OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN, CEDRAT,
--                         EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class IteratorSI from BOPDS  
    inherits Iterator from BOPDS

---Purpose:  
    -- The class BOPDS_IteratorSI is  
    --  1.to compute self-intersections between BRep sub-shapes  
    --    of each argument of an operation (see the class BOPDS_DS)
    --    in terms of theirs bounding boxes           
    --  2.provides interface to iterare the pairs of  
    --    intersected sub-shapes of given type 

uses  
    BaseAllocator from BOPCol 

is 
    Create   
    returns IteratorSI from BOPDS;
    ---C++: alias "Standard_EXPORT virtual ~BOPDS_IteratorSI();"   
    ---Purpose:  
    --- Empty contructor  
    ---   
 
    Create (theAllocator: BaseAllocator from BOPCol)  
    returns IteratorSI from BOPDS;
     ---Purpose:  
    ---  Contructor    
    ---  theAllocator - the allocator to manage the memory     
    --- 
    Intersect(me:out) 
    is redefined protected;  

    UpdateByLevelOfCheck(me:out; 
      theLevel: Integer from Standard); 
    ---Purpose:  Updates the lists of possible intersections  
    --           according to the value of <theLevel>.
    --           It defines which interferferences will be checked: 
    --           0 - only V/V; 
    --           1 - V/V and V/E; 
    --           2 - V/V, V/E and E/E; 
    --           3 - V/V, V/E, E/E and V/F;
    --           4 - V/V, V/E, E/E, V/F and E/F; 
    --           other - all interferences.
 
end IteratorSI;
