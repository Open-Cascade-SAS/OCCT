-- Created on: 2000-05-10
-- Created by: Andrey BETENEV
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1

class GroupRelationship from StepBasic
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity GroupRelationship

uses
    HAsciiString from TCollection,
    Group from StepBasic

is
    Create returns GroupRelationship from StepBasic;
	---Purpose: Empty constructor

    Init (me: mutable; aName: HAsciiString from TCollection;
                       hasDescription: Boolean;
                       aDescription: HAsciiString from TCollection;
                       aRelatingGroup: Group from StepBasic;
                       aRelatedGroup: Group from StepBasic);
	---Purpose: Initialize all fields (own and inherited)

    Name (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Name
    SetName (me: mutable; Name: HAsciiString from TCollection);
	---Purpose: Set field Name

    Description (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Description
    SetDescription (me: mutable; Description: HAsciiString from TCollection);
	---Purpose: Set field Description
    HasDescription (me) returns Boolean;
	---Purpose: Returns True if optional field Description is defined

    RelatingGroup (me) returns Group from StepBasic;
	---Purpose: Returns field RelatingGroup
    SetRelatingGroup (me: mutable; RelatingGroup: Group from StepBasic);
	---Purpose: Set field RelatingGroup

    RelatedGroup (me) returns Group from StepBasic;
	---Purpose: Returns field RelatedGroup
    SetRelatedGroup (me: mutable; RelatedGroup: Group from StepBasic);
	---Purpose: Set field RelatedGroup

fields
    theName: HAsciiString from TCollection;
    theDescription: HAsciiString from TCollection; -- optional
    theRelatingGroup: Group from StepBasic;
    theRelatedGroup: Group from StepBasic;
    defDescription: Boolean; -- flag "is Description defined"

end GroupRelationship;
