-- Created on: 1991-01-14
-- Created by: Arnaud BOUZY
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Sum from Expr

inherits PolyExpression from Expr

uses GeneralExpression from Expr,
    AsciiString from TCollection,
    NamedUnknown from Expr,
    Array1OfNamedUnknown from Expr,
    Array1OfReal from TColStd,
    SequenceOfGeneralExpression from Expr

raises OutOfRange from Standard,
    NumericError from Standard,
    NotEvaluable from Expr

is

    Create(exps : SequenceOfGeneralExpression)
    ---Purpose: Creates the sum of all the members of sequence <exps>.
    returns mutable Sum;

    Create(exp1,exp2 : GeneralExpression)
    ---Purpose: Creates the sum of <exp1> and <exp2>.
    returns mutable Sum;

    ShallowSimplified(me) 
    ---Purpose: Returns a GeneralExpression after a simplification 
    --          of the arguments of <me>.
    returns any GeneralExpression
    raises NumericError;

    Copy(me)
    ---Purpose: Returns a copy of <me> having the same unknowns and functions.
    returns mutable like me;
    
    IsIdentical(me; Other : GeneralExpression)
    ---Purpose: Tests if <me> and <Other> define the same expression.
    --          This method does not include any simplification before
    --          testing.
    returns Boolean;

    IsLinear(me)
    returns Boolean;

    Derivative(me; X : NamedUnknown)
    ---Purpose: Returns the derivative on <X> unknown of <me>. 
    returns any GeneralExpression;

    NDerivative(me; X : NamedUnknown; N : Integer)
    ---Purpose: Returns the <N>-th derivative on <X> unknown of <me>.
    --          Raises OutOfRange if <N> <= 0
    returns any GeneralExpression
    raises OutOfRange
    is redefined;

    Evaluate(me; vars : Array1OfNamedUnknown; vals : Array1OfReal)
    ---Purpose: Returns the value of <me> (as a Real) by 
    --          replacement of <vars> by <vals>.
    --          Raises NotEvaluable if <me> contains NamedUnknown not 
    --          in <vars> or NumericError if result cannot be computed.
    returns Real
    raises NotEvaluable,NumericError;

    String(me)
    ---Purpose: returns a string representing <me> in a readable way.
    returns AsciiString;

end Sum;
