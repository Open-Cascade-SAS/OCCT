-- File:	StepFEA_DummyNode.cdl
-- Created:	Thu Dec 12 17:51:04 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class DummyNode from StepFEA
inherits NodeRepresentation from StepFEA

    ---Purpose: Representation of STEP entity DummyNode

uses
    HAsciiString from TCollection,
    HArray1OfRepresentationItem from StepRepr,
    RepresentationContext from StepRepr,
    FeaModel from StepFEA

is
    Create returns DummyNode from StepFEA;
	---Purpose: Empty constructor

end DummyNode;
