-- Created on: 1993-02-22
-- Created by: Philippe DAUTRY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Parabola from PGeom
inherits Conic from PGeom 

        --- Purpose :
        --  Defines the parabola in the parameterization range  :
        --  ]-infinite,+infinite[
        --  
	--  See Also : Parabola from Geom.

uses  Ax2 from gp 

is


  Create returns mutable Parabola from PGeom;
        ---Purpose : Creates a parabola with default values.
    	---Level: Internal 


  Create (aPosition : Ax2 from gp; aFocalLength : Real)
    returns mutable Parabola from PGeom;
	---Purpose : Creates a Parabola with <aPosition> and <aFocalLength>
	--         as field values.
    	---Level: Internal 


  FocalLength (me : mutable; aFocalLength : Real);
        ---Purpose :   Set the value  of   the  field focalLength with
        --         <aFocalLength>.
    	---Level: Internal 


  FocalLength (me)  returns Real;
	---Purpose : Retruns the value of the field focalLength.
    	---Level: Internal 


fields

  focalLength : Real;

end;
