-- Created on: 1991-12-13
-- Created by: Christophe MARION
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package Intrv 

	---Purpose: 
uses
    Standard,
    TCollection

is
                                 --                  other
    enumeration Position is      --      me     **------------***
    	Before,                  --    **---*
	JustBefore,              --    **--------*
	OverlappingAtStart,      --    **--------------*
	JustEnclosingAtEnd,      --    **----------------------*
	Enclosing,               --    **------------------------------*
	JustOverlappingAtStart,  --              *---------*
	Similar,                 --              *-------------*
	JustEnclosingAtStart,    --              *---------------------*
	Inside,                  --                    *---*
	JustOverlappingAtEnd,    --                    *-------*
    	OverlappingAtEnd,        --                    *---------------*
	JustAfter,               --                            *-------*
	After                    --                                 *--*
    end Position;
    
    class Interval;
    class Intervals;
    class SequenceOfInterval instantiates Sequence from TCollection(Interval);
    
end Intrv;
