-- Created on: 1997-10-29
-- Created by: Roman BORISOV
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


package FEmTool 

	---Purpose: Tool to Finite Element methods
	
	---Level: Advanced
uses  
    TCollection, 
    TColStd, 
    math, 
    PLib,
    GeomAbs 
is  
                   
    class  Assembly; 
      
    ---Purpose: To define Criterium (or  Energy) on finite element   
    deferred  class  ElementaryCriterion;     
    class  LinearTension;      
    class  LinearFlexion;      
    class  LinearJerk;
      
    ---Purpose: To define sparse Matrix          
    deferred  class  SparseMatrix; 
    class  ProfileMatrix;

    ---Purpose: Do define one curves with Finite Element
    class  Curve;   
    
    ---Purpose:  To  define  set  of  functions  for  calculating  matrix 
    --	         elements  of  RefMatrix  by  Gauss  integration. 
    class  ElementsOfRefMatrix; 
     
    --  instantiate  classes  
      
    ---Purpose:  To define the  table  [Freedom's degree] [Dimension,Element]
    --           which gives Index  of Freedom's degree in the
    --           assembly problem.
   
    class  AssemblyTable
    instantiates Array2 from TCollection (HArray1OfInteger from  TColStd);     
    class  HAssemblyTable   
    instantiates HArray2 from TCollection (HArray1OfInteger from  TColStd,
    	    	    	                   AssemblyTable  from  FEmTool); 
					    
    ---Purpose:  To  define  list  of  segments with  non-zero  coefficients   
    --           of constraint 
        
    class  ListOfVectors  
    instantiates  List  from  TCollection  (HArray1OfReal  from  TColStd); 

    ---Purpose:  To  define  sequence  of  constraints 
    
    class  SeqOfLinConstr  
    instantiates  Sequence  from  TCollection  (ListOfVectors  from  FEmTool); 
      
     
end FEmTool;
