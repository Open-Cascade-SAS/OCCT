-- Created on: 1998-03-23
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class C2DF from TopOpeBRepTool

uses

    Curve from Geom2d,
    Face from TopoDS

is

    Create returns C2DF from TopOpeBRepTool;    
    Create(PC : Curve from Geom2d; f2d,l2d,tol : Real; F : Face from TopoDS) 
    returns C2DF from TopOpeBRepTool;
    SetPC(me : in out;PC : Curve from Geom2d; f2d,l2d,tol : Real);
    SetFace(me : in out; F : Face from TopoDS);
    PC(me; f2d,l2d,tol : out Real) returns Curve from Geom2d;
    ---C++: return const &
    Face(me) returns Face from TopoDS;
    ---C++: return const &
    IsPC(me;PC:Curve from Geom2d) returns Boolean;
    IsFace(me;F:Face from TopoDS) returns Boolean;
    
fields
    
    myPC : Curve from Geom2d;
    myf2d,myl2d,mytol : Real;
    myFace : Face from TopoDS;
    
end C2DF;
