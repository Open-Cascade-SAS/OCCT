-- Created on: 2007-05-29
-- Created by: Vlad Romashko
-- Copyright (c) 2007-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ReferenceList from PDataStd inherits Attribute from PDF

uses 

    HExtendedString from PCollection,
    HArray1OfExtendedString from PColStd

is

    Create 
    returns mutable ReferenceList from PDataStd;

    Init (me : mutable; 
    	  lower, upper : Integer from Standard);

    SetValue (me: mutable; 
    	      index : Integer from Standard; 
    	      value : HExtendedString from PCollection);

    Value (me;  
    	   index : Integer from Standard) 
    returns HExtendedString from PCollection;

    Lower (me) 
    returns Integer from Standard;      

    Upper (me) 
    returns Integer from Standard;   


fields

    myValue     :  HArray1OfExtendedString from PColStd;


end ReferenceList;
