-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package StepElement


uses

    TCollection,
    TColStd,
    MMgt,
    StepData,
    StepBasic,
    StepRepr

is 

    enumeration ElementOrder is 
	Linear,
	Quadratic,
	Cubic
    end;

    enumeration EnumeratedCurveElementPurpose is 
	Axial,
	YYBending,
	ZZBending,
	Torsion,
	XYShear,
	XZShear,
	Warping
    end;

    enumeration EnumeratedCurveElementFreedom is 
	XTranslation,
	YTranslation,
	ZTranslation,
	XRotation,
	YRotation,
	ZRotation,
	Warp,
	None
    end;

    enumeration UnspecifiedValue is 
	Unspecified
    end;

    enumeration ElementVolume is 
	Volume
    end;

    enumeration CurveEdge is 
	ElementEdge
    end;

    enumeration EnumeratedSurfaceElementPurpose is 
	MembraneDirect,
	MembraneShear,
	BendingDirect,
	BendingTorsion,
	NormalToPlaneShear
    end;

    enumeration Element2dShape is 
	Quadrilateral,
	Triangle
    end;

    enumeration EnumeratedVolumeElementPurpose is 
	StressDisplacement
    end;

    enumeration Volume3dElementShape is 
	Hexahedron,
	Wedge,
	Tetrahedron,
	Pyramid
    end;
    
    

   class AnalysisItemWithinRepresentation;
   class Curve3dElementDescriptor;
   class CurveElementEndReleasePacket;
   class CurveElementFreedom;
     class CurveElementFreedomMember;
   class CurveElementPurpose;
     class CurveElementPurposeMember;
   class CurveElementSectionDefinition;
   class CurveElementSectionDerivedDefinitions;
   class ElementAspect;
     class ElementAspectMember;
   class ElementDescriptor;
   class ElementMaterial;
   class MeasureOrUnspecifiedValue;
     class MeasureOrUnspecifiedValueMember;
   class Surface3dElementDescriptor;
   class SurfaceElementProperty;
   class SurfaceElementPurpose;
     class SurfaceElementPurposeMember;
   class SurfaceSection;
   class SurfaceSectionField;
   class SurfaceSectionFieldConstant;
   class SurfaceSectionFieldVarying;
   class UniformSurfaceSection;
   class Volume3dElementDescriptor;
   class VolumeElementPurpose;
     class VolumeElementPurposeMember;
	
	
--- Instantiations

imported Array2OfCurveElementPurposeMember;
imported transient class HArray2OfCurveElementPurposeMember;

imported Array2OfSurfaceElementPurposeMember;
imported transient class HArray2OfSurfaceElementPurposeMember;

imported Array1OfVolumeElementPurposeMember;
imported transient class HArray1OfVolumeElementPurposeMember;

imported Array2OfSurfaceElementPurpose;
imported transient class HArray2OfSurfaceElementPurpose;

imported Array1OfMeasureOrUnspecifiedValue;
imported transient class HArray1OfMeasureOrUnspecifiedValue;

imported Array1OfSurfaceSection;
imported transient class HArray1OfSurfaceSection;

imported Array1OfVolumeElementPurpose;
imported transient class HArray1OfVolumeElementPurpose;

imported Array1OfCurveElementEndReleasePacket;
imported transient class HArray1OfCurveElementEndReleasePacket;

imported Array1OfCurveElementSectionDefinition;
imported transient class HArray1OfCurveElementSectionDefinition;


imported SequenceOfElementMaterial;
imported transient class HSequenceOfElementMaterial;

imported SequenceOfCurveElementSectionDefinition;
imported transient class HSequenceOfCurveElementSectionDefinition;

imported SequenceOfCurveElementPurposeMember;
imported transient class HSequenceOfCurveElementPurposeMember;
imported Array1OfHSequenceOfCurveElementPurposeMember;
imported transient class HArray1OfHSequenceOfCurveElementPurposeMember;

imported SequenceOfSurfaceElementPurposeMember;
imported transient class HSequenceOfSurfaceElementPurposeMember;
imported Array1OfHSequenceOfSurfaceElementPurposeMember;
imported transient class HArray1OfHSequenceOfSurfaceElementPurposeMember;


end;
