-- File:        PreDefinedTextFont.cdl
-- Created:     Fri Dec  1 11:11:25 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class PreDefinedTextFont from StepVisual 

inherits PreDefinedItem from StepVisual 

uses

	HAsciiString from TCollection
is

	Create returns mutable PreDefinedTextFont;
	---Purpose: Returns a PreDefinedTextFont


end PreDefinedTextFont;
