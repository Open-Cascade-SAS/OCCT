-- File:        GaussLeastSquare.cdl
-- Created:     Mon May 13 16:24:37 1991
-- Author:      Laurent PAINNOT
--              <lpa@topsn3>
---Copyright:    Matra Datavision 1991, 1992


class GaussLeastSquare from math
    ---Purpose:
    -- This class implements the least square solution of a set of
    -- n linear equations of m unknowns (n >= m) using the gauss LU
    -- decomposition algorithm.
    -- This algorithm is more likely subject to numerical instability
    --  than math_SVD.


uses Matrix from math, 
     Vector from math, 
     IntegerVector from math,
     OStream from Standard

raises NotDone from StdFail,
       DimensionError from Standard

is

    Create(A: Matrix; MinPivot: Real = 1.0e-20)
    ---Purpose: Given an input n X m matrix A with n >= m this constructor 
    --          performs the LU decomposition with partial pivoting
    --          (interchange of rows) of the matrix AA = A.Transposed() * A;
    -- 	        This LU decomposition is stored internally and may be used 
    -- 	        to do subsequent calculation.
    --          If the largest pivot found is less than MinPivot the matrix <A>
    --          is considered as singular.

    returns GaussLeastSquare;
    
    
    IsDone(me)
    	---Purpose: Returns true if the computations are successful, otherwise returns false.e
    	---C++: inline
    returns Boolean
    is static;
    
    
    Solve(me; B: in Vector; X: out Vector)
    ---Purpose: Given the input Vector <B> this routine solves the set 
    --          of linear equations A . X = B. 
    --          Exception NotDone is raised if the decomposition of A was 
    --          not done successfully.
    --          Exception DimensionError is raised if the range of B Inv is 
    --          not equal to the rowrange of A.
    --          Exception DimensionError is raised if the range of X Inv is
    --          not equal to the colrange of A.

    raises NotDone,
    	   DimensionError
    is static;


    Dump(me; o: in out OStream)
    	---Purpose: Prints on the stream o information on the current state 
    	--          of the object.
    	--          Is used to redefine the operator <<.

    is static;

   	
fields

Done:      Boolean;
Singular:  Boolean is protected;
LU:        Matrix is protected;
A2 :       Matrix is protected;
Index:     IntegerVector is protected;
D:         Real is protected;

    
end GaussLeastSquare;
