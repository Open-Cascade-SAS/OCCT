-- Created on: 1999-03-08
-- Created by: Fabrice SERVANT
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class ArrayOfTriangles from IntPolyh

uses
    
    Triangle from IntPolyh


is


    Create;
    
    Create(nn : Integer from Standard) ; 
    
    Init(me: in out; nn: Integer from Standard) 
    is static;

    GetN(me)
    returns Integer from Standard
    ---C++: return const
    is static;
    
    NbTriangles(me)
    returns Integer from Standard
    ---C++: return const
    is static;
    
    SetNbTriangles(me : in out; endaot: Integer from Standard)
    is static;
    
    IncNbTriangles(me: in out)
    is static;
    
    Value(me; nn: Integer from Standard)
    	---C++: alias operator [] 
    	---C++: return const &      
    returns Triangle from IntPolyh
    is static;
    
    ChangeValue(me: in out;  nn: Integer from Standard)
    	---C++: alias operator [] 
    	---C++: return &
    returns Triangle from IntPolyh 
    is static;
    
    Copy(me: in out; Other : ArrayOfTriangles from IntPolyh)
    	---C++: alias operator =
    	---C++: return &
    returns ArrayOfTriangles from IntPolyh
    is static;
    
    Destroy(me:in out)
    	---C++: alias ~
    is static;
    
    Dump(me) 
    is static;
    
    DumpFleches(me) 
    is static;

     	
fields

    n, fintt : Integer from Standard;
    ptr      : Address from Standard;
    
end ArrayOfTriangles from IntPolyh;
