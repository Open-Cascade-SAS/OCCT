-- Created on: 1999-11-26
-- Created by: Andrey BETENEV
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0

class ConfigurationDesign from StepRepr
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity ConfigurationDesign

uses
    ConfigurationItem from StepRepr,
    ConfigurationDesignItem from StepRepr

is
    Create returns ConfigurationDesign from StepRepr;
	---Purpose: Empty constructor

    Init (me: mutable; aConfiguration: ConfigurationItem from StepRepr;
                       aDesign: ConfigurationDesignItem from StepRepr);
	---Purpose: Initialize all fields (own and inherited)

    Configuration (me) returns ConfigurationItem from StepRepr;
	---Purpose: Returns field Configuration
    SetConfiguration (me: mutable; Configuration: ConfigurationItem from StepRepr);
	---Purpose: Set field Configuration

    Design (me) returns ConfigurationDesignItem from StepRepr;
	---Purpose: Returns field Design
    SetDesign (me: mutable; Design: ConfigurationDesignItem from StepRepr);
	---Purpose: Set field Design

fields
    theConfiguration: ConfigurationItem from StepRepr;
    theDesign: ConfigurationDesignItem from StepRepr;

end ConfigurationDesign;
