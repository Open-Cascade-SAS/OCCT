-- File:	MakeTrimmedCone.cdl
-- Created:	Mon Sep 28 11:52:10 1992
-- Author:	Remi GILET
--		<reg@sdsun2>
---Copyright:	 Matra Datavision 1992

class MakeTrimmedCone from GC inherits Root from GC

    --- Purpose: Implements construction algorithms for a trimmed
    -- cone limited by two planes orthogonal to its axis. The
    -- result is a Geom_RectangularTrimmedSurface surface.
    -- A MakeTrimmedCone provides a framework for:
    -- -   defining the construction of the trimmed cone,
    -- -   implementing the construction algorithm, and
    -- -   consulting the results. In particular, the Value
    --   function returns the constructed trimmed cone.
uses Pnt                       from gp,
     Ax1                       from gp,
     Lin                       from gp,
     Cone                      from gp,
     RectangularTrimmedSurface from Geom,
     Real                      from Standard

raises NotDone from StdFail

is

Create(P1,P2,P3,P4 : Pnt from gp ) returns MakeTrimmedCone;
    ---Purpose: Make a RectangularTrimmedSurface <TheCone> from Geom
    --          It is trimmed by P3 and P4.
    --          Its axis is <P1P2> and the radius of its base is
    --          the distance between <P3> and <P1P2>.
    --          The distance between <P4> and <P1P2> is the radius of 
    --          the section passing through <P4>.
    --          An error iss raised if <P1>,<P2>,<P3>,<P4> are 
    --          colinear or if <P3P4> is perpendicular to <P1P2> or 
    --          <P3P4> is colinear to <P1P2>.

Create(P1,P2 : Pnt  from gp      ;
       R1,R2 : Real from Standard) returns MakeTrimmedCone;
    ---Purpose : Make a RectangularTrimmedSurface from Geom <TheCone> 
    --           from a cone and trimmed by two points P1 and P2 and 
    --           the two radius <R1> and <R2> of the sections passing 
    --           through <P1> an <P2>.
    -- Warning
    -- If an error occurs (that is, when IsDone returns
    -- false), the Status function returns:
    -- -   gce_ConfusedPoints if points P1 and P2, or P3 and P4, are coincident;
    -- -   gce_NullAngle if:
    --   -   the lines joining P1 to P2 and P3 to P4 are parallel, or
    -- -   R1 and R2 are equal (i.e. their difference is less than gp::Resolution());
    -- -   gce_NullRadius if:
    --   -   the line joining P1 to P2 is perpendicular to the line joining P3 to P4, or
    --   -   the points P1, P2, P3 and P4 are collinear;
    -- -   gce_NegativeRadius if R1 or R2 is negative; or
    -- -   gce_NullAxis if points P1 and P2 are coincident (2nd syntax only).
        
Value(me) returns RectangularTrimmedSurface from Geom
    raises NotDone
    is static;
    ---Purpose: Returns the constructed trimmed cone.
    -- StdFail_NotDone if no trimmed cone is constructed.
    ---C++: return const&

Operator(me) returns RectangularTrimmedSurface from Geom
    is static;
    ---C++: return const&
    ---C++: alias "Standard_EXPORT operator Handle_Geom_RectangularTrimmedSurface() const;"

fields

    TheCone : RectangularTrimmedSurface from Geom;
    --The solution from Geom.
    
end MakeTrimmedCone;
