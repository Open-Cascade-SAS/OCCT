-- Created on: 1992-04-14
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

generic class Segment from IntStart

    (TheVertex    as any;
     TheArc       as any;
     ThePathPoint as any) -- as PathPoint from IntStart (TheVertex,TheArc)

	---Purpose: This class defines the intersection between two implicit
	--          surfaces A and B, when this intersection is a part of an 
	--          arc of restriction .
	--          It can be bounded or  semi infinite;
	--          the extremities of these curves are vertices(ThepathPoint).


raises DomainError from Standard

is

    Create

        ---Purpose: Empty constructor.

    	returns Segment;


    SetValue(me: in out; A: TheArc)
	     
	---Purpose: Defines the concerned arc.

	---C++: inline

    	is static;
	

    SetLimitPoint(me: in out; V: ThePathPoint; First: Boolean)
    
	---Purpose: Defines the first point or the last point,
	--          depending on the value of the boolean First.

    	is static;


    Curve(me)
    
    	---Purpose: Returns the geometric curve on the surface 's domain
    	--          which is solution.

    	returns any TheArc
	---C++: return const&
	---C++: inline

    	is static;
  

    HasFirstPoint(me)
    
	---Purpose: Returns True if there is a vertex (ThePathPoint) defining
	--          the lowest valid parameter on the arc.
    
    	returns Boolean from Standard
	---C++: inline

	is static;


    FirstPoint(me)

    	---Purpose: Returns the first point.
	
    	returns ThePathPoint
	---C++: return const&	
	---C++: inline

	raises DomainError from Standard
	
	is static;



    HasLastPoint(me)
    
	---Purpose: Returns True if there is a vertex (ThePathPoint) defining
	--          the greatest valid parameter on the arc.
    
    	returns Boolean from Standard
	---C++: inline

	is static;


    LastPoint(me)

    	---Purpose: Returns the last point.
	
    	returns ThePathPoint
	---C++: return const&	
	---C++: inline

	raises DomainError from Standard
	
	is static;



fields

    arc   : TheArc;
    hasfp : Boolean from Standard;
    thefp : ThePathPoint;
    haslp : Boolean from Standard;
    thelp : ThePathPoint;

end Segment;
