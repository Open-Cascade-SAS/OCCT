-- Created on: 2000-05-10
-- Created by: Andrey BETENEV
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1

class AppliedGroupAssignment from StepAP214
inherits GroupAssignment from StepBasic

    ---Purpose: Representation of STEP entity AppliedGroupAssignment

uses
    Group from StepBasic,
    HArray1OfGroupItem from StepAP214

is
    Create returns AppliedGroupAssignment from StepAP214;
	---Purpose: Empty constructor

    Init (me: mutable; aGroupAssignment_AssignedGroup: Group from StepBasic;
                       aItems: HArray1OfGroupItem from StepAP214);
	---Purpose: Initialize all fields (own and inherited)

    Items (me) returns HArray1OfGroupItem from StepAP214;
	---Purpose: Returns field Items
    SetItems (me: mutable; Items: HArray1OfGroupItem from StepAP214);
	---Purpose: Set field Items

fields
    theItems: HArray1OfGroupItem from StepAP214;

end AppliedGroupAssignment;
