-- Created on: 1995-03-09
-- Created by: Laurent PAINNOT
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Polygon3D from DrawTrSurf inherits Drawable3D from Draw

    	---Purpose: Used to display a 3d polygon.
    	--          
    	--          Optional display of nodes.


uses Polygon3D   from Poly,
     Display     from Draw,
     Interpretor from Draw,
     OStream

is

    Create(P: Polygon3D from Poly)
    returns mutable Polygon3D from DrawTrSurf;
    
    Polygon3D(me) returns Polygon3D from Poly;
    
    ShowNodes(me: mutable; B: Boolean);
    
    ShowNodes(me) returns Boolean;
    
    DrawOn(me; dis: in out Display);
    
    Copy(me) returns mutable Drawable3D from Draw
    is redefined;
	---Purpose: For variable copy.


    Dump(me; S : in out OStream)
    is redefined;
	---Purpose: For variable dump.

    Whatis(me; I : in out Interpretor from Draw)
    is redefined;
	---Purpose: For variable whatis command. Set  as a result  the
	--          type of the variable.


fields

    myPolygon3D:  Polygon3D from Poly;
    myNodes:      Boolean;

end Polygon3D;
