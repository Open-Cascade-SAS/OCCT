-- Created on: 1993-01-09
-- Created by: CKY / Contract Toubro-Larsen ( Anand NATRAJAN )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class AssocGroupType from IGESBasic  inherits IGESEntity

        ---Purpose: defines AssocGroupType, Type <406> Form <23>
        --          in package IGESBasic
        --          Used to assign an unambiguous identification to a Group
        --          Associativity.

uses

        HAsciiString from TCollection

is

        Create returns mutable AssocGroupType;

        -- Specific Methods pertaining to the class

        Init (me : mutable; nbDataFields, aType : Integer; 
              aName : HAsciiString );
        ---Purpose : This method is used to set the fields of the class
        --           AssocGroupType
        --       - nbDataFields : number of parameter data fields = 2
        --       - aType        : type of attached associativity
        --       - aName        : identifier of associativity of type AType

        NbData (me) returns Integer;
        ---Purpose : returns the number of parameter data fields, always = 2

        AssocType (me) returns Integer;
        ---Purpose : returns the type of attached associativity

        Name (me) returns HAsciiString from TCollection;
        ---Purpose : returns identifier of instance of specified associativity

fields

--
-- Class    : IGESBasic_AssocGroupType
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class AssocGroupType.
--
-- Reminder : A AssocGroupType instance is defined by :
--            - the number of parameter data fields, always = 2
--            - the type of attached associativity
--            - the identifier of instance of specified associativity

        theNbData : Integer;
        theType   : Integer;
        theName   : HAsciiString from TCollection;

end AssocGroupType;
