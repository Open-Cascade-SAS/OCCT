-- Created on: 2002-12-15
-- Created by: data exchange team
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class ProductDefinitionFormationRelationship from StepBasic
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity ProductDefinitionFormationRelationship

uses
    HAsciiString from TCollection,
    ProductDefinitionFormation from StepBasic

is
    Create returns ProductDefinitionFormationRelationship from StepBasic;
	---Purpose: Empty constructor

    Init (me: mutable; aId: HAsciiString from TCollection;
                       aName: HAsciiString from TCollection;
                       aDescription: HAsciiString from TCollection;
                       aRelatingProductDefinitionFormation: ProductDefinitionFormation from StepBasic;
                       aRelatedProductDefinitionFormation: ProductDefinitionFormation from StepBasic);
	---Purpose: Initialize all fields (own and inherited)

    Id (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Id
    SetId (me: mutable; Id: HAsciiString from TCollection);
	---Purpose: Set field Id

    Name (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Name
    SetName (me: mutable; Name: HAsciiString from TCollection);
	---Purpose: Set field Name

    Description (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Description
    SetDescription (me: mutable; Description: HAsciiString from TCollection);
	---Purpose: Set field Description

    RelatingProductDefinitionFormation (me) returns ProductDefinitionFormation from StepBasic;
	---Purpose: Returns field RelatingProductDefinitionFormation
    SetRelatingProductDefinitionFormation (me: mutable; RelatingProductDefinitionFormation: ProductDefinitionFormation from StepBasic);
	---Purpose: Set field RelatingProductDefinitionFormation

    RelatedProductDefinitionFormation (me) returns ProductDefinitionFormation from StepBasic;
	---Purpose: Returns field RelatedProductDefinitionFormation
    SetRelatedProductDefinitionFormation (me: mutable; RelatedProductDefinitionFormation: ProductDefinitionFormation from StepBasic);
	---Purpose: Set field RelatedProductDefinitionFormation

fields
    theId: HAsciiString from TCollection;
    theName: HAsciiString from TCollection;
    theDescription: HAsciiString from TCollection;
    theRelatingProductDefinitionFormation: ProductDefinitionFormation from StepBasic;
    theRelatedProductDefinitionFormation: ProductDefinitionFormation from StepBasic;

end ProductDefinitionFormationRelationship;
