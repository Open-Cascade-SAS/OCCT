-- Created on: 1991-03-07
-- Created by: Denis Pascal
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



package GraphTools 

    ---Purpose: This package <GraphTools> provides  algorithms working
    --          on a directed graph.  Those algorithms are generic for
    --          user (Graph and Vertex)  data, and tool classes.


uses Standard,
     MMgt,
     TCollection,
     TColStd
     
is


    class ListOfSequenceOfInteger instantiates List from TCollection
                         (SequenceOfInteger from TColStd);

-- Requirements
-- ============

-- Data
--  Vertex
--  Graph
-- Tools
    generic class GraphIterator;
    generic class VertexIterator;

-- Services (Algorithms) 
-- =====================
    
    
    ---Purpose: Depth First Search (DFS)
    
    generic class DFSIterator,
                  DFSMap;


    ---Purpose: Breath First Search (BFS)

    generic class BFSIterator,
                  BFSMap;

		  
    ---Purpose: Sorted Strong Components (SC)

    generic class SortedStrgCmptsFromIterator,
                  SCMap;
		  
    generic class SortedStrgCmptsIterator;


    ---Purpose: Topological Sort (TS)

    class TSNode;

    generic class TopologicalSortFromIterator,
                  TSMap;  
		  
    generic class TopologicalSortIterator;
    
    
    ---Purpose: Connected Vertices (CV)

    generic class ConnectedVerticesFromIterator,
                  CVMap,
    	    	  ConnectMap;
		 
    generic class ConnectedVerticesIterator;


    ---Purpose: Reduced Graph (RG)
    
    class RGNode;
    
    class SC;
    
    class SCList instantiates List from TCollection
                (SC from GraphTools);

    generic class ReducedGraph,
		  RGMap,
		  SortedSCIterator,
		  AdjSCIterator;

end GraphTools;





