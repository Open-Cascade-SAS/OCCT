-- File:	IGESDraw_ReadWriteModule.cdl
-- Created:	Mon Sep  6 19:22:12 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993



class ReadWriteModule  from IGESDraw   inherits ReadWriteModule from IGESData

    ---Purpose : Defines Draw File Access Module for IGESDraw (specific parts)
    --           Specific actions concern : Read and Write Own Parameters of
    --           an IGESEntity.

uses Transient, FileReaderData,
     IGESEntity, DirPart, IGESReaderData, ParamReader, IGESWriter

raises DomainError

is

    Create returns mutable ReadWriteModule from IGESDraw;
    ---Purpose : Creates a ReadWriteModule & puts it into ReaderLib & WriterLib

    CaseIGES (me; typenum, formnum : Integer) returns Integer;
    ---Purpose : Defines Case Numbers for Entities of IGESDraw

    ReadOwnParams (me; CN : Integer; ent : mutable IGESEntity;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError;
    ---Purpose : Reads own parameters from file for an Entity of IGESDraw

    WriteOwnParams (me; CN : Integer;  ent : IGESEntity;
    	    	    IW : in out IGESWriter);
    ---Purpose : Writes own parameters to IGESWriter

end ReadWriteModule;
