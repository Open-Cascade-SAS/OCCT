-- Created on: 1993-09-06
-- Created by: Christian CAILLET
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ReadWriteModule  from IGESAppli   inherits ReadWriteModule from IGESData

    ---Purpose : Defines basic File Access Module for IGESAppli (specific parts)
    --           Specific actions concern : Read and Write Own Parameters of
    --           an IGESEntity.

uses Transient, FileReaderData,
     IGESEntity, DirPart, IGESReaderData, ParamReader, IGESWriter

raises DomainError

is

    Create returns mutable ReadWriteModule from IGESAppli;
    ---Purpose : Creates a ReadWriteModule & puts it into ReaderLib & WriterLib

    CaseIGES (me; typenum, formnum : Integer) returns Integer;
    ---Purpose : Defines Case Numbers for Entities of IGESAppli

    ReadOwnParams (me; CN : Integer; ent : mutable IGESEntity;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError;
    ---Purpose : Reads own parameters from file for an Entity of IGESAppli

    WriteOwnParams (me; CN : Integer;  ent : IGESEntity;
    	    	    IW : in out IGESWriter);
    ---Purpose : Writes own parameters to IGESWriter

end ReadWriteModule;
