-- Created on: 1994-04-18
-- Created by: Modelistation
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Segment2D from Draw inherits Drawable2D from Draw

	---Purpose: 

uses Pnt2d from gp,
    Color from Draw,
    Display from Draw,
    Interpretor from Draw

is

    Create(p1,p2 : Pnt2d; col : Color)
    returns Segment2D;
    
    DrawOn(me; dis : in out Display);
    
    First(me) returns Pnt2d from gp
	---C++: return const&
    is static;

    First(me : mutable; P : Pnt2d from gp)
    is static;

    Last(me) returns Pnt2d from gp
	---C++: return const&
    is static;

    Last(me : mutable; P : Pnt2d from gp)
    is static;
	
    Dump(me; S : in out OStream)
    is redefined;

    Whatis(me; I : in out Interpretor from Draw)
    is redefined;

fields

    myFirst : Pnt2d;
    myLast  : Pnt2d;
    myColor : Color;
    
end Segment2D;
