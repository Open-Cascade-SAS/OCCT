-- File:        SiUnit.cdl
-- Created:     Mon Dec  4 12:02:31 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWSiUnit from RWStepBasic

	---Purpose : Read & Write Module for SiUnit

uses 
    
    Check from Interface,
    StepReaderData from StepData,
    StepWriter  from StepData,
    SiUnit      from StepBasic,
    SiPrefix    from StepBasic,
    SiUnitName  from StepBasic,
    AsciiString from TCollection

is

    Create returns RWSiUnit;

    ReadStep (me; data: StepReaderData; num: Integer;
	          ach : in out Check;   ent: mutable SiUnit from StepBasic);

    WriteStep (me; SW : in out StepWriter; ent : SiUnit from StepBasic);
    
    DecodePrefix(me; aPrefix: in out SiPrefix from StepBasic;
    	    	     text   : CString from Standard)
    returns Boolean;
    
    DecodeName(me; aName: in out SiUnitName from StepBasic;
    	    	   text   : CString from Standard)
    returns Boolean;
    
    EncodePrefix(me; aPrefix: SiPrefix from StepBasic) returns AsciiString from TCollection;
    
    EncodeName(me; aName: SiUnitName from StepBasic) returns AsciiString from TCollection;

end RWSiUnit;
