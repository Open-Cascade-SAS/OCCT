-- Created on: 1995-05-10
-- Created by: Denis PASCAL
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package TDataStd 

	---Purpose:  This  package  defines   standard attributes for
	--           modelling. 
	-- These allow you to create and modify labels
	-- and attributes for many basic data types.
	-- Standard topological and visualization
	-- attributes have also been created.
	-- To find an attribute attached to a specific label,
	-- you use the GUID of the type of attribute you
	-- are looking for. To do this, first find this
	-- information using the method GetID as follows: Standard_GUID anID =
	-- MyAttributeClass::GetID();
	-- Then, use the method Find for the label as follows:
	-- Standard_Boolean HasAttribute
	-- =
	-- aLabel.Find(anID,anAttribute);
	-- Note
	-- For information on the relations between this
	-- component of OCAF and the others, refer to the OCAF User's Guide.
	
    ---  Category: GUID - AttributeID
    --           2a96b606-ec8b-11d0-bee7-080009dc3333	TDataStd_Integer 
    
    --           2a96b608-ec8b-11d0-bee7-080009dc3333	TDataStd_Name	
    --           2a96b60f-ec8b-11d0-bee7-080009dc3333	TDataStd_Real	
    --           2a96b610-ec8b-11d0-bee7-080009dc3333	TDataStd_Reference
    --           2a96b616-ec8b-11d0-bee7-080009dc3333	TDataStd_Comment  
    --           2a96b61c-ec8b-11d0-bee7-080009dc3333   TDataStd_UAttribute  	
    --           2a96b61d-ec8b-11d0-bee7-080009dc3333   TDataStd_IntegerArray        
    --           2a96b61e-ec8b-11d0-bee7-080009dc3333   TDataStd_RealArray
    --           2a96b624-ec8b-11d0-bee7-080009dc3333   TDataStd_ExtStringArray
    --           2a96b609-ec8b-11d0-bee7-080009dc3333	TDataStd_NoteBook
    --           2a96b61f-ec8b-11d0-bee7-080009dc3333   TDataStd_Directory




uses Standard,
     MMgt,
     TCollection,
     TColStd,
     TDF


is
    enumeration RealEnum is 
        ---Purpose:
	-- The terms of this enumeration define the
	-- semantics of a real number value.       
      SCALAR,
      LENGTH,
      ANGULAR
    end RealEnum;    
                  
    ---Category:  Basic  attributes
    --           ===================


    class Current;

    class Name;
    
    class Comment;
    
    class Integer; 
    
    class IntegerArray;    
    
    class Real;
    
    class RealArray;
    
    class ExtStringArray;

    class UAttribute; 
    
    
    ---Category: Attributes for organization
    --          ============================
    
    class TreeNode;
    pointer PtrTreeNode to TreeNode from TDataStd;  	    
    class ChildNodeIterator;

    class Directory;	
    

    ---Category: Other attributes
    --           ================
          
    class NoteBook;
    
    class Expression;
    
    class Relation;
    
    class Variable; 
    
    class DeltaOnModificationOfIntArray;  
     
    class DeltaOnModificationOfRealArray;  
     
    class DeltaOnModificationOfExtStringArray; 
     
    class DeltaOnModificationOfIntPackedMap; 
     
    class DeltaOnModificationOfByteArray; 
     
      
    -- Extension
    class Tick; 
    
    class AsciiString;  
    
    class IntPackedMap; 

     
    -- Lists:
    class IntegerList; 
    
    class RealList; 
    
    class ExtStringList; 
    
    class BooleanList; 
    
    class ReferenceList;


    -- Arrays:
    class BooleanArray; 
    
    class ReferenceArray; 
    
    class ByteArray;

    class NamedData;         
         					       
    imported ListOfExtendedString;
         					       
    imported ListIteratorOfListOfExtendedString;	 

      
    --  Extension
    imported ListOfByte;
    imported ListIteratorOfListOfByte;

    imported LabelArray1; 
    
    imported transient class HLabelArray1;

    imported DataMapOfStringReal;

    imported DataMapIteratorOfDataMapOfStringReal;
    imported DataMapOfStringString;
    imported DataMapIteratorOfDataMapOfStringString;
    imported DataMapOfStringByte;
    imported DataMapIteratorOfDataMapOfStringByte;
    imported DataMapOfStringHArray1OfInteger;
    imported DataMapIteratorOfDataMapOfStringHArray1OfInteger;
    imported DataMapOfStringHArray1OfReal;
    imported DataMapIteratorOfDataMapOfStringHArray1OfReal;

    class HDataMapOfStringInteger;   
    
    class HDataMapOfStringReal; 
    
    class HDataMapOfStringString;   
    
    class HDataMapOfStringByte; 
    
    class HDataMapOfStringHArray1OfInteger;  
    
    class HDataMapOfStringHArray1OfReal;  
     
    
    IDList (anIDList : in out IDList from TDF);
	---Purpose: Appends to <anIDList> the list of the attributes
	--          IDs of this package. CAUTION: <anIDList> is NOT
	--          cleared before use.



    Print (DIM : RealEnum from TDataStd; S : in out OStream) 
    	---Purpose: Prints the name of the real dimension <DIM> as a String on
    	--          the Stream <S> and returns <S>.
    	---C++: return &		
    returns OStream;   

end TDataStd;



