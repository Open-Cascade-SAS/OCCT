-- Created on: 1992-02-19
-- Created by: Jean Pierre TIRAULT
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

generic class HDoubleList from PCollection (Item as Storable) 
inherits PManaged 


raises NoSuchObject from Standard

is

	---Purpose: Definition of a double linked list
        -- Idem to the SingleList with a pointer to the previous node

	
	Create returns  mutable HDoubleList;
	---Purpose: Creation of an empty list

	IsEmpty(me) returns Boolean;
        ---Level: Public
	---Purpose: Returns True if the list contains no element.

	Construct(me : mutable; T : Item) returns mutable HDoubleList;
        ---Level: Public
	---Purpose: Adds T at the begining of me.
	---Example: before
	--   me = (A B C) 
        -- after
	--   me = (A B C)
	-- returns 
	--   (T A B C)

	Value(me) returns any Item
                raises NoSuchObject;
        ---Level: Public
	---Purpose: Value of the first node of me
	-- Raises an exception if me is empty
	---Purpose: before
	--   me = (A B C) 
        -- after
	--   me = (A B C)
	-- returns 
	--   A

	Tail(me) returns any HDoubleList
                raises NoSuchObject;
        ---Level: Public
	---Purpose: Returns the end of the list <me>.
	-- Raises an exception if me is empty.
	---Example: before
	--   me = (A B C) 
        -- after
	--   me = (A B C)
	-- returns 
	--   (B C)

	Previous(me) returns any HDoubleList
                raises NoSuchObject;
                ---Level: Public
		---Purpose: Previous node of me.
		-- Raises an exception if me is empty.
		---Example: before
                --   A list L = (A B C) with me = (B C) a sub-list of L.
                -- after
		--   L = (A B C), me = (B C)
		-- returns 
		--   (A)

	SwapTail(me : mutable; WithList : in out any HDoubleList) 
                raises NoSuchObject;
                ---Level: Public
		---Purpose: Exchanges end of me with WithList.
		-- Raises an exception if me is empty.
		---Example: before
		--   me = (A B C)
		--   WithList = (D E)
		-- after
		--   me = (A D E)
		--   WithList = (B C)

	SetValue(me : mutable; T : Item) 
                raises NoSuchObject;
                ---Level: Public
		---Purpose: Changes the value of the first node of me.
		-- Raises an exception if me is empty.
		---Example: before
		--   me = (A B C) 
                -- after
		--   me = (T B C)


	ChangeBackPointer(me : mutable; BackPointer : HDoubleList);
                ---Level: Public
		---Purpose: Modification of the backward pointer

	ChangeForwardPointer(me : mutable; ForwardPointer : 
						HDoubleList);
                ---Level: Public
		---Purpose: Modification of the forward pointer

    	ShallowCopy(me) 
                returns mutable like me 
                is redefined;
                ---Level: Advanced
	    	---C++: function call

    	ShallowDump (me; s: in out OStream) 
                is redefined;
                ---Level: Advanced
    	    	---C++: function call

    	Destroy(me : mutable);
	---C++: alias ~
       
fields 
           Data : 	Item;
           Next : 	HDoubleList;
           Before : 	HDoubleList;

end HDoubleList;
