-- File:	IGESAppli_ToolLevelToPWBLayerMap.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolLevelToPWBLayerMap  from IGESAppli

    ---Purpose : Tool to work on a LevelToPWBLayerMap. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses LevelToPWBLayerMap from IGESAppli,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolLevelToPWBLayerMap;
    ---Purpose : Returns a ToolLevelToPWBLayerMap, ready to work


    ReadOwnParams (me; ent : mutable LevelToPWBLayerMap;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : LevelToPWBLayerMap;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : LevelToPWBLayerMap;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a LevelToPWBLayerMap <ent>, from
    --           its specific (own) parameters

    DirChecker (me; ent : LevelToPWBLayerMap) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : LevelToPWBLayerMap;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : LevelToPWBLayerMap; entto : mutable LevelToPWBLayerMap;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : LevelToPWBLayerMap;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolLevelToPWBLayerMap;
