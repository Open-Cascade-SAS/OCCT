-- Created on: 1998-01-28
-- Created by: Christian CAILLET
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class SignStatus  from IGESSelect    inherits Signature  from IFSelect

    ---Purpose : Gives D.E. Status under the form i,j,k,l (4 figures)
    --           i for BlankStatus
    --           j for SubordinateStatus
    --           k for UseFlag
    --           l for Hierarchy
    --           
    --           For matching, allowed shortcuts
    --           B(Blanked) or V(Visible) are allowed instead of  i
    --           I(Independant=0), P(Physically Dep.=1), L(Logically Dep.=2) or
    --             D(Dependant=3) are allowed instead of  j
    --           These letters must be given in their good position
    --           For non-exact matching :
    --           a letter (see above), no comma : only this status is checked
    --           nothing or a star between commas : this status is OK

uses CString, Transient, AsciiString, InterfaceModel

is

    Create returns mutable SignStatus;

    Value   (me; ent : any Transient; model : InterfaceModel) returns CString;
    ---Purpose : Returns the value (see above)

    Matches (me; ent : Transient; model : InterfaceModel;
    	    	 text : AsciiString; exact : Boolean)
	returns Boolean  is redefined;
    ---Purpose : Performs the match rule (see above)

end SignStatus;
