-- Created on: 1993-01-09
-- Created by: CKY / Contract Toubro-Larsen (SIVA)
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Face from IGESSolid  inherits IGESEntity

        ---Purpose: defines Face, Type <510> Form Number <1>
        --          in package IGESSolid
        --          Face entity is a bound (partial) which has finite area

uses

        Loop              from IGESSolid,
        HArray1OfLoop from IGESSolid

raises OutOfRange

is

        Create returns Face;

            -- Specific Methods pertaining to the class

        Init (me            : mutable;
              aSurface      : IGESEntity;
              outerLoopFlag : Boolean;
              loops         : HArray1OfLoop);
        ---Purpose : This method is used to set the fields of the class Face
        --       - aSurface      : Pointer to the underlying surface
        --       - outerLoopFlag : True means the first loop is the outer loop
        --       - loops         : Array of loops bounding the face

        Surface (me) returns IGESEntity;
        ---Purpose : returns the underlying surface of the face

        NbLoops (me) returns Integer;
        ---Purpose : returns the number of the loops bounding the face

        HasOuterLoop (me) returns Boolean;
        ---Purpose : checks whether there is an outer loop or not

        Loop (me; Index : Integer) returns Loop
        raises OutOfRange;
        ---Purpose : returns the Index'th loop that bounds the face
        -- raises exception if Index < 0 or Index >= NbLoops

fields

--
-- Class    : IGESSolid_Face
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class Face.
--
-- Reminder : A Face instance is defined by :
--            a underlying surface (Surface) bounded by loops (Loops)

        theSurface   : IGESEntity;
            --  underlying surface

        hasOuterLoop : Boolean;
            -- indicator for presence of the outer loop

        theLoops     : HArray1OfLoop;
            -- array of the bounding loops

end Face;
