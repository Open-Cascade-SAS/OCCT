-- Created on: 1997-02-12
-- Created by: Alexander BRIVIN
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class OrthographicCamera from Vrml 

	---Purpose: specifies a OrthographicCamera node of VRML specifying properties of cameras. 
    	--  An orthographic camera defines a parallel projection from a viewpoint. This camera does
       	--  not diminish objects with distance, as a PerspectiveCamera does. The viewing volume for
       	--  an orthographic camera is a rectangular parallelepiped (a box). 
uses
 
    Vec         from gp, 
    SFRotation  from Vrml

is 
                                                    --  defaults  :
    Create  returns  OrthographicCamera from Vrml;  --  myPosition(0 0 1)
 						    --  myOrientation(0 0 1 0)
						    --  myFocalDistance(5)
						    --  myHeight(2)
    	    	    	    	    	    	    --  Camera looks along the negative Z-axis
    Create  ( aPosition      :  Vec         from  gp;   
    	      aOrientation   :  SFRotation  from  Vrml; 
    	      aFocalDistance :  Real        from  Standard; 
    	      aHeight        :  Real        from  Standard )
    	returns  OrthographicCamera from Vrml; 
	 
    SetPosition ( me : in out;  aPosition : Vec  from  gp );
    Position ( me )  returns Vec  from  gp;

    SetOrientation ( me : in out;  aOrientation : SFRotation  from  Vrml );
    Orientation ( me )  returns SFRotation  from  Vrml;

    SetFocalDistance ( me : in out;  aFocalDistance : Real  from  Standard );
    FocalDistance ( me )  returns Real  from  Standard;

    SetHeight ( me : in out;  aHeight : Real  from  Standard );
    Height ( me )  returns Real  from  Standard;

    Print  ( me;  anOStream: in out OStream from Standard) returns OStream from Standard;
    ---C++:  return  & 
    
fields
 
    myPosition      :  Vec         from  gp;        -- Location of viewpoint
    myOrientation   :  SFRotation  from  Vrml;      -- Orientation (rotation with respect to (0,0,-1) vector)
    myFocalDistance :  Real        from  Standard;  -- Distance from viewpoint to point of focus.
    myHeight        :  Real        from  Standard;  -- Height of view volume

end OrthographicCamera;

