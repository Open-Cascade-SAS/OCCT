-- Created on: 1998-06-30
-- Created by: Christian CAILLET
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ProductDefinitionWithAssociatedDocuments  from StepBasic
    inherits ProductDefinition  from StepBasic

uses
     HAsciiString from TCollection,
     ProductDefinitionFormation from StepBasic,
     ProductDefinitionContext from StepBasic,
     Document from StepBasic,
     HArray1OfDocument from StepBasic

is

    Create returns ProductDefinitionWithAssociatedDocuments;

    Init (me : mutable;
    	  aId : HAsciiString;
    	  aDescription : HAsciiString;
    	  aFormation : ProductDefinitionFormation;
	  aFrame : ProductDefinitionContext;
	  aDocIds : HArray1OfDocument);

    DocIds (me) returns HArray1OfDocument;
    SetDocIds (me : mutable; DocIds : HArray1OfDocument);
    NbDocIds (me) returns Integer;
    DocIdsValue (me; num : Integer) returns Document;
    SetDocIdsValue (me : mutable; num : Integer; adoc : Document);

fields

    theDocIds : HArray1OfDocument;

end ProductDefinitionWithAssociatedDocuments;
