-- Created on: 1997-05-28
-- Created by: Xavier BENVENISTE
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class CheckBSplineCurve from GeomLib

	---Purpose: this class is used to  construct the BSpline curve
	--          from an Approximation ( ApproxAFunction from AdvApprox).
    	

uses
    Pnt	            from gp,
    BSplineCurve    from Geom,
    BSplineCurve    from Geom2d

raises

    NotDone    from StdFail,
    OutOfRange from Standard
    
is

    Create( Curve : BSplineCurve from Geom ;
    	    Tolerance        : Real from Standard ;
            AngularTolerance : Real from Standard) 
    returns CheckBSplineCurve from GeomLib;
    
    IsDone(me) returns Boolean from Standard
	---C++: inline
    is static;
    
    NeedTangentFix(me; FirstFlag : in out Boolean from Standard ;
    	         SecondFlag : in out Boolean from Standard) ;
    FixTangent  (me : in out ; FirstFlag : Boolean from Standard ;
              		       LastFlag  : Boolean from Standard)  ;	 
	
    FixedTangent  (me : in out ; FirstFlag : Boolean from Standard ;
              		       LastFlag  : Boolean from Standard) 
    ---Purpose:  modifies the curve
    -- by fixing the first or the last tangencies 
    -- 
    returns BSplineCurve from Geom
    raises
    	OutOfRange from Standard,
    	---Purpose: if Index3D not in the Range [1,Nb3dSpaces]
	NotDone    from StdFail
	---Purpose: if the Approx is not Done
    is static;
 

fields

    myCurve            : BSplineCurve from Geom ;
    myDone             : Boolean from Standard ;
    myFixFirstTangent  : Boolean from Standard ;
    myFixLastTangent   : Boolean from Standard ;
    myAngularTolerance : Real from Standard ;
    myTolerance        : Real from Standard ;
    myFirstPole        : Pnt from gp ;
    	-- the second pole that controls first tangency
    myLastPole         : Pnt from gp ;
    	-- the before last pole that controls last tangency

end CheckBSplineCurve;
