-- Created on: 1993-01-21
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Iterator from TopoDS 

	---Purpose: Iterates on the underlying shape underlying a given
	-- TopoDS_Shape object, providing access to its
	-- component sub-shapes. Each component shape is
	-- returned as a TopoDS_Shape with an orientation,
	-- and a compound of the original values and the relative values.

uses
    Shape                     from TopoDS,
    ListIteratorOfListOfShape from TopoDS,
    Location                  from TopLoc,
    Orientation               from TopAbs

raises
    NoMoreObject from Standard,
    NoSuchObject from Standard

is
    Create returns Iterator from TopoDS;
    ---C++: inline
	---Purpose: Creates an empty Iterator.


    Create(S : Shape from TopoDS;
    	   cumOri : Boolean = Standard_True;
    	   cumLoc : Boolean = Standard_True) returns Iterator from TopoDS;
    ---C++: inline
	---Purpose: Creates an Iterator on <S> sub-shapes.
	--      Note:
	-- - If cumOri is true, the function composes all
	--   sub-shapes with the orientation of S.
	-- - If cumLoc is true, the function multiplies all
	--   sub-shapes by the location of S, i.e. it applies to
	--   each sub-shape the transformation that is associated with S.

    Initialize(me : in out; S      : Shape from TopoDS;
    	                    cumOri : Boolean = Standard_True;
    	                    cumLoc : Boolean = Standard_True)
	---Purpose: Initializes this iterator with shape S.
	-- Note:
	-- - If cumOri is true, the function composes all
	--   sub-shapes with the orientation of S.
	-- - If cumLoc is true, the function multiplies all
	--   sub-shapes by the location of S, i.e. it applies to
	--   each sub-shape the transformation that is associated with S.
    is static;
    
    More(me) returns Boolean
	---Purpose: Returns true if there is another sub-shape in the
	-- shape which this iterator is scanning.
    ---C++: inline
    is static;
    
    Next(me : in out)
	---Purpose: Moves on to the next sub-shape in the shape which
	-- this iterator is scanning.
	-- Exceptions
	-- Standard_NoMoreObject if there are no more sub-shapes in the shape.
    raises
    	NoMoreObject from Standard
    is static;
    
    Value(me) returns Shape from TopoDS
	---Purpose: Returns the current sub-shape in the shape which
	-- this iterator is scanning.
	-- Exceptions
	-- Standard_NoSuchObject if there is no current sub-shape.
    raises
    	NoSuchObject from Standard
	---C++: return const &
    ---C++: inline
    is static;

    
fields
    myShape       : Shape                     from TopoDS;
    myShapes      : ListIteratorOfListOfShape from TopoDS;
    myOrientation : Orientation               from TopAbs;
    myLocation    : Location                  from TopLoc;

end Iterator;
