-- Created on: 1999-03-11
-- Created by: data exchange team
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class RevolvedFaceSolid from StepShape 
inherits SweptFaceSolid from StepShape 
	

uses
    	Axis1Placement from StepGeom, 
	Real from Standard, 
	HAsciiString from TCollection,
	FaceSurface from StepShape 

is
    	Create returns mutable RevolvedFaceSolid;
	---Purpose: Returns a RevolvedFaceSolid


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aSweptArea : mutable FaceSurface from StepShape) is redefined ;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aSweptArea : mutable FaceSurface from StepShape;
	      aAxis : mutable Axis1Placement from StepGeom;
	      aAngle : Real from Standard);

	-- Specific Methods for Field Data Access --

	SetAxis(me : mutable; aAxis : mutable Axis1Placement);
	Axis (me) returns mutable Axis1Placement;
	SetAngle(me : mutable; aAngle : Real);
	Angle (me) returns Real;


fields

    	axis : Axis1Placement from StepGeom;
	angle : Real from Standard;

end RevolvedFaceSolid;
