-- File:	BinMDataStd_NamedDataDriver.cdl
-- Created:	Mon Jul  2 10:16:56 2007
-- Author:	Sergey ZARITCHNY
--		<sergey.zaritchny@opencascade.com>
---Copyright:	Open CasCade SA 2007


class NamedDataDriver from BinMDataStd inherits ADriver from BinMDF

	---Purpose: 

uses
    MessageDriver    from CDM,
    SRelocationTable from BinObjMgt,
    RRelocationTable from BinObjMgt,
    Persistent       from BinObjMgt,
    Attribute        from TDF

is
    Create (theMessageDriver:MessageDriver from CDM)
    returns mutable NamedDataDriver from BinMDataStd;

    NewEmpty (me)
    returns mutable Attribute from TDF
    is redefined;

    Paste(me; Source     : Persistent from BinObjMgt;
              Target     : mutable Attribute from TDF;
              RelocTable : out RRelocationTable from BinObjMgt)
    returns Boolean from Standard is redefined;

    Paste(me; Source     : Attribute from TDF;
              Target     : in out Persistent from BinObjMgt;
              RelocTable : out SRelocationTable from BinObjMgt)
    is redefined;

end NamedDataDriver;
