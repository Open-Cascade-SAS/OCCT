-- Created on: 2003-06-04
-- Created by: Galina KULIKOVA
-- Copyright (c) 2003-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



package RWStepDimTol 

	---Purpose: Packsge contains tools for parsing and formatting GD&T entities.

    uses
    	TCollection,
    	RWStepRepr, 
    	RWStepShape,
    	RWStepVisual,
    	RWStepBasic,
    	TColStd,
	StepData,
    	Interface, 
	StepDimTol,
    	MMgt

    is
    	class RWAngularityTolerance;
    	class RWCircularRunoutTolerance;
    	class RWConcentricityTolerance;
    	class RWCylindricityTolerance;
    	class RWCoaxialityTolerance;
    	class RWFlatnessTolerance;
    	class RWLineProfileTolerance;
    	class RWParallelismTolerance;
    	class RWPerpendicularityTolerance;
    	class RWPositionTolerance;
    	class RWRoundnessTolerance;
    	class RWStraightnessTolerance;
    	class RWSurfaceProfileTolerance;
    	class RWSymmetryTolerance;
    	class RWTotalRunoutTolerance;
    
    	class RWGeometricTolerance;
    	class RWGeometricToleranceRelationship;
    	class RWGeometricToleranceWithDatumReference;
    	class RWModifiedGeometricTolerance;
     
    	class RWDatum;
    	class RWDatumFeature;
    	class RWDatumReference;
    	class RWCommonDatum;
    	class RWDatumTarget;
    	class RWPlacedDatumTargetFeature;
    	
	class RWGeoTolAndGeoTolWthDatRefAndModGeoTolAndPosTol;


end RWStepDimTol;
