-- Created on: 1999-11-29
-- Created by: Peter KURNEV
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class VertexInfo from TopOpeBRepBuild 

	---Purpose: 

uses
    Vertex  from  TopoDS,  
    Edge    from  TopoDS,
    SequenceOfInteger  from  TColStd, 
    IndexedMapOfOrientedShape from TopTools,
    ListOfShape  from TopTools
--raises

is
    Create     returns VertexInfo from TopOpeBRepBuild; 
     
    SetVertex    (me:out;  aV:Vertex  from  TopoDS); 
     
    Vertex       (me)  returns  Vertex  from  TopoDS;  
    ---C++: return const & 
     
    SetSmart     (me:out;  aFlag: Boolean  from  Standard);
     
    Smart        (me)  returns Boolean  from  Standard; 
     
    NbCases    (me) returns  Integer  from  Standard; 
     
    FoundOut   (me) returns  Integer  from  Standard; 
     
    AddIn        (me:out;  anE:  Edge  from  TopoDS);	      
     
    AddOut       (me:out;  anE:  Edge  from  TopoDS);	      

    SetCurrentIn (me:out;  anE:  Edge  from  TopoDS);	 
     
    EdgesIn    (me) returns IndexedMapOfOrientedShape from TopTools;    
    ---C++: return const & 
     
    EdgesOut   (me) returns IndexedMapOfOrientedShape from TopTools;      
    ---C++: return const & 

    ChangeEdgesOut   (me:out) returns IndexedMapOfOrientedShape from TopTools;      
    ---C++: return &  
    
    Dump       (me); 
   
    CurrentOut (me:out)  returns  Edge from  TopoDS; 
    ---C++: return const &  
     
    AppendPassed  (me:out; anE:  Edge  from  TopoDS); 
     
    RemovePassed  (me:out);  
     
    ListPassed    (me)  returns  ListOfShape  from TopTools;
    ---C++: return const &  
     
    Prepare(me:  out;  aL  :   ListOfShape  from TopTools);
    
fields
    myVertex         :  Vertex  from  TopoDS; 
    myCurrent        :  Edge  from  TopoDS;  
    myCurrentIn      :  Edge  from  TopoDS;  

    mySmart          :  Boolean  from  Standard; 
    
    myEdgesIn        :  IndexedMapOfOrientedShape from TopTools; 
    myEdgesOut       :  IndexedMapOfOrientedShape from TopTools;  
    myLocalEdgesOut  :  IndexedMapOfOrientedShape from TopTools; 
    myEdgesPassed    :  ListOfShape  from TopTools; 
    
    myFoundOut  :  Integer from Standard;    
    
end VertexInfo;








