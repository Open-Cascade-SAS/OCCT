-- Created on: 1998-01-22
-- Created by: Sergey ZARITCHNY
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MinRadiusDimension from AIS inherits EllipseRadiusDimension from AIS

	---Purpose:--  Ellipse  Min  radius  dimension  of  a  Shape  which   
    	--  can  be  Edge  or  Face  (planar  or  cylindrical(surface  of   
    	--  extrusion  or  surface  of  offset)) 	 

uses
 
     Shape                 from TopoDS,
     Elips                 from gp,
     Pnt                   from gp, 
     Pln                   from gp,  
     Ellipse               from Geom, 
     Plane                 from Geom, 
     Surface               from Geom,
     Presentation          from Prs3d,
     PresentationManager3d from PrsMgr,
     Selection             from SelectMgr,
     Projector             from Prs3d,
     Transformation        from Geom,
     ExtendedString        from TCollection,    
     ArrowSide             from DsgPrs, 
     KindOfSurface         from AIS,
     KindOfDimension       from AIS 


raises ConstructionError from Standard

is
 
     
    Create (aShape      : Shape          from TopoDS;
	    aVal        : Real           from Standard;
	    aText       : ExtendedString from TCollection)    
	    ---Purpose: Max  Ellipse  radius dimension 
	    --  Shape  can  be  edge  ,  planar  face  or  cylindrical  face 
    	    --  
    returns mutable MinRadiusDimension from AIS;

    Create (aShape      : Shape          from TopoDS;
	    aVal        : Real           from Standard;
	    aText       : ExtendedString from TCollection;	    
	    aPosition   : Pnt            from gp;
	    aSymbolPrs  : ArrowSide      from DsgPrs;    
    	    anArrowSize : Real           from Standard = 0.0)
	    ---Purpose:  Max  Ellipse  radius dimension with  position
	    --  Shape  can  be  edge  ,  planar  face  or  cylindrical  face 
    	    --   
    returns mutable MinRadiusDimension  from AIS;



              
-- Methods from PresentableObject

    Compute(me                  : mutable;
    	    aPresentationManager: PresentationManager3d from PrsMgr;
    	    aPresentation       : mutable Presentation from Prs3d;
    	    aMode               : Integer from Standard= 0) 
    is redefined private;
    
    Compute(me:mutable;
    	        aProjector: Projector from Prs3d;
                aPresentation: mutable Presentation from Prs3d)
    is redefined static private;     
    
    Compute(me            : mutable;
    	    aProjector    : Projector from Prs3d;
    	    aTrsf         : Transformation from Geom;
	    aPresentation : mutable Presentation from Prs3d)
    is redefined;
    ---Purpose: computes the presentation according to a point of view
    --          given by <aProjector>. 
    --          To be Used when the associated degenerated Presentations 
    --          have been transformed by <aTrsf> which is not a Pure
    --          Translation. The HLR Prs can't be deducted automatically
    --          WARNING :<aTrsf> must be applied
    --           to the object to display before computation  !!!

-- Methods from SelectableObject

    ComputeSelection(me         : mutable;
    	    	     aSelection : mutable Selection from SelectMgr;
    	    	     aMode      : Integer from Standard)
    is redefined private;

--
--     Computation private methods
--

    ComputeEllipse(me: mutable;
    	    	     	aPresentation : mutable Presentation from Prs3d)
    is private; 
     
    ComputeArcOfEllipse(me: mutable;
    	    	     	aPresentation : mutable Presentation from Prs3d  )
    is private; 

fields 

    myApexP       :  Pnt  from  gp;  
    myApexN       :  Pnt  from  gp; 
    myEndOfArrow  :  Pnt  from  gp; 
    
end MinRadiusDimension;
