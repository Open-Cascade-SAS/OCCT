-- Created on: 1999-09-08
-- Created by: Andrey BETENEV
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MeasureRepresentationItem from StepRepr 
    inherits RepresentationItem from StepRepr 

	---Purpose: Implements a measure_representation_item entity
	--          which is used for storing validation properties
	--          (e.g. area) for shapes

uses
    HAsciiString       from TCollection,
    Unit               from StepBasic,
    MeasureWithUnit    from StepBasic,
    MeasureValueMember from StepBasic
    
is
    Create returns mutable MeasureRepresentationItem;
        ---Purpose: Creates empty object
    
    Init (me : mutable;
	  aName : mutable HAsciiString from TCollection;
	  aValueComponent : MeasureValueMember from StepBasic;
	  aUnitComponent : Unit from StepBasic);
        ---Purpose: Init all fields

    SetMeasure (me: mutable; Measure: MeasureWithUnit from StepBasic);
    Measure (me) returns MeasureWithUnit from StepBasic;
    
fields
    myMeasure: MeasureWithUnit from StepBasic;

end MeasureRepresentationItem;

