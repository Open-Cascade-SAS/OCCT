-- Created on: 1994-09-05
-- Created by: Gilles DEBARBOUILLE
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class CompositVariableInstance from Dynamic

inherits

    AbstractVariableInstance from Dynamic
	---Purpose: This  class corresponds to  the instanciation of a
	--          variable group. It allows the setting of more than
	--          one variable in  a variable instance. It is useful
	--          when a  method takes  a collection  of homogeneous
	--          objects as   argument. For   example a wire  needs
	--          edges as argument.
   
uses

    Variable     from Dynamic,
    VariableNode from Dynamic


is

    Create returns mutable CompositVariableInstance from Dynamic;
    
    ---Level: Advanced 
    
    ---Purpose: Creates  a new  empty  instance of   CompositVariable-
    --          Instance.
    
    Variable(me : mutable ; avariable : Variable from Dynamic)
    
    ---Purpose: Sets <avariable> into the collection of variable.
    
    is redefined;
    
    FirstVariableNode(me) returns VariableNode from Dynamic
    
    ---Purpose: Returns the first VariableNode  useful to explore  the
    --          list of variables addressed by <me>.
    
    is static;

fields

    thefirstvariablenode : VariableNode from Dynamic;

end CompositVariableInstance;
