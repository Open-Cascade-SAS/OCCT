-- Created on: 2002-12-12
-- Created by: data exchange team
-- Copyright (c) 2002-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


package RWStepFEA

uses

	StepData, Interface, TCollection, TColStd, StepFEA

is

    class RWAlignedCurve3dElementCoordinateSystem;
    class RWArbitraryVolume3dElementCoordinateSystem;
    class RWCurve3dElementProperty;
    class RWCurve3dElementRepresentation;
    class RWCurveElementEndOffset;
    class RWCurveElementEndRelease;
    class RWCurveElementInterval;
    class RWCurveElementIntervalConstant;
    class RWCurveElementLocation;
    class RWDummyNode;
    class RWElementGeometricRelationship;
    class RWElementGroup;
    class RWElementRepresentation;
    class RWFeaAreaDensity;
    class RWFeaAxis2Placement3d;
    class RWFeaGroup;
    class RWFeaLinearElasticity;
    class RWFeaMassDensity;
    class RWFeaMaterialPropertyRepresentation;
    class RWFeaMaterialPropertyRepresentationItem;
    class RWFeaModel;
    class RWFeaModel3d;
    class RWFeaMoistureAbsorption;
    class RWFeaParametricPoint;
    class RWFeaRepresentationItem;
    class RWFeaSecantCoefficientOfLinearThermalExpansion;
    class RWFeaShellBendingStiffness;
    class RWFeaShellMembraneBendingCouplingStiffness;
    class RWFeaShellMembraneStiffness;
    class RWFeaShellShearStiffness;
    class RWFeaTangentialCoefficientOfLinearThermalExpansion;
    class RWGeometricNode;
    class RWNode;
    class RWNodeGroup;
    class RWNodeRepresentation;
    class RWNodeSet;
    class RWNodeWithSolutionCoordinateSystem;
    class RWNodeWithVector;
    class RWParametricCurve3dElementCoordinateDirection;
    class RWParametricCurve3dElementCoordinateSystem;
    class RWParametricSurface3dElementCoordinateSystem;
    class RWSurface3dElementRepresentation;
    class RWVolume3dElementRepresentation;
    class RWFeaModelDefinition;
    class RWFreedomAndCoefficient;
    class RWFreedomsList;
    class RWNodeDefinition;
    class RWAlignedSurface3dElementCoordinateSystem;
    class RWConstantSurface3dElementCoordinateSystem;
    class RWCurveElementIntervalLinearlyVarying;    -- added 23.01.2003
    class RWFeaCurveSectionGeometricRelationship;   -- added 23.01.2003
    class RWFeaSurfaceSectionGeometricRelationship; -- added 23.01.2003

end;
