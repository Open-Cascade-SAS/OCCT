-- Created on: 1994-04-18
-- Created by: Modelistation
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Circle2D from Draw inherits Drawable2D from Draw

	---Purpose: 

uses
    Circ2d from gp,
    Color from Draw,
    Display from Draw

is

    Create(C : Circ2d from gp; A1,A2 : Real; col : Color)
    returns Circle2D;
    
    DrawOn(me; dis : in out Display);

fields

    myCirc  : Circ2d from gp;
    myA1    : Real;
    myA2    : Real;
    myColor : Color;
    
end Circle2D;

