-- Created on: 1997-08-22
-- Created by: VAUTHIER Jean-Claude
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Sphere from QANewBRepNaming inherits TopNaming from QANewBRepNaming

    ---Purpose: To load the Sphere results 

uses 
 
    MakeSphere from BRepPrimAPI,
    Label      from TDF,
    TypeOfPrimitive3D from QANewBRepNaming

is
     
    Create returns Sphere from QANewBRepNaming;
      
    Create(ResultLabel : Label from TDF) 
    returns Sphere from QANewBRepNaming;
      
    Init(me : in out; ResultLabel : Label from TDF);
     
    
    Load (me; mkSphere : in out MakeSphere from BRepPrimAPI; Type : TypeOfPrimitive3D from QANewBRepNaming);

    Bottom (me)
    ---Purpose: Returns the label of the bottom
    --          face of the Sphere.
    returns Label from TDF;

    Top (me)
    ---Purpose: Returns the label of the top
    --          face of the Sphere.
    returns Label from TDF;

    Lateral (me)
    ---Purpose: Returns the label of the lateral
    --          face of the Sphere.
    returns Label from TDF;

    StartSide (me)
    ---Purpose: Returns the label of the first
    --          side of the Sphere.
    returns Label from TDF;
        
    EndSide (me)
    ---Purpose: Returns the label of the second
    --          side of the Sphere.
    returns Label from TDF;

    Meridian (me)
    ---Purpose: Returns the label of the meridian
    --          edges of the Sphere.
    returns Label from TDF;

    Degenerated (me)
    ---Purpose: Returns the label of the degenerated
    --          edges of the Sphere.
    returns Label from TDF;

end Sphere;
