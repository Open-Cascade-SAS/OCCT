-- File:	GeomTools_SurfaceSet.cdl
-- Created:	Mon Jul 19 15:21:50 1993
-- Author:	Remi LEQUETTE
--		<rle@nonox>
---Copyright:	 Matra Datavision 1993



class SurfaceSet from GeomTools 

	---Purpose: Stores a set of Surfaces from Geom.

uses
    Surface               from Geom,
    IndexedMapOfTransient from TColStd,
    ProgressIndicator     from Message
    
raises
    OutOfRange from Standard

is

    Create returns SurfaceSet from GeomTools;
	---Purpose: Returns an empty set of Surfaces.
	
    Clear(me : in out)
	---Purpose: Clears the content of the set.
    is static;
	
    Add(me : in out; S : Surface from Geom) returns Integer
	---Purpose: Incorporate a new Surface in the  set and returns
	--          its index.
    is static;
    
    Surface(me; I : Integer) returns Surface from Geom
	---Purpose: Returns the Surface of index <I>.
    raises
    	OutOfRange from Standard
    is static;

    Index(me; S : Surface from Geom) returns Integer
	---Purpose: Returns the index of <L>.
    is static;
    
    Dump(me; OS : in out OStream)
	---Purpose: Dumps the content of me on the stream <OS>.
    is static;
	
    Write(me; OS : in out OStream)
	---Purpose: Writes the content of  me  on the stream <OS> in a
	--          format that can be read back by Read.
    is static;
	
    Read(me : in out; IS : in out IStream)
	---Purpose: Reads the content of me from the  stream  <IS>. me
	--          is first cleared.
	--          
    is static;
	
    --
    -- 	class methods to write an read surfaces
    -- 	
    
    PrintSurface(myclass; S  : Surface from Geom;
    	    	    	  OS : in out OStream;
			  compact : Boolean = Standard_False);
	---Purpose: Dumps the surface on the stream,  if compact is True
	--          use the compact format that can be read back.
	
    ReadSurface(myclass; IS : in out IStream;
    	    	         S  : in out Surface from Geom)
    returns IStream;
	---Purpose: Reads the surface  from  the stream.  The  surface  is
	--          assumed   to have  been  writtent  with  the Print
	--          method (compact = True).
	--          
	---C++: return &
	
    SetProgress(me : in out; PR : ProgressIndicator from Message);

    GetProgress(me) returns ProgressIndicator from Message;

fields

    myMap : IndexedMapOfTransient from TColStd;
    myProgress : ProgressIndicator from Message;

end SurfaceSet;


