-- File:        GeneralModule.cdl
-- Created:     Thu Dec  7 14:30:07 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class GeneralModule from RWStepAP214  inherits GeneralModule from StepData
	---Purpose : Defines General Services for StepAP214 Entities
	--           (Share,Check,Copy; Trace already inherited)
	--           Depends (for case numbers) of Protocol from StepAP214

uses Transient,  HAsciiString from TCollection,
     EntityIterator from Interface,
     ShareTool      from Interface,
     Check          from Interface,
     CopyTool       from Interface,
     InterfaceModel from Interface

is

    Create returns mutable GeneralModule from RWStepAP214;
    ---Purpose : Creates a GeneralModule

    FillSharedCase (me; CN : Integer; ent : Transient;
                        iter : in out EntityIterator);
    ---Purpose : Specific filling of the list of Entities shared by an Entity
    --           <ent>, according to a Case Number <CN> (provided by StepAP214
    --           Protocol).

    CheckCase (me; CN : Integer; ent : Transient; shares : ShareTool; ach : in out Check);
    ---Purpose : Specific Checking of an Entity <ent>

    CopyCase (me; CN : Integer; entfrom : Transient; entto : mutable Transient; TC : in out CopyTool);
    ---Purpose : Specific Copy ("Deep") from <entfrom> to <entto> (same type)
    --           by using a CopyTool which provides its working Map.
    --           Use method Transferred from CopyTool to work


    NewVoid (me; CN : Integer; ent : out mutable Transient) returns Boolean;

    CategoryNumber (me; CN : Integer; ent : Transient; shares : ShareTool)
    returns Integer  is redefined;

    Name (me; CN : Integer; ent : Transient; shares : ShareTool from Interface)
    returns HAsciiString from TCollection  is redefined;
    ---Purpose : Returns the name of a STEP Entity according to its type

end GeneralModule;
