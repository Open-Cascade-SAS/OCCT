-- Created on: 1993-01-09
-- Created by: CKY / Contract Toubro-Larsen ( Anand NATRAJAN )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ExternalRefFileName from IGESBasic  inherits IGESEntity

        ---Purpose: defines ExternalRefFileName, Type <416> Form <0-2>
        --          in package IGESBasic
        --          Used when single definition from the reference file is
        --          required or for external logical references where an
        --          entity in one file relates to an entity in another file

uses

        HAsciiString from TCollection

is

        Create returns mutable ExternalRefFileName;

        -- Specific Methods pertaining to the class

        Init (me : mutable; aFileIdent, anExtName : HAsciiString);
        ---Purpose : This method is used to set the fields of the class
        --           ExternalRefFileName
        --       - aFileIdent : External Reference File Identifier
        --       - anExtName  : External Reference Entity Symbolic Name

    	SetForEntity (me : mutable; mode : Boolean);
	---Purpose : Changes FormNumber to be 2 if <mode> is True (For Entity)
	--           or 0 if <mode> is False (For Definition)

        FileId (me) returns HAsciiString from TCollection;
        ---Purpose : returns External Reference File Identifier

        ReferenceName (me) returns HAsciiString from TCollection;
        ---Purpose : returns External Reference Entity Symbolic Name

fields

--
-- Class    : IGESBasic_ExternalRefFileName
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class ExternalRefFileName.
--
-- Reminder : A ExternalRefFileName instance is defined by :
--            - External Reference File Identifier
--            - External Reference Entity Symbolic Name

        theExtRefFileIdentifier : HAsciiString from TCollection;
        theExtRefEntitySymbName : HAsciiString from TCollection;

end ExternalRefFileName;
