-- Created on: 1993-06-08
-- Created by: Laurent BOURESCHE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Tool from BRepSweep -- as Tool from Sweep

    ---Purpose: Provides  the  indexation and type  analysis  services
    --          required by the TopoDS generating Shape of BRepSweep.
    --          

uses

    Shape from TopoDS,
    IndexedMapOfShape from TopTools,
    ShapeEnum from TopAbs,
    Orientation from TopAbs

raises 

    OutOfRange from Standard

is

    Create(aShape: Shape from TopoDS);
	---Purpose: Initialize the tool  with <aShape>.  The IndexTool
	--          must prepare an indexation for  all  the subshapes
	--          of this shape.

    NbShapes(me) returns Integer
	---Purpose: Returns the number of subshapes in the shape.
    is static;

    Index(me; aShape : Shape from TopoDS) returns Integer
	---Purpose: Returns the index of <aShape>.
    is static;
    
    Shape(me; anIndex : Integer from Standard) returns Shape from TopoDS
	---Purpose: Returns the Shape at Index anIdex.
    is static;
    
    Type(me; aShape : Shape from TopoDS) returns ShapeEnum from TopAbs
	---Purpose: Returns the type of <aShape>.
    is static;

    Orientation (me; aShape : Shape from TopoDS) 
    returns Orientation from TopAbs
	---Purpose: Returns the Orientation of <aShape>.
    is static;

    SetOrientation (me; 
    	    	    aShape : in out Shape from TopoDS; 
    	    	    Or     : Orientation  from  TopAbs) 
	---Purpose: Set the Orientation of <aShape> with Or.
    is static;

fields

    myMap : IndexedMapOfShape from TopTools;
    
end Tool from BRepSweep;



