-- Created on: 1993-01-11
-- Created by: CKY / Contract Toubro-Larsen ( SIVA )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class OrdinateDimension from IGESDimen  inherits IGESEntity

        ---Purpose: defines IGES Ordinate Dimension, Type <218> Form <0, 1>,
        --          in package IGESDimen
        -- Note   : The ordinate dimension entity is used to
        --          indicate dimensions from a common base line.
        --          Dimensioning is only permitted along the XT
        --          or YT axis.

uses

        LeaderArrow from IGESDimen,
        WitnessLine from IGESDimen,
        GeneralNote from IGESDimen

is

        Create returns OrdinateDimension;

            -- --specific-- --

        Init(me       : mutable;
             aNote    : GeneralNote;
             aType    : Boolean;
             aLine    : WitnessLine;
             anArrow  : LeaderArrow);
        -- This method is used to set fields of the
        -- class OrdinateDimension
        --       - aNote    : Note for the dimension
        --       - aType    : Type (Witness line or leader arrow)
        --                    (Ignored if form no. = 1)
        --       - aLine    : Witness line used for the dimension
        --       - anArrow  : Leader arrow used for the dimension

        IsLine(me) returns Boolean;
        ---Purpose : returns True if Witness Line and False if Leader (only for Form 0)

        IsLeader(me) returns Boolean;
        ---Purpose : returns True if Leader and False if Witness Line (only for Form 0)

        Note(me) returns GeneralNote;
        ---Purpose : returns the General Note entity associated.

        WitnessLine(me) returns WitnessLine;
        ---Purpose : returns the Witness Line associated or Null handle

        Leader(me) returns LeaderArrow;
        ---Purpose : returns the Leader associated or Null handle

fields

--
-- Class    : IGESDimen_OrdinateDimension
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class OrdinateDimension.
--
-- Reminder : A OrdinateDimension instance is defined by :
--            - A General Note
--            - A Boolean field determining whether a Witness Line
--                                or Leader is present
--            - A Witness Line
--            - A Leader Arrow
--

        theNote        : GeneralNote;
        isItLine       : Boolean;     --True if Witness Line, False if Leader
        theWitnessLine : WitnessLine;
        theLeader      : LeaderArrow;

end OrdinateDimension;
