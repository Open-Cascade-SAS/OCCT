-- Created on: 1994-01-14
-- Created by: Gilles DEBARBOUILLE
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MaterialDefinition from Materials

inherits

    FuzzyDefinitionsDictionary from Dynamic 
     
    
	---Purpose: This  inherited  class  is  useful  to create  the
	--          abstract description  of  a material,  in  term of
	--          authorized properties.

uses

    Parameter from Dynamic

    
is

    Create returns mutable MaterialDefinition from Materials;
    
    ---Level: Internal 

    ---Purpose: Creates the exhaustive definition of a material.

    Switch(me ; aname , atype , avalue : CString from Standard) returns Parameter from Dynamic
    
    ---Level: Internal 

    ---Purpose: Starting with the identifier of the parameter <aname>,
    --          the type  of parameter <atype>  and a  string <avalue>
    --          which describes  the values  useful  for  this type of
    --          parameters,  creates and returns  a  Parameter  object
    --          from Dynamic.
    
    is redefined;
    
--fields

end MaterialDefinition;
