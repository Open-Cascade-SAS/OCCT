-- File:	QualifiedLin.cdl
-- Created:	Mon Apr 15 15:19:09 1991
-- Author:	Philippe DAUTRY
--		<fid@phobox>
---Copyright:	 Matra Datavision 1991


class QualifiedLin

from GccEnt

inherits Storable from Standard

    	--- Purpose: Describes a qualified 2D line.
    	-- A qualified 2D line is a line (gp_Lin2d line) with a
    	-- qualifier which specifies whether the solution of a
    	-- construction algorithm using the qualified line (as an argument):
    	-- -   is 'enclosed' by the line, or
    	-- -   is built so that both the line and it are external to one another, or
    	-- -   is undefined (all solutions apply).
    	-- Note: the interior of a line is defined as the left-hand
    	-- side of the line in relation to its orientation (i.e. when
    	-- moving from the start to the end of the curve).       
        
        
uses Position from GccEnt, 
     Lin2d    from gp

is

Create(Qualified : Lin2d    from gp        ;
       Qualifier : Position from GccEnt ) 
returns QualifiedLin from GccEnt;
    	---Purpose:
    	-- Constructs a qualified line by assigning the qualifier
    	-- Qualifier to the line Qualified.
    	-- Qualifier may be:
    	-- -   GccEnt_enclosed if the solution is enclosed by the line, or
	-- -   GccEnt_outside if both the solution and the line are external to one another, or
    	-- -   GccEnt_unqualified if all solutions apply.
    	-- Note : the interior of a line is defined as the left-hand
    	-- side of the line in relation to its orientation.

Qualified(me) returns Lin2d from gp
is static;
    	---Purpose: Returns a 2D line to which the qualifier is assigned.
    
Qualifier(me) returns Position from GccEnt
is static;
    	---Purpose:
    	-- Returns the qualifier of this qualified line, if it is "enclosed" or
    	--   "outside", or
    	-- -   GccEnt_noqualifier if it is unqualified.
    
IsUnqualified(me) returns Boolean from Standard
is static;
    	---Purpose: Returns true if the solution is unqualified and false in 
    	--          the other cases.

IsEnclosed(me) returns Boolean from Standard
is static;
    	---Purpose: Returns true if the solution is Enclosed in the Lin2d and false in 
    	--          the other cases.

IsOutside(me) returns Boolean from Standard
is static;
    	---Purpose: Returns true if the solution is Outside the Lin2d and false in 
    	--          the other cases.

fields

TheQualifier : Position from GccEnt;
TheQualified : Lin2d    from gp;

--friends

--Unqualified(Obj : Lin2d) from GccEnt,
--Enclosed   (Obj : Lin2d) from GccEnt,
--Outside    (Obj : Lin2d) from GccEnt

end QualifiedLin;
