-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class PolyLoop from StepShape 

inherits Loop from StepShape 
-- WARNING : Multiple EXPRESS inheritance
-- Not yet automaticly managed
-- inherits GeometricRepresentationItem from StepShape 

uses

	HArray1OfCartesianPoint from StepGeom,
	CartesianPoint from StepGeom,
	HAsciiString from TCollection
is

	Create returns mutable PolyLoop;
	---Purpose: Returns a PolyLoop


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aPolygon : mutable HArray1OfCartesianPoint from StepGeom) is virtual;

	-- Specific Methods for Field Data Access --

	SetPolygon(me : mutable; aPolygon : mutable HArray1OfCartesianPoint);
	Polygon (me) returns mutable HArray1OfCartesianPoint;
	PolygonValue (me; num : Integer) returns mutable CartesianPoint;
	NbPolygon (me) returns Integer;

fields

	polygon : HArray1OfCartesianPoint from StepGeom;

end PolyLoop;
