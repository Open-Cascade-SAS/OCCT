-- File:	StdSelect_Shape.cdl
-- Created:	Fri Mar 27 14:46:27 1998
-- Author:	Robert COUBLANC
--		<rob@robox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1998


private class Shape from StdSelect inherits PresentableObject from PrsMgr

	---Purpose: Presentable shape only for purpose of display for BRepOwner...

uses
    Projector             from Prs3d,
    Transformation        from Geom,
    PresentationManager2d from PrsMgr,
    GraphicObject         from Graphic2d,    
    Shape                 from TopoDS,
    PresentationManager3d from PrsMgr,
    Presentation          from Prs3d

is
    Create(Sh:Shape from TopoDS) returns mutable Shape from StdSelect;
    
    Compute(me:mutable;
    	        aPresentationManager: PresentationManager3d from PrsMgr;
                aPresentation: mutable Presentation from Prs3d;
                aMode: Integer from Standard = 0)
    is redefined static;
    
    Compute(me:mutable;
    	        aProjector: Projector from Prs3d;
                aPresentation: mutable Presentation from Prs3d)
    is redefined static private;     

    Compute(me:mutable;
    	    aPresentationManager: PresentationManager2d from PrsMgr;
            aPresentation: mutable GraphicObject from Graphic2d;
            aMode: Integer from Standard = 0)
    is redefined static private;	

    Compute(me            : mutable;
    	    aProjector    : Projector from Prs3d;
    	    aTrsf         : Transformation from Geom;
	    aPresentation : mutable Presentation from Prs3d)
    is redefined;
    	---Purpose: computes the presentation according to a point of view
    	--          given by <aProjector>. 
    	--          To be Used when the associated degenerated Presentations 
    	--          have been transformed by <aTrsf> which is not a Pure
    	--          Translation. The HLR Prs can't be deducted automatically
    	--          WARNING :<aTrsf> must be applied
    	--           to the object to display before computation  !!!

    Shape(me) returns Shape from TopoDS;
    	---C++: inline
    	---C++: return const&

    Shape(me:mutable;sh : Shape from TopoDS);
    	---C++: inline

fields
    mysh : Shape  from TopoDS;
end Shape;
