-- Created by: Peter KURNEV
-- Copyright (c) 2010-2014 OPEN CASCADE SAS
-- Copyright (c) 2007-2010 CEA/DEN, EDF R&D, OPEN CASCADE
-- Copyright (c) 2003-2007 OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN, CEDRAT,
--                         EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class WireEdgeSet from BOPAlgo 

	---Purpose: 

uses
    Face   from TopoDS, 
    Shape  from TopoDS, 
    ListOfShape from BOPCol,
    BaseAllocator from BOPCol 
    
--raises

is 
    Create   
    	returns WireEdgeSet from BOPAlgo;  
    ---C++: inline  
    ---C++: alias " virtual ~BOPAlgo_WireEdgeSet();"  
     
    Create (theAllocator: BaseAllocator from BOPCol)   
    	returns WireEdgeSet from BOPAlgo;   
    ---C++: inline  
     
    Clear(me:out);
    ---C++: inline   
 
    SetFace(me:out; 
    	    aF:Face from TopoDS); 
    ---C++: inline        
    
    Face(me) 
	 returns Face from TopoDS; 
    ---C++: return const &  
    ---C++: inline    
    
    AddStartElement(me:out; 
    	    sS: Shape from TopoDS);  
    ---C++: inline       
    
    StartElements(me)  
    	returns ListOfShape from BOPCol;
    ---C++: return const & 
    ---C++: inline   
    
    AddShape(me:out; 
    	    sS:Shape from TopoDS); 
    ---C++: inline        
    
    Shapes(me)  
    	returns ListOfShape from BOPCol;
    ---C++: return const & 
    ---C++: inline   
    
fields
    myFace         : Face from TopoDS is protected; 
    myStartShapes  : ListOfShape from BOPCol is protected;
    myShapes       : ListOfShape from BOPCol is protected;  

end WireEdgeSet;
