-- Created on: 1997-09-22
-- Created by: VAUTHIER Jean-Claude
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Chamfer from QANewBRepNaming inherits TopNaming from QANewBRepNaming

    ---Purpose: To load the Chamfer results

uses 
 
    MakeChamfer from BRepFilletAPI,
    Shape       from TopoDS,
    Label       from TDF

is
 
    Create returns Chamfer from QANewBRepNaming; 

    Create(ResultLabel : Label from TDF) 
    returns Chamfer from QANewBRepNaming; 

    Init(me : in out; ResultLabel :  Label from TDF);


    Load (me; part      : in     Shape       from TopoDS;
    	      mkChamfer : in out MakeChamfer from BRepFilletAPI);

    FacesFromEdges (me) 
    ---Purpose: Returns the label of faces generated from edges
    returns Label from TDF;
    
    ModifiedFaces (me)
    ---Purpose: Returns the label of modified faces 
    returns Label from TDF;

    DeletedFaces (me)
    ---Purpose: Returns the label of deleted faces 
    returns Label from TDF;

end Chamfer;
