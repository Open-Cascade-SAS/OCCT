-- Created on: 1991-07-19
-- Created by: Isabelle GRIGNON
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


private class MyGaussFunction from CPnts 
inherits Function from math

uses
    RealFunction from CPnts

is

    Create returns MyGaussFunction;
	---C++: inline

    Init(me : in out;
    	   F : RealFunction from CPnts;
           D : Address from Standard);
	---Purpose: F  is a pointer on a  function  D is a client data
	--          
	--          Each value is computed with F(D)
    
    Value(me: in out; X : Real; F : out Real)
    returns Boolean
    is static;

fields

    myFunction : RealFunction from CPnts;
    myData     : Address      from Standard;

end MyGaussFunction;
