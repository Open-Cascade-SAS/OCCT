-- File:	BRepExtrema_ExtCC.cdl
-- Created:	Tue Feb  8 09:03:52 1994
-- Author:	Laurent PAINNOT
--		<lpa@phylox>
---Copyright:	 Matra Datavision 1994


class ExtCC from BRepExtrema

uses
    Integer from Standard,
    Real    from Standard,
    Boolean from Standard,
    Edge    from TopoDS,
    HCurve  from BRepAdaptor,
    ExtCC   from Extrema,
    Pnt     from gp
     
raises 
    NotDone      from StdFail,
    OutOfRange   from Standard,
    TypeMismatch from Standard

is
    Create returns ExtCC from BRepExtrema;

    Create(E1 : Edge from TopoDS;
           E2 : Edge from TopoDS)
    	---Purpose: It calculates all the distances.
    returns ExtCC from BRepExtrema;

    Initialize(me: in out; E2 : Edge from TopoDS)
    	---Purpose: 
    is static;
    
    Perform(me: in out; E1 : Edge from TopoDS)
    	---Purpose: An exception is raised if the fields have not been
    	--          initialized.
    raises TypeMismatch from Standard
    is static;
    
    IsDone(me) returns Boolean from Standard
    	---Purpose: True if the distances are found.
    is static;
    
    NbExt(me) returns Integer from Standard
    	---Purpose: Returns the number of extremum distances.
    raises NotDone from StdFail
    is static;

    IsParallel(me) returns Boolean from Standard
    	---Purpose: Returns True if E1 and E2 are parallel.
    raises NotDone from StdFail
    is static;
    
    SquareDistance(me; N : Integer from Standard) returns Real from Standard
    	---Purpose: Returns the value of the <N>th extremum square distance.
    raises NotDone    from StdFail,
    	   OutOfRange from Standard
    is static;
    
    ParameterOnE1(me; N : Integer from Standard) returns Real from Standard
    	---Purpose: Returns the parameter  on the first edge  of the  <N>th
    	--          extremum distance.
    raises NotDone    from StdFail,
    	   OutOfRange from Standard
    is static;
    
    PointOnE1(me; N : Integer from Standard) returns Pnt from gp
    	---Purpose: Returns the Point of the <N>th extremum distance 
    	--          on the edge E1.
    raises NotDone    from StdFail, 
    	   OutOfRange from Standard
    is static;
    
    ParameterOnE2(me; N : Integer from Standard) returns Real from Standard
    	---Purpose: Returns the parameter  on the second edge  of the  <N>th
    	--          extremum distance.
    raises NotDone    from StdFail,
    	   OutOfRange from Standard
    is static;
    
    PointOnE2(me; N : Integer from Standard) returns Pnt from gp
    	---Purpose: Returns the Point of the <N>th extremum distance 
    	--          on the edge E2.
    raises NotDone    from StdFail, 
    	   OutOfRange from Standard
    is static;
    
    
    TrimmedSquareDistances(me; dist11, distP12, distP21, distP22: out Real;
                     P11, P12, P21, P22: out Pnt)
    	---Purpose: if the edges is a trimmed curve,
    	--          dist11 is a square distance between the point on E1
    	--          of parameter FirstParameter and the point of 
    	--          parameter FirstParameter on E2.

    is static;

    
fields
    myExtrem  : ExtCC   from Extrema;
    myHC      : HCurve  from BRepAdaptor;    
end ExtCC;
