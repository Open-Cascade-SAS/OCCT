-- Created on: 1994-08-03
-- Created by: Christophe MARION
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class OutLiner from HLRTopoBRep inherits TShared from MMgt

uses
    Integer        from Standard,
    Shape          from TopoDS,
    Face           from TopoDS,
    Projector      from HLRAlgo,
    Data           from HLRTopoBRep,
    MapOfShapeTool from BRepTopAdaptor
is
    Create
    returns mutable OutLiner from HLRTopoBRep;

    Create (OriSh : Shape from TopoDS)
    returns mutable OutLiner from HLRTopoBRep;

    Create (OriS : Shape from TopoDS;
            OutS : Shape from TopoDS)
    returns mutable OutLiner from HLRTopoBRep;

    OriginalShape(me : mutable; OriS : Shape from TopoDS)
    	---C++: inline
    is static;

    OriginalShape(me : mutable) returns Shape from TopoDS
    	---C++: inline
    	---C++: return &
    is static;

    OutLinedShape(me : mutable; OutS : Shape from TopoDS)
    	---C++: inline
    is static;

    OutLinedShape(me : mutable) returns Shape from TopoDS
    	---C++: inline
    	---C++: return &
    is static;

    DataStructure(me : mutable) returns Data from HLRTopoBRep
    	---C++: inline
    	---C++: return &
    is static;

    Fill(me : mutable;
         P     :        Projector      from HLRAlgo;
	 MST   :in out  MapOfShapeTool from BRepTopAdaptor;
         nbIso :        Integer        from Standard)
    is static;
    
    ProcessFace(me : mutable; F :        Face           from TopoDS;
                              S : in out Shape          from TopoDS;
                              M : in out MapOfShapeTool from BRepTopAdaptor)  
	---Purpose: Builds faces from F and add them to S.
    is static private;

    BuildShape(me : mutable; M : in out MapOfShapeTool from BRepTopAdaptor)
    is static private;
    
fields
    myOriginalShape : Shape from TopoDS;
    myOutLinedShape : Shape from TopoDS;
    myDS            : Data  from HLRTopoBRep;

end OutLiner;
