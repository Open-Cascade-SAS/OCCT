-- Created on: 1995-09-05
-- Created by: Christian CAILLET
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class SelectFlag  from IFSelect  inherits SelectExtract

    ---Purpose : A SelectFlag queries a flag noted in the bitmap of the Graph.
    --           The Flag is designated by its Name. Flag Names are defined
    --           by Work Session and, as necessary, other functional objects
    --           
    --           WorkSession from IFSelect defines flag "Incorrect"
    --           Objects which control application running define some others

uses AsciiString from TCollection, InterfaceModel, Graph, EntityIterator

is

    Create (flagname : CString) returns mutable SelectFlag;
    ---Purpose : Creates a Select Flag, to query a flag designated by its name

    FlagName (me) returns CString;
    ---Purpose : Returns the name of the flag

    RootResult (me; G : Graph) returns EntityIterator  is redefined;
    ---Purpose : Returns the list of selected entities. It is redefined to
    --           work on the graph itself (not queried by sort)
    --           
    --           An entity is selected if its flag is True on Direct mode,
    --           False on Reversed mode
    --           
    --           If flag does not exist for the given name, returns an empty
    --           result, whatever the Direct/Reversed sense

    Sort (me; rank : Integer; ent : Transient; model : InterfaceModel)
        returns Boolean;
    ---Purpose : Returns always False because RootResult has done the work


    ExtractLabel (me) returns AsciiString from TCollection;
    ---Purpose : Returns a text defining the criterium, includes the flag name

fields

    thename : AsciiString from TCollection;

end SelectFlag;
