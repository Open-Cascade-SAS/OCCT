-- File:        SurfaceStyleElementSelect.cdl
-- Created:     Fri Dec  1 11:11:11 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993



class SurfaceStyleElementSelect from StepVisual inherits SelectType from StepData

	-- <SurfaceStyleElementSelect> is an EXPRESS Select Type construct translation.
	-- it gathers : SurfaceStyleFillArea, SurfaceStyleBoundary, SurfaceStyleSilhouette, SurfaceStyleSegmentationCurve, SurfaceStyleControlGrid, SurfaceStyleParameterLine
	-- Rev4 : only remain SurfaceStyleFillArea, SurfaceStyleBoundary, SurfaceStyleParameterLine

uses

	SurfaceStyleFillArea,
	SurfaceStyleBoundary,
--	SurfaceStyleSilhouette,
--	SurfaceStyleSegmentationCurve,
--	SurfaceStyleControlGrid,
	SurfaceStyleParameterLine
is

	Create returns SurfaceStyleElementSelect;
	---Purpose : Returns a SurfaceStyleElementSelect SelectType

	CaseNum (me; ent : Transient) returns Integer;
	---Purpose: Recognizes a SurfaceStyleElementSelect Kind Entity that is :
	--        1 -> SurfaceStyleFillArea
	--        2 -> SurfaceStyleBoundary
	--        3 -> SurfaceStyleParameterLine
	--        4 -> SurfaceStyleSilhouette
	--        5 -> SurfaceStyleSegmentationCurve
	--        6 -> SurfaceStyleControlGrid
	--        0 else

	SurfaceStyleFillArea (me) returns any SurfaceStyleFillArea;
	---Purpose : returns Value as a SurfaceStyleFillArea (Null if another type)

	SurfaceStyleBoundary (me) returns any SurfaceStyleBoundary;
	---Purpose : returns Value as a SurfaceStyleBoundary (Null if another type)

	SurfaceStyleParameterLine (me) returns any SurfaceStyleParameterLine;
	---Purpose : returns Value as a SurfaceStyleParameterLine (Null if another type)


end SurfaceStyleElementSelect;

