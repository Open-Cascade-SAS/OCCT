-- Created on: 1993-08-24
-- Created by: Bruno DUMORTIER
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Sphere from ProjLib inherits Projector from ProjLib

	---Purpose: Projects elementary curves on a sphere.

uses
    CurveType  from GeomAbs,
    Sphere     from gp,
    Lin        	   from gp,
    Circ       	   from gp,
    Elips      	   from gp,
    Parab      	   from gp,
    Hypr       	   from gp,
    Lin2d      from gp,
    Circ2d     from gp,
    Elips2d    from gp,
    Parab2d    from gp,
    Hypr2d     from gp

raises
    NoSuchObject from Standard

is

    Create returns Sphere from ProjLib;
	---Purpose: Undefined projection.

    Create(Sp : Sphere from gp) returns Sphere from ProjLib;
	---Purpose: Projection on the sphere <Sp>.

    Create(Sp : Sphere  from gp;
           C  : Circ from gp) returns Sphere from ProjLib;
	---Purpose: Projection of the circle <C> on the sphere <Sp>.



    Init(me : in out;
    	 Sp : Sphere from gp)
    is static;
	 
     Project(me : in out;
     	     L  : Lin from gp)
     is redefined;
 
    Project(me : in out;
    	    C  : Circ from gp)
    is redefined;

     Project(me : in out;
     	     E  : Elips from gp)
     is redefined;
 
     Project(me : in out;
     	     P  : Parab from gp)
     is redefined;
 
     Project(me : in out;
     	     H  : Hypr from gp)
     is redefined;
	     
    SetInBounds(me: in out;
    	    	U : Real from Standard)
    	---Purpose: Set the point of parameter U on C in the natural
    	--          restrictions of the sphere.
    is static;		
    

fields

    mySphere : Sphere from gp;

end Sphere;
