-- Created on: 1996-09-04
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Pipe from LocOpe 

	---Purpose: Defines a  pipe  (near from   Pipe from BRepFill),
	--          with modifications provided for the Pipe feature.

uses Pipe from BRepFill,

     ListOfShape               from TopTools,
     DataMapOfShapeListOfShape from TopTools,
     Curve                     from  Geom,      
     Shape                     from TopoDS,
     Wire                      from TopoDS,     
     SequenceOfPnt             from TColgp,
     SequenceOfCurve           from TColGeom
     

raises NoSuchObject from Standard,
       DomainError  from Standard

is

    Create (Spine   : Wire from TopoDS;
    	    Profile : Shape from TopoDS)
	    
    	returns Pipe from LocOpe;


    Spine(me)
    
    	returns Shape from TopoDS
	---C++: inline
	---C++: return const &
	is static;


    Profile(me)
    
    	returns Shape from TopoDS
	---C++: inline
	---C++: return const &
	is static;


    FirstShape(me)
    
    	returns Shape from TopoDS
	---C++: inline
	---C++: return const &
	is static;


    LastShape(me)
    
    	returns Shape from TopoDS
	---C++: inline
	---C++: return const &
	is static;


    Shape(me)
    
    	returns Shape from TopoDS
	---C++: return const &
	is static;


    Shapes(me: in out; S: Shape from TopoDS)
    
    	returns ListOfShape from TopTools
	---C++: return const &
    	raises NoSuchObject from Standard,
	       -- The exception is raised if S is not a subshape of the profile
               DomainError  from Standard
	       -- The exception is raised if S is neither a vertex nor
	       -- an edge
	is static;


    Curves(me: in out; Spt: SequenceOfPnt from TColgp)

	---C++: return const &
    	returns SequenceOfCurve from TColGeom
	is static;

    BarycCurve(me: in out) 
     
    	returns  Curve  from  Geom 
	is  static;

fields

    myPipe : Pipe                      from BRepFill;
    myMap  : DataMapOfShapeListOfShape from TopTools;
    myRes  : Shape                     from TopoDS;
    myGShap: ListOfShape               from TopTools;
    myCrvs : SequenceOfCurve           from TColGeom;
    myFirstShape : Shape             from TopoDS;
    myLastShape  : Shape             from TopoDS;

end Pipe;
