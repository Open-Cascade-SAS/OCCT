-- Created on: 1992-05-05
-- Created by: Remi GILET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package GCE2d

uses gp,
     Geom2d,
     gce,
     StdFail


    ---Level : Public. 
    --  All methods of all  classes will be public.



is

private deferred class Root;

---------------------------------------------------------------------------
--          Constructions of 2d geometrical elements from Geom2d.
---------------------------------------------------------------------------

class MakeLine;

class MakeCircle;

class MakeHyperbola;

class MakeEllipse;

class MakeParabola;

class MakeSegment;

class MakeArcOfCircle;

class MakeArcOfEllipse;

class MakeArcOfParabola;

class MakeArcOfHyperbola;

---------------------------------------------------------------------------
--              Constructions of Transformation from Geom2d.
---------------------------------------------------------------------------

class MakeTranslation;
 
class MakeMirror;

class MakeRotation;

class MakeScale;

    
end GCE2d;



