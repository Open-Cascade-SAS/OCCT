-- Created on: 1993-01-12
-- Created by: Philippe DAUTRY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



package BRepSweep

    ---Purpose: This package implements the package Sweep for the BRep
    --          structure.

uses

    Standard,
    Quantity,
    TCollection, 
    TColStd,
    gp, 
    Geom,
    TopAbs, 
    TopLoc, 
    TopTools, 
    TopoDS, 
    TopExp, 
    BRep,
    Sweep

is

    class Builder;
	---Purpose: Implements the Builder required for Sweep.

    class Tool;
	---Purpose: Provides an indexation of the subShapes of a Shape
	--          from TopoDS.
	
    class Iterator;
	---Purpose: Iterator on the subShapes of a shape.
	

    deferred class NumLinearRegularSweep
    	instantiates LinearRegularSweep from Sweep(
    	Shape              from TopoDS,     -- Resulting topological objects.
    	Shape              from TopoDS,     -- Generating Shape.
    	NumShape           from Sweep,      -- Directing Wire.
    	Builder            from BRepSweep,
    	Tool               from BRepSweep,  -- GenTool
	NumShapeTool       from Sweep,      -- DirTool
    	Iterator           from BRepSweep,  -- Resulting objects Iterator
    	Iterator           from BRepSweep,  -- GenIterator
	NumShapeIterator   from Sweep);     -- DirSubEdgeIterator

    deferred class Trsf;
    --- This class is inherited  from LinearRegularSweep to  implement
    --  the simple swept primitives built moving a Shape with a Trsf.

    class Translation;
    --- This class is inherited from Trsf to implement the translation
    --  sweep.

    class Rotation;
    --- This class is  inherited  from Trsf to implement  the rotation
    --  sweep.

    class Prism;
    --- This class provides simple methods to build prism.

    class Revol;
    --- This class provides simple methods to build Revol.

end BRepSweep;
