-- File:	IGESSolid_SpecificModule.cdl
-- Created:	Tue Sep  7 11:14:37 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class SpecificModule  from IGESSolid  inherits  SpecificModule from IGESData

    ---Purpose : Defines Services attached to IGES Entities : Dump, for IGESSolid

uses Messenger from Message, IGESEntity, IGESDumper

is

    Create returns mutable SpecificModule from IGESSolid;
    ---Purpose : Creates a SpecificModule from IGESSolid & puts it into SpecificLib

    OwnDump (me; CN : Integer; ent : IGESEntity;
    	      dumper : IGESDumper;  S : Messenger from Message; own : Integer);
    ---Purpose : Specific Dump (own parameters) for IGESSolid

end SpecificModule;
