-- File:	BRepLProp_SurfaceTool.cdl
-- Created:	Thu Feb 24 10:40:20 1994
-- Author:	Laurent BOURESCHE
--		<lbo@nonox>
---Copyright:	 Matra Datavision 1994

class SurfaceTool from BRepLProp

uses Pnt     from gp,
     Vec     from gp,
     Surface from BRepAdaptor

is

    Value(myclass; S : Surface; U, V : Real; P : out Pnt);
    ---Purpose: Computes the point <P> of parameter <U> and <V> on the 
    --          Surface <S>.
     	
    D1   (myclass; S : Surface; U, V : Real; P : out Pnt; D1U, D1V : out Vec);
    ---Purpose: Computes the point <P> and first derivative <D1*> of 
    --          parameter <U> and <V> on the Surface <S>.

    D2   (myclass; S : Surface; U, V : Real; 
              P : out Pnt; D1U, D1V, D2U, D2V, DUV : out Vec);
    ---Purpose: Computes the point <P>, the first derivative <D1*> and second
    --          derivative <D2*> of parameter <U> and <V> on the Surface <S>.
              
   DN     (myclass; S : Surface; U, V : Real;  IU,  IV  :  Integer) 
   returns  Vec;
     
    Continuity(myclass; S : Surface) returns Integer;
    ---Purpose: returns the order of continuity of the Surface <S>.
    --          returns 1 : first derivative only is computable
    --          returns 2 : first and second derivative only are computable.

    Bounds(myclass; S : Surface; U1, V1, U2, V2 : out Real);
    ---Purpose: returns the bounds of the Surface.

end SurfaceTool;


