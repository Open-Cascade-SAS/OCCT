-- File:	StdSchema.cdl
-- Created:	Sep 7 14:00:00 2000
-- Author:	TURIN Anatoliy
---Copyright:	Matra Datavision 2000

schema StdSchema

is
    package PDataXtd;
    package PNaming;    
    package PPrsStd;
    
end StdSchema;

