-- Created on: 1991-07-24
-- Created by: Michel CHAUVAT
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Modified by skv - Thu Sep 30 15:19:59 2004 OCC593


private class FuncExtPS from Extrema

 inherits FunctionSetWithDerivatives from math
    ---Purpose: 
    --
    -- Functional for search of extremum of the distance between point P and 
    -- surface S, starting from approximate solution (u0, v0).
    --          
    -- The class inherits math_FunctionSetWithDerivatives and thus is intended
    -- for use in math_FunctionSetRoot algorithm .
    --          
    -- Denoting derivatives of the surface S(u,v) by u and v, respectively, as 
    -- Su and Sv, the two functions to be nullified are:
    --          
    -- F1(u,v) = (S - P) * Su
    -- F2(u,v) = (S - P) * Sv
    --          
    -- The derivatives of the functional are:
    --          
    -- Duf1(u,v) = Su^2    + (S-P) * Suu;
    -- Dvf1(u,v) = Su * Sv + (S-P) * Suv
    -- Duf2(u,v) = Sv * Su + (S-P) * Suv = Dvf1
    -- Dvf2(u,v) = Sv^2    + (S-P) * Svv
    --
    -- Here * denotes scalar product, and ^2 is square power. 

uses    POnSurf           from Extrema,
	SequenceOfPOnSurf from Extrema,
	SequenceOfReal    from TColStd,
	Pnt               from gp,
	Vector            from math,
	Matrix            from math,
	Surface           from Adaptor3d,
    	SurfacePtr        from Adaptor3d

raises  OutOfRange from Standard

is
    Create returns FuncExtPS;

    Create (P: Pnt; S: Surface from Adaptor3d) returns FuncExtPS;
    	---Purpose:

    Initialize(me: in out; S: Surface from Adaptor3d)
    	---Purpose: sets the field mysurf of the function.
    is static;
    
    SetPoint(me: in out; P: Pnt)
    	---Purpose: sets the field mysurf of the function.
    is static;

    ------------------------------------------------------------
    -- In all next methods, an exception is raised if the fields 
    -- were not initialized.

    NbVariables (me) returns Integer;

    NbEquations (me) returns Integer;

    Value (me: in out; UV: Vector; F: out Vector) returns Boolean;
    	---Purpose: Calculate Fi(U,V).

    Derivatives (me: in out; UV: Vector; DF: out Matrix)
    	returns Boolean;
    	---Purpose: Calculate Fi'(U,V).

    Values (me: in out; UV: Vector; F: out Vector; DF: out Matrix)
    	returns Boolean;
    	---Purpose: Calculate Fi(U,V) and Fi'(U,V).

    GetStateNumber (me: in out) returns Integer
    	---Purpose: Save the found extremum.
    	is redefined;

    NbExt (me) returns Integer;
    	---Purpose: Return the number of found extrema.

    SquareDistance (me; N: Integer) returns Real
    	---Purpose: Return the value of the Nth distance.
    	raises  OutOfRange;
	    	-- if N < 1 or N > NbExt(me).

    Point (me; N: Integer) returns POnSurf
        ---C++: return const &
    	---Purpose: Returns the Nth extremum.
    	raises  OutOfRange;
	    	-- if N < 1 or N > NbExt(me).

fields
    myP    : Pnt from gp;
    myS    : SurfacePtr from Adaptor3d;

    myU    : Real;          -- current value of U
    myV    : Real;          -- current value of V
    myPs   : Pnt from gp;   -- current point

    mySqDist: SequenceOfReal    from TColStd;
    myPoint: SequenceOfPOnSurf from Extrema;
    myPinit: Boolean;
    mySinit: Boolean;

end FuncExtPS;
