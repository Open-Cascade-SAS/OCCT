-- Created on: 1993-06-14
-- Created by: Martine LANGLOIS
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MakeAxis1Placement from GeomToStep inherits Root from GeomToStep

    ---Purpose: This class implements the mapping between classes 
    --          Axis1Placement from Geom and Ax1 from gp, and the class
    --          Axis1Placement from StepGeom which describes an
    --          Axis1Placement from Prostep. 
    --         
  
uses Ax1 from gp,
     Ax2d from gp,
     Axis1Placement from Geom,
     AxisPlacement from Geom2d,
     Axis1Placement from StepGeom
     
raises NotDone from StdFail
     
is 

Create ( A : Ax1 from gp ) returns MakeAxis1Placement;

Create ( A : Ax2d from gp ) returns MakeAxis1Placement;

Create ( A : Axis1Placement from Geom ) returns MakeAxis1Placement;

Create ( A : AxisPlacement from Geom2d ) returns MakeAxis1Placement;

Value (me) returns Axis1Placement from StepGeom
    raises NotDone
    is static;
    ---C++: return const&

fields

    theAxis1Placement : Axis1Placement from StepGeom;
    	-- The solution from StepGeom
    	
end MakeAxis1Placement;


