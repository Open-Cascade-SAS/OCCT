-- Created on: 2001-07-17
-- Created by: Julia DOROVSKIKH <jfa@hotdox.nnov.matra-dtv.fr>
-- Copyright (c) 2001-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Persistent from XmlObjMgt

uses
    Element from XmlObjMgt,
    DOMString from XmlObjMgt

is
    Create      returns Persistent from XmlObjMgt;
      ---Purpose: empty constructor

    Create (theElement : Element from XmlObjMgt)
                returns Persistent from XmlObjMgt;
      ---Purpose: constructor

    Create (theElement : Element from XmlObjMgt;
            theRef     : DOMString from XmlObjMgt)
                returns Persistent from XmlObjMgt;
      ---Purpose: constructor from sub-element of Element referenced by theRef

    CreateElement (me:in out; theParent: out Element   from XmlObjMgt;
                              theType:       DOMString from XmlObjMgt;
                              theID:         Integer   from Standard);
      ---Purpose: myElement := <theType id="theID"/>

    SetId (me:in out; theId: Integer from Standard)
    is static;
      ---Level: Internal

    Element (me) returns Element from XmlObjMgt;
      ---C++: inline
      ---C++: return const &
      ---C++: alias "inline operator const XmlObjMgt_Element&() const;"
      ---Purpose: return myElement

    Element (me:in out) returns Element from XmlObjMgt;
      ---C++: inline
      ---C++: return &
      ---C++: alias "inline operator XmlObjMgt_Element&();"
      ---Purpose: return myElement

    Id(me) returns Integer from Standard
    is static;
      ---C++: inline
      ---Level: Internal

fields
    myElement: Element from XmlObjMgt;
    myID     : Integer from Standard;

end Persistent;
