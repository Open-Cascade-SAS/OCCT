-- Created on: 1993-05-05
-- Created by: Christian CAILLET
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class Protocol  from IGESDimen  inherits  Protocol from IGESData

    ---Purpose : Description of Protocol for IGESDimen

uses Type, Protocol from Interface

is

    Create returns mutable Protocol from IGESDimen;

    NbResources (me) returns Integer  is redefined;
    ---Purpose : Gives the count of Resource Protocol. Here, two
    --           (Protocols from IGESGraph and IGESGeom)

    Resource (me; num : Integer) returns Protocol from Interface  is redefined;
    ---Purpose : Returns a Resource, given a rank.

    TypeNumber (me; atype : any Type) returns Integer  is redefined;
    ---Purpose : Returns a Case Number, specific of each recognized Type
    --           This Case Number is then used in Libraries : the various
    --           Modules attached to this class of Protocol must use them
    --           in accordance (for a given value of TypeNumber, they must
    --           consider the same Type as the Protocol defines)

end Protocol;
