-- File:        Axis1Placement.cdl
-- Created:     Fri Dec  1 11:11:14 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class Axis1Placement from StepGeom 

inherits Placement from StepGeom 

uses

	Direction from StepGeom, 
	Boolean from Standard, 
	HAsciiString from TCollection, 
	CartesianPoint from StepGeom
is

	Create returns mutable Axis1Placement;
	---Purpose: Returns a Axis1Placement


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aLocation : mutable CartesianPoint from StepGeom) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aLocation : mutable CartesianPoint from StepGeom;
	      hasAaxis : Boolean from Standard;
	      aAxis : mutable Direction from StepGeom) is virtual;

	-- Specific Methods for Field Data Access --

	SetAxis(me : mutable; aAxis : mutable Direction);
	UnSetAxis (me:mutable);
	Axis (me) returns mutable Direction;
	HasAxis (me) returns Boolean;

fields

	axis : Direction from StepGeom;   -- OPTIONAL can be NULL
	hasAxis : Boolean from Standard;

end Axis1Placement;
