-- Created on: 1993-03-01
-- Created by: Philippe DAUTRY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class TrimmedCurve from PGeom inherits BoundedCurve from PGeom

        ---Purpose :
        --  Defines a portion of a curve limited by two values of 
        --  parameters inside the parametric domain of the curve.
        --  
	---See Also : TrimmedCurve from Geom.


uses Curve from PGeom

is


  Create returns mutable TrimmedCurve from PGeom;
	---Purpose: Creates a TrimmedCurve with default values.
    	---Level: Internal 


  Create (
    	aBasisCurve: Curve from PGeom;
    	aFirstU, aLastU: Real from Standard)
     returns mutable TrimmedCurve from PGeom;
        ---Purpose : Creates a TrimmedCurve with these field values.
    	---Level: Internal 


  FirstU(me : mutable; aFirstU: Real from Standard);
        ---Purpose : Set the value of the field firstU with <aFirstU>.
    	---Level: Internal 


  FirstU(me) returns Real from Standard;
        ---Purpose : Returns the value of the field firstU.
    	---Level: Internal 


  LastU(me : mutable; aLastU: Real from Standard);
        ---Purpose : Set the value of the field lastU with <aLastU>.
    	---Level: Internal 


  LastU(me) returns Real from Standard;
        ---Purpose : Returns the value of the field lastU.
    	---Level: Internal 


  BasisCurve (me: mutable; aBasisCurve: Curve from PGeom);
        ---Purpose : Set the value of the field basisCurve with <aBasisCurve>.
        --  This curve can be a trimmed curve.
    	---Level: Internal 


  BasisCurve (me) returns Curve from PGeom;
        ---Purpose : Returns the value of the field basisCurve. 
        --  This curve can be a trimmed curve.
    	---Level: Internal 


fields

    basisCurve : Curve from PGeom;
    firstU     : Real from Standard;
    lastU      : Real from Standard;

end;
