-- Created on: 1993-04-06
-- Created by: Philippe DAUTRY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package PGeom2d 

        ---Purpose :  This  package contains   the definition   of the
        --         geometric persistent objects such as point, vector,
        --         axis placement, curves, surfaces.
        --  
        --  All these entities are defined in 2D space.
        --  This package gives the possibility :
        --    . to create geometric objects with given or default field values,
        --    . to set field values,
        --    . to get field values.


uses PColStd, gp, PColgp, GeomAbs

is


  class Transformation from PGeom2d;


  deferred class Geometry from PGeom2d;


     deferred class Point from PGeom2d;
              class  CartesianPoint from PGeom2d;


     deferred class Vector from PGeom2d;
              class Direction from PGeom2d;
              class VectorWithMagnitude from PGeom2d;
     

     class AxisPlacement from PGeom2d;


     deferred class Curve from PGeom2d;

              class Line from PGeom2d;

              deferred class Conic from PGeom2d;
                       class Circle from PGeom2d;
                       class Ellipse from PGeom2d;
                       class Hyperbola from PGeom2d;
                       class Parabola from PGeom2d;

              deferred class BoundedCurve from PGeom2d;
                       class BezierCurve from PGeom2d;
                       class BSplineCurve from PGeom2d;
                       class TrimmedCurve from PGeom2d;

              class  OffsetCurve from PGeom2d;

end PGeom2d;
