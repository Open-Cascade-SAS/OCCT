-- Created on: 1998-01-17
-- Created by: Julia GERASIMOVA
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class EqualRadiusPresentation from DsgPrs 

	---Purpose: A framework to define display of equality in radii.

uses
    Presentation from Prs3d,
    Drawer from Prs3d,
    Pnt from gp,
    Plane from Geom
    
is
    Add( myclass; aPresentation : Presentation from Prs3d;
    	    	  aDrawer       : Drawer from Prs3d;
		  FirstCenter   : Pnt from gp;
		  SecondCenter  : Pnt from gp;
		  FirstPoint    : Pnt from gp;
		  SecondPoint   : Pnt from gp; 
		  Plane         : Plane from Geom );
	---Purpose: Adds the points FirstCenter, SecondCenter,
    	-- FirstPoint, SecondPoint, and the plane Plane to the
    	-- presentation object aPresentation.
    	-- The display attributes of these elements is defined by
    	-- the attribute manager aDrawer.
    	-- FirstCenter and SecondCenter are the centers of the
    	-- first and second shapes respectively, and FirstPoint
    	-- and SecondPoint are the attachment points of the radii to arcs.
    	    	    
end EqualRadiusPresentation;
