-- Created on: 1993-06-02
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred generic class SOBFunction from IntStart 
    (TheArc as any)

inherits FunctionWithDerivative from math 


	---Purpose: Template class for the function on an arc of restriction
	--          used in the SearchOnBoundaries class.

uses Pnt from gp


is


    Set(me: in out; A: TheArc)
    
    	is static;


    Value(me: in out; X: Real from Standard; F: out Real from Standard)
    
    	returns Boolean from Standard;
    
    Derivative(me: in out; X: Real from Standard; D: out Real from Standard)
    
    	returns Boolean from Standard;
    
    Values(me: in out; X: Real from Standard; F,D: out Real from Standard)
    
    	returns Boolean from Standard;
    

    GetStateNumber(me: in out)

    	returns Integer from Standard

    	is redefined;
	
	
    Valpoint(me; Index: Integer from Standard)
    
    	returns Pnt from gp
	
	is static;
    

end SOBFunction;
