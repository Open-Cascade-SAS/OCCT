-- Created on: 1995-05-04
-- Created by: Dieter THIEMANN
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MakeParabola from GeomToStep inherits Root from GeomToStep

    ---Purpose: This class implements the mapping between the class
    --          Parabola from Geom and the class Parabola from
    --          StepGeom which describes a Parabola from ProSTEP


uses Parabola from Geom,
     Parabola from Geom2d,
     Parabola from StepGeom
     
raises NotDone from StdFail

is

Create ( C : Parabola from Geom2d) returns MakeParabola;

Create ( C : Parabola from Geom) returns MakeParabola;


Value (me) returns Parabola from StepGeom
    raises NotDone
    is static;
    ---C++: return const&


fields

    theParabola : Parabola from StepGeom;
    	-- The solution from StepGeom

end MakeParabola;
