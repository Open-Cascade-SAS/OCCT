-- File:	MakeTranslation.cdl
-- Created:	Mon Sep 28 11:52:25 1992
-- Author:	Remi GILET
--		<reg@sdsun2>
---Copyright:	 Matra Datavision 1992

class MakeTranslation

from GC

    	---Purpose: This class mplements elementary construction algorithms for a
    	-- translation in 3D space. The result is a
    	-- Geom_Transformation transformation.
    	-- A MakeTranslation object provides a framework for:
    	-- -   defining the construction of the transformation,
    	-- -   implementing the construction algorithm, and
    	-- -   consulting the result.

uses Pnt            from gp,
     Transformation from Geom,
     Vec            from gp,
     Real           from Standard
     
is

Create(Vect : Vec from gp) returns MakeTranslation;
    	---Purpose: Constructs a translation along the vector " Vect "        
Create(Point1 : Pnt from gp;
       Point2 : Pnt from gp) returns MakeTranslation;
    	---Purpose: Constructs a translation along the vector (Point1,Point2)
    	--  defined from the point Point1 to the point Point2.
    
Value(me) returns Transformation from Geom
    is static;
    	---Purpose:  Returns the constructed transformation.
    	---C++: return const&

Operator(me) returns Transformation from Geom
    is static;
    	---C++: return const&
    	---C++: alias "Standard_EXPORT operator Handle_Geom_Transformation() const;"

fields

    TheTranslation : Transformation from Geom;

end MakeTranslation;

