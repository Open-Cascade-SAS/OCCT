-- Created on: 1993-07-27
-- Created by: Jean Louis FRENKEL
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class PseudoColorImage from Image inherits DIndexedImage from Image

	---Purpose : A PseudoColorImage is a DIndexedImage associated with a
	--	     ColorMap . The ColoMap is set at Creation time and then
	--	     never be changed. Each Pixel in the Image ,as a IndexPixel
	--	     from Aspect, match a ColoMap Entry with the same value.

uses
    ColorMap 		from Aspect,
    Color    		from Quantity,
    IndexPixel 		from Aspect ,
    Array1OfColor 	from Quantity,
    HArray1OfColor 	from Quantity,
    LookupTable  	from Image,
    Image 		from Image,
    TypeOfImage 	from Image
    
is

    Create( x,y,dx,dy   : in Integer from Standard ;
            aColorMap   : ColorMap   from Aspect )
    	returns mutable PseudoColorImage from Image;
	---Level: Public
	---Purpose : Creates a PseudoColorImage object.
	--	       The default Background Pixel is set to 0 .
	--	       All the Image is initialised with Background Pixel
    
    Create( x,y,dx,dy   : in Integer from Standard ;
            aColorMap   : ColorMap   from Aspect ;
	    BackPixel   : IndexPixel from Aspect )
    	returns mutable PseudoColorImage from Image;
	---Level: Public
	---Purpose : Creates a PseudoColorImage object and set the 
	--	       Background Pixel.
	--	       All the Image is initialised with Background Pixel
    
    Type    ( me : immutable )  returns TypeOfImage from Image ;
	---Level: Public
	---Purpose : Returns the Image Type.

    ColorMap( me ) returns immutable ColorMap from Aspect;
	---Level: Public
	---Purpose : returns the Image ColorMap .

    PixelColor( me : immutable ; X,Y : in Integer from Standard ) 
	returns Color from Quantity ;
    	---C++: return const &
	---Level: Public
	---Purpose : Returns the Pixel Color .

    RowColor  ( me : immutable ; Y : in Integer from Standard )
	returns HArray1OfColor from Quantity is redefined ;
	---Level: Public
	---Purpose : Return the PixelRow Color in a HArray1 of Color.

    RowColor  ( me       : immutable ; 
		Y        : in Integer from Standard ;
		aArray1  : in out Array1OfColor from Quantity ) is redefined ;
	---Level: Public
	---Purpose : Stores the PixelRow Color in a Array1 .

    Squeeze( 	me 		: immutable ; 
		BasePixel 	: IndexPixel from Aspect ) 
	returns PseudoColorImage from Image ;
	---Level: Public
	---Purpose : Creates a new Image with continuous Pixel and a continuous 
	--              ColorMap whith only used Image color starting from
	--		BasePixel .

    SqueezedLookupTable( 
		me 		: immutable ; 
		BasePixel 	: IndexPixel from Aspect ;
		aLookup		: in out LookupTable from Image ) ;
	---Level: Public
	---Purpose: Creates a LookupTable that can be used to create a
	--	    new Image with continuous Pixel and a continuous 
	--	    ColorMap with only used Image color starting
	--	    from BasePixel .

    Lookup( me : mutable ; 
	    aLookup : in LookupTable from Image ) ;
	---Level: Public
	---Purpose : Pass a PseudoColorImage through a lookupTable

    Extrema( me : immutable ; Min, Max : in out IndexPixel from Aspect );
	---Level: Public
	---Purpose: Find the maximum and minimum Pixel Value of an Image.

    Threshold( me : mutable ; Min, Max : IndexPixel from Aspect ;
			      Map      : IndexPixel from Aspect );
	---Level: Public
	---Purpose: This method changes the value of any Pixel beetwen the 
	--	    range (Min->Max) to the Pixel Map value. All Pixel values
	--	    outside the range are passed through without changed .

    Rescale( me : mutable ; Scale, Offset : Real from Standard ) ;
	---Level: Public
	---Purpose : Map the Image Pixel Value from one range to another range.
	--	     This method perform the mapping by multiplying each
	--	     Pixel Value by Scale and then adding Offset to the result.

    Dup   ( me : immutable ) returns mutable Image from Image;
	---Level: Public
	---Purpose : Duplicate a Image.

    -- ******************* Redefined method  *************************** 

--	ShallowCopy (me) returns mutable like me  ;
	---Level: Public
--	    ---Purpose: Returns a copy at the first level of <me>. The objects 
--	    --         referenced are not copied. Entities copied by 
--	    --         ShallowCopy are equal.
--	    ---C++:  function call

--	DeepCopy (me) returns mutable like me  ;
	---Level: Public
--	    ---Purpose: Returns a deep copy of <me>. The objects 
--	    --          referenced are copied. Entities copied by 
--	    --          DeepCopy are similar (c.f the Method IsSimilar).
--	    ---C++:  function call

fields
    myColorMap: ColorMap from Aspect;
    
end PseudoColorImage from Image;
