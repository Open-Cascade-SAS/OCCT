-- Created on: 1993-04-28
-- Created by: Laurent PAINNOT
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred generic class TheSurfTool from AppCont(Surf as any)

    ---Purpose: Template for describing a continuous surface.


uses Pnt           from gp,
     Vec           from gp

is


    D0(myclass; S: Surf; U, V: Real; Pt: out Pnt);
    	---Purpose: returns the point of the surface at <U, V>.


    D1(myclass; S: Surf; U, V: Real; Pt: out Pnt; V1U, V1V: out Vec);
    	---Purpose: returns the derivative and the point values of the surface
    	--          at the parameters <U, V> .

end TheSurfTool;
