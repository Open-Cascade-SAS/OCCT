-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Product from StepBasic 

inherits TShared from MMgt

uses

	HAsciiString from TCollection, 
	HArray1OfProductContext from StepBasic, 
	ProductContext from StepBasic
is

	Create returns mutable Product;
	---Purpose: Returns a Product

	Init (me : mutable;
	      aId : mutable HAsciiString from TCollection;
	      aName : mutable HAsciiString from TCollection;
	      aDescription : mutable HAsciiString from TCollection;
	      aFrameOfReference : mutable HArray1OfProductContext from StepBasic) is virtual;

	-- Specific Methods for Field Data Access --

	SetId(me : mutable; aId : mutable HAsciiString);
	Id (me) returns mutable HAsciiString;
	SetName(me : mutable; aName : mutable HAsciiString);
	Name (me) returns mutable HAsciiString;
	SetDescription(me : mutable; aDescription : mutable HAsciiString);
	Description (me) returns mutable HAsciiString;
	SetFrameOfReference(me : mutable; aFrameOfReference : mutable HArray1OfProductContext);
	FrameOfReference (me) returns mutable HArray1OfProductContext;
	FrameOfReferenceValue (me; num : Integer) returns mutable ProductContext;
	NbFrameOfReference (me) returns Integer;

fields

	id : HAsciiString from TCollection;
	name : HAsciiString from TCollection;
	description : HAsciiString from TCollection;
	frameOfReference : HArray1OfProductContext from StepBasic;

end Product;
