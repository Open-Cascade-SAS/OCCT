-- Created on: 1995-01-31
-- Created by: Mister rmi
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

--Modified by   rob 11-mar-98 : Implement virtual methods from Graphic3d_Structure
--                              to optimize HLR Display...

class Prs from PrsMgr inherits Presentation from Prs3d

uses
    Array2OfReal          from TColStd,
    StructureManager      from Graphic3d,
    Structure             from Graphic3d,
    DataStructureManager  from Graphic3d,
    TypeOfPresentation3d  from PrsMgr,
    PresentationPointer   from PrsMgr
    
is
    Create (theStructManager        : StructureManager from Graphic3d;
            thePresentation         : PresentationPointer from PrsMgr;
            theTypeOfPresentation3d : TypeOfPresentation3d from PrsMgr)
    returns Prs from PrsMgr;

    Compute (me: mutable)
    is redefined static;

    Compute(me : mutable; aProjector: DataStructureManager from Graphic3d)
    returns Structure from Graphic3d
    is redefined static;

    Compute ( me	: mutable;
	      aProjector: DataStructureManager from Graphic3d;
	      AMatrix	: Array2OfReal from TColStd )
    returns Structure from Graphic3d is 
    redefined static;
    ---Purpose: the "degenerated" Structure is displayed with
    --          a transformation defined by <AMatrix>
    --          which is not a Pure Translation.
    --          We have to take in account this Transformation
    --          in the computation of hidden line removal...
    --          returns a filled Graphic Structure.



    Compute(me              : mutable; 
    	    aProjector      : DataStructureManager from Graphic3d;
	    ComputedStruct  : in out Structure from Graphic3d)
    is redefined static;
    ---Purpose: No need to return a structure, just to fill
    --          <ComputedStruct> ....


    Compute ( me	: mutable;
	      aProjector: DataStructureManager from Graphic3d;
	      AMatrix	: Array2OfReal from TColStd ;
    	      aStructure: in out Structure from Graphic3d )
    is redefined static;
    ---Purpose: No Need to return a Structure, just to
    --          Fill <aStructure>. The Trsf has to be taken in account
    --          in the computation (Rotation Part....)

    

fields 
    myPresentation3d: PresentationPointer from PrsMgr;
end Prs from PrsMgr;
