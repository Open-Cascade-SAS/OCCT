-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ApprovalPersonOrganization from StepBasic 

inherits TShared from MMgt

uses

	PersonOrganizationSelect from StepBasic, 
	Approval from StepBasic, 
	ApprovalRole from StepBasic
is

	Create returns ApprovalPersonOrganization;
	---Purpose: Returns a ApprovalPersonOrganization

	Init (me : mutable;
	      aPersonOrganization : PersonOrganizationSelect from StepBasic;
	      aAuthorizedApproval : Approval from StepBasic;
	      aRole : ApprovalRole from StepBasic) is virtual;

	-- Specific Methods for Field Data Access --

	SetPersonOrganization(me : mutable; aPersonOrganization : PersonOrganizationSelect);
	PersonOrganization (me) returns PersonOrganizationSelect;
	SetAuthorizedApproval(me : mutable; aAuthorizedApproval : Approval);
	AuthorizedApproval (me) returns Approval;
	SetRole(me : mutable; aRole : ApprovalRole);
	Role (me) returns ApprovalRole;

fields

	personOrganization : PersonOrganizationSelect from StepBasic; -- a SelectType
	authorizedApproval : Approval from StepBasic;
	role : ApprovalRole from StepBasic;

end ApprovalPersonOrganization;
