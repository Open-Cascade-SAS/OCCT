-- Created on: 1995-01-26
-- Created by: Mister rmi
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class SensitiveSegment from Select2D 
inherits SensitiveEntity from Select2D


	---Purpose: A framework to define sensitive areas along a line segment.

uses
    Pnt2d from gp,
    EntityOwner from SelectBasics,
    ListOfBox2d from SelectBasics    

is


    Create (OwnerId      : EntityOwner from SelectBasics;
    	    FirstP,LastP : Pnt2d from gp;
    	    MaxRect      : Integer = 3)
     returns mutable SensitiveSegment;
    	---Purpose: Constructs the sensitive line segment object defined
    	-- by the owner OwnerId, the 2D starting and ending
    	-- points FirstPoint and LastPoint and the maximum
    	-- number of sensitive bounding boxes MaxRect.
    	-- The parameters can be modified using the functions provided.	    
	    
    Set (me:mutable; MaxRect : Integer) is static;
    	---Purpose: Sets the maximum number of 2D sensitive bounding boxes - MaxRect.
    
    
    
    StartPoint (me : mutable ; aPt : Pnt2d from gp) is static;
    	---Level: Public 
    	---C++: inline
    	---Purpose: changes the start Point of the Segment;
    


    EndPoint (me : mutable ; aPt : Pnt2d from gp) is static;
    	---Level: Public 
    	---C++: inline
    	---Purpose: changes the end point of the segment
    
    
    StartPoint (me) returns Pnt2d from gp;
    	---Level: Public 
    	---Purpose: gives the 3D start Point of the Segment
    	---C++: return const&
    	---C++: inline
    
    
    EndPoint(me) returns Pnt2d from gp;
    	---Level: Public 
    	---Purpose: Returnes the 3D start Point of the Segment
    	---C++: return const&
    	---C++: inline
    
    
    Areas   (me:mutable;aSeq : in out ListOfBox2d from SelectBasics) is static;
    
    
    Matches (me   : mutable; 
    	     X,Y  : Real from Standard;
    	     aTol : Real from Standard;
    	     DMin : out Real from Standard)
    returns Boolean is static;

    Matches (me  :mutable; 
             XMin,YMin,XMax,YMax : Real from Standard;
             aTol: Real from Standard) 
    returns Boolean
    is static;
    

    MaxBoxes(me) returns Integer is redefined static;
    	---Level: Public 
    	---Purpose: Returns the max number of sensitive aeas describing the sensitive segment
    	---C++: inline

fields

    mymaxrect : Integer;
    mystart   : Pnt2d from gp;
    myend     : Pnt2d from gp;

end SensitiveSegment;
