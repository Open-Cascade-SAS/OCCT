-- Created on: 1995-01-31
-- Created by: Dieter THIEMANN
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ActorWrite from STEPControl
    inherits ActorOfFinderProcess  from Transfer
    
    ---Purpose : This class performs the transfer of a Shape from TopoDS
    --           to AP203 or AP214 (CD2 or DIS)


uses FinderProcess, TransientProcess, Binder, Finder, StepModel from StepData,
     Shape from TopoDS,
     StepModelType from STEPControl,
     Axis2Placement3d from StepGeom,
     ShapeRepresentation from StepShape,
     ShapeDefinitionRepresentation from StepShape,
     HAsciiString from TCollection,
     ContextTool from STEPConstruct,
     Part from STEPConstruct,
     HSequenceOfShape from TopTools, -- For non-manifold topology processing (ssv; 13.11.2010)
     NonManifoldSurfaceShapeRepresentation from StepShape -- For non-manifold topology processing (ssv; 13.11.2010)

is

    Create  returns mutable ActorWrite from STEPControl;

    Recognize (me : mutable; start : Finder) returns Boolean  is redefined;

    Transfer (me : mutable; start : Finder; FP : mutable FinderProcess)
    	returns mutable Binder is redefined;
    -- enchains : TransferShape , MakeProductData , and manages mode
    --   "simple" or in Assembly

    TransferSubShape (me : mutable; start : Finder;
                     SDR : ShapeDefinitionRepresentation from StepShape;
                     AX1 : out Axis2Placement3d from StepGeom;
                      FP : mutable FinderProcess;
              shapeGroup : HSequenceOfShape from TopTools = NULL;
              isManifold : Boolean = Standard_True)
    	returns mutable Binder;

    TransferShape (me : mutable; start : Finder;
                  SDR : ShapeDefinitionRepresentation from StepShape;
    	    	       FP : mutable FinderProcess;
		       shapeGroup : HSequenceOfShape from TopTools = NULL;
		       isManifold : Boolean = Standard_True)		      
    	returns mutable Binder;

    TransferCompound (me : mutable; start : Finder;
	              SDR : ShapeDefinitionRepresentation from StepShape;
    	    	      FP : mutable FinderProcess)
    	returns mutable Binder;

--    InitProductData  (me: mutable) returns Part from STEPConstruct;

--    MakeProductData  (me : mutable;
--        SR      : ShapeRepresentation from StepShape;
--    	SDRTool : Part from STEPConstruct;
--	model   : StepModel from StepData;
--        addPRPC : Boolean)
--    	    returns mutable Binder;


    SetMode (me : mutable; M : StepModelType from STEPControl);	

    Mode (me) returns StepModelType from STEPControl;

    SetGroupMode (me : mutable; mode : Integer);
    -- Default is 0 (no group item)
    -- 1 for REPRESENTATION_RELATIONSHIP with ITEM_DEFINED_TRANSFORMATION
    -- other positive values if needed (not implemented)

    GroupMode (me) returns Integer;

    SetTolerance (me : mutable; Tol : Real);
    --  Tol <= 0 means Unset

    IsAssembly (me; S: in out Shape from TopoDS) returns Boolean is virtual;
    	---Purpose: Customizable method to check whether shape S should
	--          be written as assembly or not
	--          Default implementation uses flag GroupMode and analyses
	--          the shape itself
	--          NOTE: this method can modify shape
	
    getNMSSRForGroup (me; 
                      shapeGroup : HSequenceOfShape from TopTools;
                      FP : mutable FinderProcess;
                      isNMSSRCreated : in out Boolean)
    returns NonManifoldSurfaceShapeRepresentation from StepShape
    is private;
    ---Purpose: Non-manifold shapes are stored in NMSSR group
    --          (NON_MANIFOLD_SURFACE_SHAPE_REPRESENTATION).
    --          Use this method to get the corresponding NMSSR (or
    --          to create a new one if doesn't exist yet)
    --          (ssv; 13.11.2010)

fields

    mygroup  :  Integer;
    mytoler  :  Real;
    myContext:  ContextTool from STEPConstruct;
    
end ActorWrite;
