-- Created on: 1992-12-15
-- Created by: Jean Louis FRENKEL
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



generic class CurvePresentation from Prs3d 
    	           ( anyCurve as any; 
    	             CurveTool as any) -- as CurveTool from Adaptor3d

inherits Root from Prs3d

uses
    Presentation from Prs3d,
    Drawer from Prs3d,
    Length from Quantity

is

    --- Purpose:
    --  

    Add(myclass; aPresentation: Presentation from Prs3d; 
    	    	 aCurve: anyCurve;
    	    	 aDrawer: Drawer from Prs3d);

    Add(myclass; aPresentation: Presentation from Prs3d; 
    	    	 aCurve: anyCurve;
                 U1,U2 : Real from Standard;
    	    	 aDrawer: Drawer from Prs3d);

    Add(myclass; aPresentation: Presentation from Prs3d; 
    	    	 aCurve: anyCurve;
    	    	 aDeflection: Real from Standard);

    Add(myclass; aPresentation: Presentation from Prs3d; 
    	    	 aCurve: anyCurve;
                 U1,U2 : Real from Standard;
    	    	 aDeflection: Real from Standard);

		 
    Match(myclass; X,Y,Z: Length from Quantity;
                   aDistance: Length from Quantity;
    	    	   aCurve: anyCurve;
    	    	   aDrawer: Drawer from Prs3d) 
    returns Boolean from Standard;

    Match(myclass; X,Y,Z: Length from Quantity;
                   aDistance: Length from Quantity;
    	    	   aCurve: anyCurve;
                   U1,U2 : Real from Standard;
    	    	   aDrawer: Drawer from Prs3d)
    returns Boolean from Standard;

    Match(myclass; X,Y,Z: Length from Quantity;
                   aDistance: Length from Quantity;
    	    	   aCurve: anyCurve;
    	    	   aDeflection: Real from Standard)
    returns Boolean from Standard;

    Match(myclass; X,Y,Z: Length from Quantity;
                   aDistance: Length from Quantity;
        	   aCurve: anyCurve;
                   U1,U2 : Real from Standard;
    	    	   aDeflection: Real from Standard)
    returns Boolean from Standard;

		 
end CurvePresentation from Prs3d;



