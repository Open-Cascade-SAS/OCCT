-- Created on: 2000-11-16
-- Created by: Peter KURNEV
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Tools from BOPTools 

	---Purpose:  
	---  The class contains handy static functions 
	---  dealing with the topology 
	 
uses 
    Pnt  from  gp ,  
    	
    Shape   from  TopoDS, 
    Vertex  from  TopoDS, 
    Edge    from  TopoDS, 
    Face    from  TopoDS,

    Range   from IntTools, 
    Context from IntTools, 
    Curve   from IntTools, 

    PaveBlock from BOPTools, 
     
    IndexedMapOfShape from TopTools 

is  
    
    
	 
    MakeNewVertex  (myclass;  
        	    aP1 : Pnt  from  gp;  
		    aTol: Real from Standard;
		    aNewVertex:out Vertex from TopoDS); 
    	---Purpose: 
    	--- Make a vertex using 3D-point <aP1> and 3D-tolerance value <aTol>  
    	---
    MakeNewVertex  (myclass;  
        	    aV1,aV2:   Vertex from TopoDS; 
		    aNewVertex:out Vertex from TopoDS); 						 
    	---Purpose: 
    	--- Make a vertex using couple of vertices  <aV1, aV2>     
    	---
    MakeNewVertex  (myclass;  
        	    aE1: Edge from TopoDS; 
		    aP1: Real from Standard; 
    	    	    aE2: Edge from TopoDS; 
		    aP2: Real from Standard; 
    	    	    aNewVertex:out Vertex from TopoDS); 	    			 
    	---Purpose: 
    	--- Make a vertex in place of intersection between two edges 
    	--- <aE1, aE2> with parameters <aP1, aP2>     
    	---
    MakeNewVertex  (myclass;  
        	    aE1: Edge from TopoDS; 
		    aP1: Real from Standard; 
    	    	    aF2: Face from TopoDS; 
    	    	    aNewVertex:out Vertex from TopoDS); 	
    	---Purpose: 
    	--- Make a vertex in place of intersection between the edge <aE1> 
    	--- with parameter <aP1> and the face <aF2> 
    	---
    PointOnEdge    (myclass;   
    	    	    aEdge: Edge from TopoDS; 
		    aPrm: Real from Standard; 
    	    	    aP:out Pnt  from  gp);
    	---Purpose: 
    	--- Compute a 3D-point on the edge <aEdge> at parameter <aPrm> 
    	---
    MakeSplitEdge  (myclass;  
        	    aE1: Edge from TopoDS; 
		    aV1: Vertex from TopoDS;	     
   	    	    aP1: Real from Standard; 
    	    	    aV2: Vertex from TopoDS; 
		    aP2: Real from Standard; 
    	    	    aNewEdge:out Edge from TopoDS); 	 
    	---Purpose: 
    	--- Make the edge from base edge <aE1> and two vertices <aV1,aV2>  
    	--- at parameters <aP1,aP2>  
    	---
    MakeSectEdge   (myclass;  
        	    aIC: Curve  from IntTools; 
		    aV1: Vertex from TopoDS;	     
   	    	    aP1: Real from Standard; 
    	    	    aV2: Vertex from TopoDS; 
		    aP2: Real from Standard; 
    	    	    aNewEdge:out Edge from TopoDS); 	    
    	---Purpose: 
    	--- Make the edge from 3D-Curve <aIC>  and two vertices <aV1,aV2>  
    	--- at parameters <aP1,aP2>  
    	---
    UpdateVertex   (myclass;  
        	    aIC: Curve  from IntTools; 
    	    	    aT : Real from Standard;  
		    aV : Vertex from TopoDS); 
    	---Purpose:   
    	--- Update the tolerance value for vertex  <aV> 
    	--- taking into account the fact that <aV> lays on   
    	--- the curve <aIC>   
    	---
    UpdateVertex   (myclass;  
        	    aE : Edge from TopoDS;  
    	    	    aT : Real from Standard;  
		    aV : Vertex from TopoDS); 	     
    	---Purpose:  
    	--- Update the tolerance value for vertex  <aV> 
    	--- taking into account the fact that <aV> lays on   
    	--- the edge <aE>   
    	---
    UpdateVertex   (myclass;  
    	    	    aVF : Vertex from TopoDS; 
		    aVN : Vertex from TopoDS); 	
    	---Purpose:  
    	--- Update the tolerance value for vertex  <aVN> 
    	--- taking into account the fact that <aVN> should   
    	--- cover tolerance zone of <aVF>    
    	---
    IsBlocksCoinside(myclass;   
    	    	     aPB1: PaveBlock from BOPTools; 
		     aPB2: PaveBlock from BOPTools) 
    	    returns Boolean from Standard;         
    	---Purpose:  
    	--- Returns TRUE if PaveBlocks  <aPB1>,<aPB2> coinside in 3D       
    	--- taking into account corresp. tolerances' values of vertices, 
    	--- edges     
    	---
    IsBlockInOnFace(myclass;   
    	    	     aPB : PaveBlock from BOPTools; 
		     aF  : Face from TopoDS;  
    	    	     aContext: Context from IntTools)  
    	    returns Boolean from Standard;  	     
    	---Purpose:  
    	--- Returns TRUE if PaveBlock <aPB> lays on the face <aF>, i.e 
    	--- the <PB> is IN or ON in 2D of <aF>               
    	---
    MapShapes      (myclass; 
		     aS : Shape from TopoDS; 
		     aM :out IndexedMapOfShape from TopTools); 		      
    	---Purpose:  
    	--- Get a  Map <aM> containing the shape itself and all its subshapes   
    	---
    CorrectRange   (myclass;  
    	    	     aE1:   Edge from TopoDS;    
    	    	     aE2:   Edge from TopoDS;   
		     aSR:   Range from IntTools;  		      
		     aNewSR:out  Range from IntTools);  
    	---Purpose:  
    	--- Correct shrunk range <aSR> taking into account 3D-curve      
    	--- resolution and corresp. tolerances' values of <aE1>, <aE2>   
    	---
    CorrectRange   (myclass;  
    	    	     aE:   Edge from TopoDS;    
    	    	     aF:   Face from TopoDS;   
		     aSR:  Range from IntTools;  		      
		     aNewSR:out  Range from IntTools); 
    	---Purpose:  
    	--- Correct shrunk range <aSR> taking into account 3D-curve      
    	--- resolution and corresp. tolerances' values of <aE>, <aF>
    	---
    CopySource (myclass;  
    	    	    aSourceShape:  Shape from TopoDS;   
       	    	    aDestShape:out Shape from TopoDS);  
    	---Purpose: 
    	--- Make a copy of <aSourceShape> 
	---
     
end Tools;
