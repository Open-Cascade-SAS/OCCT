-- Created on: 1995-02-22
-- Created by: Mister rmi
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

--Modified by Rob Jan 13 th  98 : Compute Depth on EyeLine for
--                                Each Kind of SensitiveEntity. 
--                                (Deferred Method to be implemented)


package Select3D 

	---Purpose: The Select3D package provides the following services
    	-- -   definition of standard   3D sensitive primitives such as points, curves and faces.
    	-- -   recovery of the bounding boxes in the 2D graphic selection space, if required.
    	-- -   a 3D-2D projector.

uses
    Standard,
    TCollection,
    TColStd,
    TColgp,
    gp,
    Bnd,
    Poly,
    TopLoc,
    Geom,
    SelectBasics,
    SelectMgr,
    V3d,
    Graphic3d

is

    imported BndBox3d;
    imported BVHPrimitiveContent;
    imported InteriorSensitivePointSet;
    imported EntitySequence;
    imported Pnt;
    imported PointData;
    imported SelectingVolumeManager;
    imported SensitiveBox;
    imported SensitiveCircle;
    imported SensitiveCurve;
    imported transient class SensitiveEntity;
    imported SensitiveFace;
    imported SensitiveGroup;
    imported SensitivePoint;
    imported SensitivePoly;
    imported SensitiveSegment;
    imported SensitiveSet;
    imported SensitiveTriangle;
    imported SensitiveTriangulation;
    imported SensitiveWire;
    imported TypeOfSensitivity;

end Select3D;
