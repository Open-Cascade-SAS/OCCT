-- Created on: 1997-12-10
-- Created by: Denis PASCAL
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Variable from PDataStd inherits Attribute from PDF

	---Purpose: Persistant variable
	--          ===================

uses HAsciiString from PCollection
is

    Create returns mutable Variable from PDataStd;

    
    Create (constant : Boolean from Standard)
    returns mutable Variable from PDataStd;
    
    Constant (me : mutable; status : Boolean from Standard);    
    Constant (me)
    returns Boolean from Standard;

    Unit(me:mutable; unit : HAsciiString from PCollection);
    Unit(me) 
    returns HAsciiString from PCollection;

fields

    isConstant : Boolean      from Standard;
    myUnit     : HAsciiString from PCollection;

end Variable;
