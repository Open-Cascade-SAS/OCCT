-- Created on: 1999-11-26
-- Created by: Andrey BETENEV
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0

class VersionedActionRequest from StepBasic
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity VersionedActionRequest

uses
    HAsciiString from TCollection

is
    Create returns VersionedActionRequest from StepBasic;
	---Purpose: Empty constructor

    Init (me: mutable; aId: HAsciiString from TCollection;
                       aVersion: HAsciiString from TCollection;
                       aPurpose: HAsciiString from TCollection;
                       hasDescription: Boolean;
                       aDescription: HAsciiString from TCollection);
	---Purpose: Initialize all fields (own and inherited)

    Id (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Id
    SetId (me: mutable; Id: HAsciiString from TCollection);
	---Purpose: Set field Id

    Version (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Version
    SetVersion (me: mutable; Version: HAsciiString from TCollection);
	---Purpose: Set field Version

    Purpose (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Purpose
    SetPurpose (me: mutable; Purpose: HAsciiString from TCollection);
	---Purpose: Set field Purpose

    Description (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Description
    SetDescription (me: mutable; Description: HAsciiString from TCollection);
	---Purpose: Set field Description
    HasDescription (me) returns Boolean;
	---Purpose: Returns True if optional field Description is defined

fields
    theId: HAsciiString from TCollection;
    theVersion: HAsciiString from TCollection;
    thePurpose: HAsciiString from TCollection;
    theDescription: HAsciiString from TCollection; -- optional
    defDescription: Boolean; -- flag "is Description defined"

end VersionedActionRequest;
