-- Created on: 1993-01-12
-- Created by: Philippe DAUTRY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package BRepSweep

    ---Purpose: This package implements the package Sweep for the BRep
    --          structure.

uses

    Standard,
    Quantity,
    TCollection, 
    TColStd,
    gp, 
    Geom,
    TopAbs, 
    TopLoc, 
    TopTools, 
    TopoDS, 
    TopExp, 
    BRep,
    Sweep

is

    class Builder;
	---Purpose: Implements the Builder required for Sweep.

    class Tool;
	---Purpose: Provides an indexation of the subShapes of a Shape
	--          from TopoDS.
	
    class Iterator;
	---Purpose: Iterator on the subShapes of a shape.
	

    deferred class NumLinearRegularSweep
    	instantiates LinearRegularSweep from Sweep(
    	Shape              from TopoDS,     -- Resulting topological objects.
    	Shape              from TopoDS,     -- Generating Shape.
    	NumShape           from Sweep,      -- Directing Wire.
    	Builder            from BRepSweep,
    	Tool               from BRepSweep,  -- GenTool
	NumShapeTool       from Sweep,      -- DirTool
    	Iterator           from BRepSweep,  -- Resulting objects Iterator
    	Iterator           from BRepSweep,  -- GenIterator
	NumShapeIterator   from Sweep);     -- DirSubEdgeIterator

    deferred class Trsf;
    --- This class is inherited  from LinearRegularSweep to  implement
    --  the simple swept primitives built moving a Shape with a Trsf.

    class Translation;
    --- This class is inherited from Trsf to implement the translation
    --  sweep.

    class Rotation;
    --- This class is  inherited  from Trsf to implement  the rotation
    --  sweep.

    class Prism;
    --- This class provides simple methods to build prism.

    class Revol;
    --- This class provides simple methods to build Revol.

end BRepSweep;
