-- Created on: 2001-05-08
-- Created by: Peter KURNEV
-- Copyright (c) 2001-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Curve from BOPTools 

	---Purpose:  
    	--  Class holds the  structure for storing information about  
    	--- intersection curve and set of paves on it     
    	---     

uses 
    ListOfInteger from  TColStd,  
    Curve           from IntTools, 
    PaveSet         from BOPTools, 
    PaveBlock       from BOPTools, 
    ListOfPaveBlock from BOPTools 
    

is
    Create   
    	returns Curve from BOPTools; 
    	---Purpose:  
    	--- Empty constructor 
    	---
    Create  (aIC:Curve from IntTools) 
    	returns Curve from BOPTools; 
    	---Purpose:  
    	--- Constructor 
    	---
    SetCurve(me:out; 
    	     aIC:Curve from IntTools); 
    	---Purpose:  
    	--- Modifier 
    	---
    Curve(me)
    	returns Curve from IntTools; 
    	---C++:  return const &  
    	---Purpose:  
    	--- Selector 
    	---
    Set(me:out) 
    	returns PaveSet from BOPTools; 
    	---C++:  return &  
    	---Purpose:  
    	--- Selector 
    	--- 
    AppendNewBlock(me:out;   
    	    	aPB:PaveBlock from BOPTools);      
    	---Purpose:  
    	--- Adds the PaveBlock  <aPB> to the pave set    
    	---
    NewPaveBlocks(me) 
    	returns ListOfPaveBlock from BOPTools; 
    	---C++:  return const & 
    	---Purpose:  
    	--- Returns the PaveBlock-s attached to the curve      
    	---
    TechnoVertices (me:out) 
    	returns ListOfInteger from TColStd; 
    	---C++:  return &  
    	---Purpose:  
    	--- Returns indices TechnoVertices attached to the curve      
    	---

fields
    myCurve  : Curve           from IntTools;
    myPaveSet: PaveSet         from BOPTools;
    myNewPBs : ListOfPaveBlock from BOPTools;   
    myTechnoVertices    : ListOfInteger from  TColStd; 

end Curve;
