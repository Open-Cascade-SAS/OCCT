-- Created on: 1999-12-08
-- Created by: Vladislav ROMASHKO
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package QANewDBRepNaming

    ---Purpose: To test topological naming

uses 
 
    Draw,
    TCollection, 
    TDF,
    TNaming,
    TopoDS,
    gp

is

    AllCommands       (Di : in out Interpretor from Draw);

    PrimitiveCommands (DI : in out Interpretor from Draw);
--    OffsetCommands    (DI : in out Interpretor from Draw);
--    FilletCommands    (DI : in out Interpretor from Draw);
    FeatureCommands   (DI : in out Interpretor from Draw);
    
end QADBRepNaming;
