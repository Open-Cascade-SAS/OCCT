-- Created on: 2004-09-03
-- Created by: Oleg FEDYAEV
-- Copyright (c) 2004-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ArgumentAnalyzer from BOPAlgo
  inherits Algo from BOPAlgo
    ---Purpose: check the validity of argument(s) for Boolean Operations
    
uses
    Shape       from TopoDS,
    Operation   from BOPAlgo, 
    CheckStatus from BOPAlgo,
    ShapeEnum  from TopAbs,
    ListOfCheckResult  from BOPAlgo,
    DataMapOfShapeReal from BOPCol
    
is
    Create
       returns ArgumentAnalyzer;
    ---C++: alias "Standard_EXPORT virtual ~BOPAlgo_ArgumentAnalyzer();"
    ---Purpose: empty constructor

    SetShape1(me: in out; TheShape: Shape from TopoDS);
    ---Purpose: sets object shape

    SetShape2(me: in out; TheShape: Shape from TopoDS);
    ---Purpose: sets tool shape

    GetShape1(me)
    returns Shape from TopoDS;
    ---C++: return const &
    ---Purpose: returns object shape;

    GetShape2(me)
    returns Shape from TopoDS;
    ---C++: return const &
    ---Purpose: returns tool shape

    ---options
    OperationType(me: in out)
    returns Operation from BOPAlgo;
    ---C++: return &
    ---Purpose: returns ref

    StopOnFirstFaulty(me: in out)
    returns Boolean from Standard;
    ---C++: return &
    ---Purpose: returns ref

    ArgumentTypeMode(me: in out)
    returns Boolean from Standard;
    ---C++: return &
    ---C++: inline
    ---Purpose: Returns (modifiable) mode 
    --          that means checking types of shapes. 
     
    Prepare(me: in out) 
    is protected; 
    ---Purpose: Prepares data;

    SelfInterMode(me: in out)
    returns Boolean from Standard;
    ---C++: return &
    ---C++: inline
    ---Purpose: Returns (modifiable) mode that means
    --          checking of self-intersection of shapes.

    SmallEdgeMode(me: in out)
    returns Boolean from Standard;
    ---C++: return &
    ---C++: inline
    ---Purpose: Returns (modifiable) mode that means
    --          checking of small edges.

    RebuildFaceMode(me: in out)
    returns Boolean from Standard;
    ---C++: return &
    ---C++: inline
    ---Purpose: Returns (modifiable) mode that means
    --          checking of possibility to split or rebuild faces.

    TangentMode(me: in out)
    returns Boolean from Standard;
    ---C++: return &
    ---C++: inline
    ---Purpose: Returns (modifiable) mode that means
    --          checking of tangency between subshapes.

    MergeVertexMode(me: in out)
    returns Boolean from Standard;
    ---C++: return &
    ---C++: inline
    ---Purpose: Returns (modifiable) mode that means
    --          checking of problem of merging vertices.
 
    MergeEdgeMode(me: in out)
    returns Boolean from Standard;
    ---C++: return &
    ---C++: inline
    ---Purpose: Returns (modifiable) mode that means
    --          checking of problem of merging edges.

    ContinuityMode(me: in out)
    returns Boolean from Standard;
    ---C++: return &
    ---C++: inline
    ---Purpose: Returns (modifiable) mode that means
    --          checking of problem of continuity of the shape.

    CurveOnSurfaceMode(me: in out) 
    returns Boolean from Standard;
    ---C++: return &
    ---C++: inline
    ---Purpose: Returns (modifiable) mode that means
    --          checking of problem of invalid curve on surface.

    ---
    Perform(me: out);
    ---Purpose: performs analysis

    HasFaulty(me)
    returns Boolean from Standard;
    ---Purpose: result of test

    GetCheckResult(me)
    returns ListOfCheckResult from BOPAlgo;
    ---C++: return const &
    ---Purpose: returns a result of test

    --- protected	
    TestTypes(me: out)
    is protected;

    TestSelfInterferences(me: out)
    is protected;

    TestSmallEdge(me: out)
    is protected;

    TestRebuildFace(me: out)
    is protected;

    TestTangent(me: out)
    is protected;

    TestMergeSubShapes(me: out; theType: ShapeEnum from TopAbs)
    is protected;

    TestMergeVertex(me: out)
    is protected;

    TestMergeEdge(me: out)
    is protected;

    TestContinuity(me: out)
    is protected; 
     
    TestCurveOnSurface(me: out) 
    is protected;

--  TestMergeFace(me: out)
--  is protected;  

    SetFuzzyValue(me:out; 
      theFuzz : Real from Standard);
    ---C++: inline
    ---Purpose: Sets the additional tolerance

    FuzzyValue(me)
    returns Real from Standard;
    ---C++: inline
    ---Purpose: Returns the additional tolerance 

    UpdateTolerances(me:out)
    is protected; 
    ---Purpose: Updates the shapes tolerance values.

    SetDefaultTolerances(me:out)
    is protected; 
    ---Purpose: Reverts the tolerance values for all entities to default values.

fields

    myShape1             : Shape     from TopoDS;
    myShape2             : Shape     from TopoDS;
    myStopOnFirst        : Boolean   from Standard;
    myOperation          : Operation from BOPAlgo;
    myArgumentTypeMode   : Boolean   from Standard;
    mySelfInterMode      : Boolean   from Standard;
    mySmallEdgeMode      : Boolean   from Standard;
    myRebuildFaceMode    : Boolean   from Standard;
    myTangentMode        : Boolean   from Standard;
    myMergeVertexMode    : Boolean   from Standard;
    myMergeEdgeMode      : Boolean   from Standard;
    myContinuityMode     : Boolean   from Standard; 
    myCurveOnSurfaceMode : Boolean   from Standard; 
    myEmpty1, myEmpty2   : Boolean   from Standard; 
    myResult             : ListOfCheckResult from BOPAlgo;
    myFuzzyValue         : Real      from Standard;
    myToleranceMap       : DataMapOfShapeReal from BOPCol;

end ArgumentAnalyzer;
