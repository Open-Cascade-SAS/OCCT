-- Created on: 1993-03-02
-- Created by: Philippe DAUTRY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class OffsetSurface from PGeom inherits Surface from PGeom

        ---Purpose : This class implements  the basis services for  an
        --         offset surface in 3D space.
        --         

uses Surface from PGeom

is


  Create returns mutable OffsetSurface from PGeom;
    ---Purpose: Creates an OffsetSurface with default values.
    	---Level: Internal 


  Create (
    	    aBasisSurface : Surface from PGeom;
    	    aOffsetValue : Real from Standard)
     returns mutable OffsetSurface from PGeom;
        ---Purpose :  <aBasisSurface>    is  the   basis      surface,
        --         <aOffsetValue> is the distance between <me> and the
        --         basis  surface at any  point.    <aOffsetDirection>
        --         defines  the  fixed  reference  direction   (offset
        --         direction).
    	---Level: Internal 


  BasisSurface (me : mutable; aBasisSurface : Surface from PGeom);
	---Purpose: Set the field basisSurface with <aBasisSurface>.
    	---Level: Internal 
      

  BasisSurface (me) returns Surface from PGeom;
        ---Purpose : The basis surface can be an offset surface.
    	---Level: Internal 


  OffsetValue (me : mutable; aOffsetValue : Real from Standard);
        ---Purpose : Set the field offsetValue with <aOffsetValue>.
    	---Level: Internal 


  OffsetValue (me) returns Real from Standard;
        ---Purpose : Returns the value of the field offsetValue.
    	---Level: Internal 


fields

  basisSurface : Surface from PGeom;
  offsetValue  : Real from Standard;

end;
