-- Created on: 1996-01-29
-- Created by: Christian CAILLET
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class SignType  from IFSelect  inherits Signature

    ---Purpose : This Signature returns the cdl Type of an entity, under two
    --           forms :
    --           - complete dynamic type (package and class)
    --           - class type, without package name

uses CString, Transient, InterfaceModel

is

    Create (nopk : Boolean = Standard_False) returns mutable SignType;
    ---Purpose : Returns a SignType
    --           <nopk> false (D) : complete dynamic type (name = Dynamic Type)
    --           <nopk> true : class type without pk (name = Class Type)

    Value (me; ent : any Transient; model : InterfaceModel) returns CString;
    ---Purpose : Returns the Signature for a Transient object, as its Dynamic
    --           Type, with or without package name, according starting option

fields

    thenopk : Boolean;

end SignType;
