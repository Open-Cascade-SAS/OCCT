-- Created on: 2001-03-06
-- Created by: Christian CAILLET
-- Copyright (c) 2001-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class SignColor  from IGESSelect    inherits Signature  from IFSelect

    ---Purpose : Gives Color attached to an entity
    --           Several forms are possible, according to <mode>
    --           1 : number : "Dnn" for entity, "Snn" for standard, "(none)" for 0
    --           2 : name : Of standard color, or of the color entity, or "(none)"
    --               (if the color entity has no name, its label is taken)
    --           3 : RGB values, form R:nn,G:nn,B:nn
    --           4 : RED value   : an integer
    --           5 : GREEN value : an integer
    --           6 : BLUE value  : an integer
    --           Other computable values can be added if needed :
    --           CMY values, Percentages for Hue, Lightness, Saturation

uses CString, Transient, AsciiString, InterfaceModel

is

    Create (mode : Integer) returns SignColor;
    ---Purpose : Creates a SignColor
    --           mode : see above for the meaning
    --           modes 4,5,6 give a numeric integer value
    --           Name is initialised according to the mode

    Value   (me; ent : any Transient; model : InterfaceModel) returns CString;
    ---Purpose : Returns the value (see above)

fields

    themode : Integer;

end SignColor;
