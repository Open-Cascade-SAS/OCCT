-- Created on: 1995-03-17
-- Created by: Mister rmi
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Modification: DCB 14-07-98
--    SetColorIndices() method has been added to avoid exception
--    after V2d_Viewer::SetColorMap() call.

private class CircularGrid from V2d inherits CircularGrid from Aspect

uses
    ViewerPointer from V2d,
    View from V2d,
    GraphicObject from Graphic2d,
    CircularGraphicGrid from V2d,
    NameOfColor from Quantity
is
    Create(aViewer: ViewerPointer from V2d;
           aColorIndex1: Integer from Standard;
           aColorIndex2: Integer from Standard)
    returns mutable CircularGrid from V2d;

    SetColorIndices (me: mutable;
                     aColorIndex1: Integer from Standard;
                     aColorIndex2: Integer from Standard);

    Display(me: mutable)
    is redefined static;

    Erase(me)
    is redefined static;

    IsDisplayed(me)
    returns Boolean from Standard
    is redefined static;

    UpdateDisplay(me:mutable)
    is redefined static protected;

fields
    myViewer: ViewerPointer from V2d;
    myGraphicObject: GraphicObject from Graphic2d;
    myColorIndex1: Integer from Standard;
    myColorIndex2: Integer from Standard;
    myGrid: CircularGraphicGrid from V2d;

end CircularGrid from V2d;
