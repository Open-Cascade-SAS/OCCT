-- File:	Extrema_GExtCC.cdl
-- Created:	Wed Jul  6 14:37:10 1994
-- Author:	Laurent PAINNOT
--		<lpa@metrox>
---Copyright:	 Matra Datavision 1994


generic class GExtCC from Extrema (Curve1    as any;
    	    	    	    	   Tool1     as any;
    	    	    	    	   Curve2    as any;
    	    	    	    	   Tool2     as any)

	---Purpose: It calculates all the distance between two curves.
	--          These distances can be maximum or minimum.

uses POnCurv           from Extrema,
     SequenceOfPOnCurv from Extrema,
     ExtElC            from Extrema,
     Pnt               from gp,
     HArray1OfPnt      from TColgp,
     SequenceOfReal    from TColStd,
     ListOfTransient   from TColStd


raises  InfiniteSolutions from StdFail,
    	NotDone           from StdFail,
    	OutOfRange        from Standard
	
    class CCache instantiates CurveCache from Extrema (Curve1, Pnt from gp, HArray1OfPnt from TColgp);

    class ECC instantiates GenExtCC from Extrema
        (Curve1,
         Tool1,
         Curve2,
         Tool2,
         CCache,
         HArray1OfPnt from TColgp,
         POnCurv,
         Pnt,
         Vec);


is

    Create (TolC1: Real = 1.0e-10; TolC2: Real = 1.0e-10) returns GExtCC;
    

    Create (C1: Curve1;  C2: Curve2;
            TolC1: Real = 1.0e-10; TolC2: Real = 1.0e-10) returns GExtCC;
      	---Purpose: It calculates all the distances.


    Create (C1: Curve1;
    	    C2: Curve2;
	    U1: Real  from Standard;
	    U2: Real  from Standard;
	    V1: Real  from Standard;
	    V2: Real  from Standard;
            TolC1: Real = 1.0e-10;
            TolC2: Real = 1.0e-10) returns GExtCC;
      	---Purpose: It calculates all the distances.


    SetCurve (me: in out; theRank: Integer; C: Curve1);
        ---Purpose:

    SetCurve (me: in out; theRank: Integer; C: Curve1; Uinf, Usup: Real);
        ---Purpose:

    SetRange (me: in out; theRank: Integer; Uinf, Usup: Real);
        ---Purpose:

    SetTolerance (me: in out; theRank: Integer; Tol: Real);
        ---Purpose:

    Perform(me: in out);
    

    IsDone (me) returns Boolean
    	---Purpose: Returns True if the distances are found.
    	is static;

    NbExt (me) returns Integer
    	---Purpose: Returns the number of extremum distances.
    	raises  NotDone from StdFail,
	    	-- if IsDone(me)=False.
    	    	InfiniteSolutions from StdFail
		-- if IsParallel(me)= True.
    	is static;


    IsParallel (me) returns Boolean
    	---Purpose: Returns True if the two curves are parallel.
    	raises  NotDone from StdFail
	    	-- if IsDone(me)=False.
    	is static;


    SquareDistance (me; N: Integer =1) returns Real
    	---Purpose: Returns the value of the Nth extremum square distance.
    	raises  NotDone from StdFail,
	    	-- if IsDone(me)=False.
    	    	InfiniteSolutions from StdFail,
		-- if IsParallel(me)= True and N > 1.
    	    	OutOfRange
		-- if N < 1 or N > NbExt(me)
    	is static;

    Points (me; N: Integer; P1,P2: out POnCurv)
    	---Purpose: Returns the points of the Nth extremum distance.
    	--          P1 is on the first curve, P2 on the second one.
    	raises  NotDone from StdFail,
	    	-- if IsDone(me)=False.
    	    	InfiniteSolutions from StdFail,
		-- if IsParallel(me)= True.
    	    	OutOfRange
		-- if N < 1 or N > NbExt(me)
    	is static;

    TrimmedSquareDistances(me; dist11, distP12, distP21, distP22: out Real;
                     P11, P12, P21, P22: out Pnt)
    	---Purpose: if the curve is a trimmed curve,
    	--          dist11 is a square distance between the point on C1
    	--          of parameter FirstParameter and the point of 
    	--          parameter FirstParameter on C2.

    is static;
    
    Results(me: in out; AlgExt: ExtElC from Extrema;
    	    Ut11, Ut12, Ut21, Ut22: Real)

    is static protected;    	

    Results(me: in out;AlgExt: ECC;
    	    Ut11, Ut12, Ut21, Ut22: Real)

    is static protected;


    

fields
    myECC:    ECC from Extrema;
    myDone:   Boolean;
    myIsPar:  Boolean;
    mypoints: SequenceOfPOnCurv from Extrema;
    mySqDist: SequenceOfReal    from TColStd;
    mynbext:  Integer;
    inverse:  Boolean;
    myC:     Address from Standard [2];
    myInf: Real [2];
    mySup: Real [2];
    myTol:  Real [2];
    myCacheLists: ListOfTransient from TColStd [2]; -- lists of Handle(Extrema_CCache)
    P1f:      Pnt;
    P1l:      Pnt;
    P2f:      Pnt;
    P2l:      Pnt;
    mydist11: Real;
    mydist12: Real;
    mydist21: Real;
    mydist22: Real;
    


end GExtCC;
