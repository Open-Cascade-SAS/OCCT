-- File:        StepVisual.cdl
-- Created:     Mon Dec  4 12:02:22 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




package RWStepVisual 

uses

	StepData, Interface, TCollection, TColStd, StepVisual

is


--class ReadWriteModule;

--class GeneralModule;

-- Removed from Rev2 to Rev4 : class RWAnnotationCurveOccurrence;
-- Removed from Rev2 to Rev4 : class RWAnnotationFillArea;
-- Removed from Rev2 to Rev4 : class RWAnnotationFillAreaOccurrence;
-- Removed from Rev2 to Rev4 : class RWAnnotationOccurrence;
-- Removed from Rev2 to Rev4 : class RWAnnotationSubfigureOccurrence;
-- Removed from Rev2 to Rev4 : class RWAnnotationSymbol;
-- Removed from Rev2 to Rev4 : class RWAnnotationSymbolOccurrence;
-- Removed from Rev2 to Rev4 : class RWAnnotationText;
-- Removed from Rev2 to Rev4 : class RWAnnotationTextOccurrence;
class RWAreaInSet;
class RWBackgroundColour;
class RWCameraImage;
class RWCameraModel;
class RWCameraModelD2;
class RWCameraModelD3;
class RWCameraUsage;
class RWColour;
class RWColourRgb;
class RWColourSpecification;
class RWContextDependentInvisibility;
class RWContextDependentOverRidingStyledItem;
-- Removed from CC1-Rev2 to CC1-Rev4, re-added CC2-Rev4 :
class RWCompositeText;
-- Removed from Rev2 to Rev4 : class RWCompositeTextWithAssociatedCurves;
-- Removed from Rev2 to Rev4 : class RWCompositeTextWithBlankingBox;
-- Removed from CC1-Rev2 to CC1-Rev4, re-added CC2-Rev4 :
class RWCompositeTextWithExtent;

class RWCurveStyle;
class RWCurveStyleFont;
class RWCurveStyleFontPattern;
-- Removed from Rev2 to Rev4 : class RWDefinedSymbol;
-- Removed from Rev2 to Rev4 : class RWDimensionCurve;
-- Removed from Rev2 to Rev4 : class RWDimensionCurveTerminator;
-- Removed from Rev2 to Rev4 : class RWDraughtingAnnotationOccurrence;
-- Removed from Rev2 to Rev4 : class RWDraughtingCallout;
class RWDraughtingModel; -- added for CAX-IF TR3
class RWDraughtingPreDefinedColour;
class RWDraughtingPreDefinedCurveFont;
-- Removed from Rev2 to Rev4 : class RWDraughtingSubfigureRepresentation;
-- Removed from Rev2 to Rev4 : class RWDraughtingSymbolRepresentation;
-- Removed from Rev2 to Rev4 : class RWDraughtingTextLiteralWithDelineation;
-- Removed from Rev2 to Rev4 : class RWDrawingDefinition;
-- Removed from Rev2 to Rev4 : class RWDrawingRevision;
--moved to RWStepBasic: class RWExternalSource;
class RWExternallyDefinedCurveFont;
-- Removed from Rev2 to Rev4 : class RWExternallyDefinedHatchStyle;
--moved to RWStepBasic: class RWExternallyDefinedItem;
-- Removed from Rev2 to Rev4 : class RWExternallyDefinedSymbol;
-- Removed from Rev2 to Rev4 : class RWExternallyDefinedTextFont;
-- Removed from Rev2 to Rev4 : class RWExternallyDefinedTileStyle;
class RWFillAreaStyle;
class RWFillAreaStyleColour;
-- Removed from Rev2 to Rev4 : class RWFillAreaStyleHatching;
-- Removed from Rev2 to Rev4 : class RWFillAreaStyleTileSymbolWithStyle;
-- Removed from Rev2 to Rev4 : class RWFillAreaStyleTiles;
class RWInvisibility;
class RWMechanicalDesignGeometricPresentationArea;
class RWMechanicalDesignGeometricPresentationRepresentation;
-- Removed from Rev2 to Rev4 : class RWMechanicalDesignPresentationArea;
class RWOverRidingStyledItem;
class RWPlanarBox;
class RWPlanarExtent;
class RWPointStyle;
class RWPreDefinedColour;
class RWPreDefinedCurveFont;
class RWPreDefinedItem;
-- Removed from Rev2 to Rev4 : class RWPreDefinedSymbol;
-- Removed from Rev2 to Rev4 : class RWPreDefinedTextFont;
class RWPresentationArea;
class RWPresentationLayerAssignment;
class RWPresentationRepresentation;
class RWPresentationSet;
class RWPresentationSize;
class RWPresentationStyleAssignment;
class RWPresentationStyleByContext;
class RWPresentationView;
-- Removed from Rev2 to Rev4 : class RWProductDataRepresentationView;
class RWStyledItem;
class RWSurfaceSideStyle;
class RWSurfaceStyleBoundary;
class RWSurfaceStyleControlGrid;
class RWSurfaceStyleFillArea;
class RWSurfaceStyleParameterLine;
class RWSurfaceStyleSegmentationCurve;
class RWSurfaceStyleSilhouette;
class RWSurfaceStyleUsage;
-- Removed from Rev2 to Rev4 : class RWSymbolColour;
-- Removed from Rev2 to Rev4 : class RWSymbolRepresentation;
-- Removed from Rev2 to Rev4 : class RWSymbolRepresentationMap;
-- Removed from Rev2 to Rev4 : class RWSymbolStyle;
-- Removed from Rev2 to Rev4 : class RWSymbolTarget;
class RWTemplate;
class RWTemplateInstance;
-- Removed from Rev2 to Rev4 : class RWTerminatorSymbol;
-- Removed from CC1-Rev2 to CC1-Rev4, re-added CC2-Rev4 :
class RWTextLiteral;
-- Removed from Rev2 to Rev4 : class RWTextLiteralWithAssociatedCurves;
-- Removed from Rev2 to Rev4 : class RWTextLiteralWithBlankingBox;
-- Removed from Rev2 to Rev4 : class RWTextLiteralWithDelineation;
-- Removed from Rev2 to Rev4 : class RWTextLiteralWithExtent;
-- Removed from CC1-Rev2 to CC1-Rev4, re-added CC2-Rev4 :
class RWTextStyle;
class RWTextStyleForDefinedFont;
class RWTextStyleWithBoxCharacteristics;
-- Removed from Rev2 to Rev4 : class RWTextStyleWithMirror;
class RWViewVolume;

    -- Added from Rev2 to Rev4
class RWPresentedItemRepresentation;
class RWPresentationLayerUsage;


	---Package Method ---

--	Init;
	---Purpose: enforced the initialisation of the  libraries

end RWStepVisual;
