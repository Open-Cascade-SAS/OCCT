-- Created on: 2001-09-19
-- Created by: admin of fao FACTORY
-- Copyright (c) 2001-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

private class NamespaceDef from XmlLDrivers

uses    AsciiString from TCollection

is
    Create returns NamespaceDef from XmlLDrivers;
    
    Create (thePrefix: AsciiString from TCollection;
            theURI   : AsciiString from TCollection)
        returns NamespaceDef from XmlLDrivers;

    Prefix (me) returns AsciiString from TCollection;
    ---C++: return const &

    URI (me) returns AsciiString from TCollection;
    ---C++: return const &

fields

    myPrefix :  AsciiString     from TCollection;
    myURI    :  AsciiString     from TCollection;

end NamespaceDef;
