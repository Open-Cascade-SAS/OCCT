-- Created on: 1997-10-08
-- Created by: Olga KOULECHOVA
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


deferred class RibSlot from BRepFeat inherits MakeShape from BRepBuilderAPI

        ---Purpose:  Provides functions to build mechanical features.
            -- Mechanical features include ribs - protrusions and grooves (or slots) - depressions along
            -- planar (linear) surfaces or revolution surfaces. The semantics of mechanical features is built
            -- around giving thickness to a contour. This thickness can either be unilateral - on one side
            -- of the contour - or bilateral - on both sides.
            -- As in the semantics of form features, the thickness is defined by construction of shapes
            -- in specific contexts. The development contexts differ, however,in case of mechanical features.
            -- Here they include extrusion:
            -- -   to a limiting face of the basis shape
            -- -   to or from a limiting plane
            -- -   to a height.

uses Shape                     from TopoDS,
     Face                      from TopoDS,
     Wire                      from TopoDS,
     Edge                      from TopoDS,
     Vertex                    from TopoDS,
     ShapeModification         from BRepBuilderAPI,
     DataMapOfShapeListOfShape from TopTools,
     ListOfShape               from TopTools,
     SequenceOfCurve           from TColGeom,
     Plane                     from Geom,
     Curve                     from Geom,
     DataMapOfShapeShape       from TopTools,
     
     Gluer                     from LocOpe,
     HBuilder                  from TopOpeBRepBuild,
     PerfSelection             from BRepFeat,
     Pnt                       from gp,
     Dir                       from gp,
     StatusError               from BRepFeat,
     --modified by NIZNHY-PKV Thu Mar 21 17:09:08 2002  f 
     BooleanOperation          from BRepAlgoAPI
     --modified by NIZNHY-PKV Thu Mar 21 17:09:11 2002  t
is

    Initialize;
    
        ---Purpose: Redefines the empty constructor.
        ---C++: inline


---  Methods redefined from BRepBuilderAPI_MakeShape

    IsDeleted(me : in out ; F: Shape from TopoDS) 
    returns Boolean from Standard 
    is redefined;
            ---Purpose: Returns true if F a TopoDS_Shape of type edge or face has been deleted.   
    
    Modified(me: in out; F: Shape from TopoDS)
            ---Purpose: Returns the list of generated Faces F. This list may be empty.
            ---C++:     return const &
    returns ListOfShape from TopTools
    is redefined;
    

    Generated(me: in out; S: Shape from TopoDS)
            ---Purpose: Returns a list TopTools_ListOfShape of the faces S created in the shape.
        ---C++:     return const &
    returns ListOfShape from TopTools
    is redefined;


    FirstShape (me)
            ---Purpose: Returns the list  of shapes created  at the bottom  of
            --          the created form.  It may be an empty list.
    returns ListOfShape from TopTools;
             ---C++: return const&


    LastShape (me)
            ---Purpose: Returns  the list of shapes  created at the top of the
            --          created form.  It may be an empty list.
    returns ListOfShape from TopTools;
             ---C++: return const&

    LFPerform(me: in out)
            ---Purpose: General perform method...

            is static protected;

    FacesForDraft(me)
            ---Purpose: Returns a list of the limiting and glueing faces
            -- generated by the feature. These faces did not originally exist in the basis shape.
            -- The list provides the information necessary for
            -- subsequent addition of a draft to a face. It may be an empty list.
            -- If a face has tangent edges, no draft is possible, and the tangent edges must
            -- subsequently be removed if you want to add a draft to the face.
    returns ListOfShape from TopTools;
             ---C++: return const&

    NewEdges(me)
            ---Purpose: Returns a list of the limiting and glueing edges
            -- generated by the feature. These edges did not originally exist in the basis shape.
            -- The list provides the information necessary for
            -- subsequent addition of fillets. It may be an empty list.
    returns ListOfShape from TopTools;
             ---C++: return const&

    TgtEdges(me)
            ---Purpose: Returns a list of the tangent edges among the
            -- limiting and glueing edges generated by the
            -- feature. These edges did not originally exist in
            -- the basis shape and are tangent to the face
            -- against which the feature is built.
            -- The list provides the information necessary for
            -- subsequent addition of fillets. It may be an empty list.
            -- If an edge is tangent, no fillet is possible, and
            -- the edge must subsequently be removed if you want to add a fillet.
    returns ListOfShape from TopTools;
             ---C++: return const&

    CheckPoint(me: in out;
                   e        : Edge  from TopoDS;
               bnd      : Real  from Standard;
               Pln      : Plane from Geom)
    returns Pnt from gp
    is static protected;


    Normal(me: in out;
               F : Face from TopoDS;
           P : Pnt from gp)
    returns Dir from gp
    is static protected;
    
            
    IntPar(myclass; 
               C    : Curve from Geom;
           P    : Pnt   from gp)
    returns Real from Standard;
    
    
    EdgeExtention(me: in out;
                          e         : in out Edge from TopoDS;
                  bnd       : Real from Standard;
                  FirstLast : Boolean from Standard)
    is static protected;
    
    
    ChoiceOfFaces(myclass;
                          faces : in out ListOfShape from TopTools;
                  cc    : Curve from Geom;
                  par   : Real  from Standard;
                  bnd   : Real  from Standard;
                  Pln   : Plane from Geom)
    returns Face from TopoDS;


    HeightMax(me: in out; 
                  theSbase  : Shape from TopoDS;
              theSUntil : Shape from TopoDS;
              p1        : in out Pnt   from gp;
              p2        : in out Pnt   from gp)
    returns Real from Standard
    is static protected;
        
    ExtremeFaces(me: in out;
                         RevolRib  : Boolean from Standard;
                 bnd       : Real    from Standard;
                 Pln       : Plane   from Geom;
                 FirstEdge : in out Edge from TopoDS;
                 LastEdge  : in out Edge from TopoDS;
                 FirstFace : in out Face from TopoDS;
                 LastFace  : in out Face from TopoDS;
                 FirstVertex : in out Vertex  from TopoDS;
                 LastVertex  : in out Vertex  from TopoDS;
                 OnFirstFace : in out Boolean from Standard;
                 OnLastFace  : in out Boolean from Standard;
                 PtOnFirstEdge : in out Boolean from Standard;
                 PtOnLastEdge  : in out Boolean from Standard;
                 OnFirstEdge : in out Edge from TopoDS;
                 OnLastEdge  : in out Edge from TopoDS)                        
    returns Boolean from Standard
    is static protected;
    
             
    PtOnEdgeVertex(me: in out;
                           RevolRib  : Boolean from Standard;
                   shape     : Shape   from TopoDS;
                   point     : Pnt     from gp;
                   FirstVertex : Vertex  from TopoDS;
                   LastVertex  : Vertex  from TopoDS;
                   PtOnEdge  : in out Boolean from Standard;
                   OnEdge    : in out Edge    from TopoDS;
                   PtOnVertex  : in out Boolean from Standard;
                   OnVertex    : in out Vertex  from TopoDS)
    is static protected;
    
    
    SlidingProfile(me: in out;
                           Prof      : in out Face from TopoDS;
                   RevolRib  : Boolean from Standard;
                   myTol     : Real from Standard;
                   Concavite : in out Integer from Standard;
                   myPln     : Plane   from Geom;
                   BndFace   : Face from TopoDS;
                   CheckPnt  : Pnt  from gp;
                   FirstFace : Face from TopoDS;
                   LastFace  : Face from TopoDS;
                   FirstVertex : Vertex  from TopoDS;
                   LastVertex  : Vertex  from TopoDS;
                   FirstEdge : Edge from TopoDS;
                   LastEdge  : Edge from TopoDS)
    returns Boolean from Standard
    is static protected;
    
        
    NoSlidingProfile(me: in out;
                             Prof      : in out Face from TopoDS;
                     RevolRib  : Boolean from Standard;
                     myTol     : Real from Standard;
                     Concavite : in out Integer from Standard;
                     myPln     : Plane   from Geom;
                     bnd       : Real from Standard;
                     BndFace   : Face from TopoDS;
                     CheckPnt  : Pnt  from gp;
                     FirstFace : Face from TopoDS;
                     LastFace  : Face from TopoDS;
                     FirstVertex : Vertex  from TopoDS;
                     LastVertex  : Vertex  from TopoDS;
                     FirstEdge : Edge from TopoDS;
                     LastEdge  : Edge from TopoDS;
                     OnFirstFace : Boolean from Standard;
                     OnLastFace  : Boolean from Standard)
    returns Boolean from Standard
    is static protected;
    
        
    UpdateDescendants(me: in out; G: Gluer from LocOpe)
    
    is static protected;
            ---Purpose: Updates the data structures of descendant
            -- shapes during the glueing operation.Returns the modified, generated
            --   and deleted faces during the course of the glueing operation.

    UpdateDescendants(me: in out; 
                       B        : HBuilder from TopOpeBRepBuild;
                       SResult  : Shape    from TopoDS;
                       SkipFace : Boolean  from Standard = Standard_False)
    
    is static protected;
 
--modified by NIZNHY-PKV Thu Mar 21 18:42:53 2002  f
    UpdateDescendants(me: in out;  
                   aBOP: BooleanOperation from BRepAlgoAPI;   
               SResult  : Shape    from TopoDS;
               SkipFace : Boolean  from Standard = Standard_False)
            is static protected;
--modified by NIZNHY-PKV Thu Mar 21 18:42:50 2002  t

    CurrentStatusError(me)
    returns StatusError from BRepFeat;

fields

    myFirstPnt : Pnt                      from gp is protected;
    myLastPnt  : Pnt                      from gp is protected;
    myFuse    : Boolean                   from Standard is protected;
    mySliding : Boolean                   from Standard is protected;
    myMap     : DataMapOfShapeListOfShape from TopTools is protected;
    myLFMap   : DataMapOfShapeListOfShape from TopTools is protected;
    myFShape  : Shape                     from TopoDS   is protected;
    myLShape  : Shape                     from TopoDS   is protected;
    
    myPerfSelection: PerfSelection        from BRepFeat is protected;
    
    myWire    : Wire                      from TopoDS is protected;
    mySbase   : Shape                     from TopoDS is protected;
    mySkface  : Face                      from TopoDS is protected;
    myPbase   : Face                      from TopoDS is protected;
    myGShape  : Shape                     from TopoDS is protected;
    mySUntil  : Shape                     from TopoDS is protected;
    myGluedF  : DataMapOfShapeShape       from TopTools is protected;
    myNewEdges: ListOfShape               from TopTools is protected; 
    myTgtEdges: ListOfShape               from TopTools is protected;
    myFacesForDraft: ListOfShape          from TopTools is protected;
    
    myStatusError : StatusError           from BRepFeat is protected;
       
end RibSlot;
