-- Created on: 1997-04-11
-- Created by: VAUTHIER Jean-Claude
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class NamedShape from PNaming inherits Attribute from PDF

	---Purpose: This is the persistent attribute of the
	--          topological naming.

uses

    HArray1OfShape1 from PTopoDS,
    HArray1OfInteger from PColStd


is


    Create returns mutable NamedShape from PNaming;
	---Purpose: Creates a mutable NamedShape from PNaming.

    
    NbShapes(me) returns Integer;
	---Purpose: Returns the number of shapes.


    OldShapes(me : mutable; theShapes : HArray1OfShape1 from PTopoDS);
	---Purpose: Sets the field <myOldShapes>.
    
    OldShapes(me) returns HArray1OfShape1 from PTopoDS;
	---Purpose: Returns the field <myOldShapes>.
    

    NewShapes(me : mutable; theShapes : HArray1OfShape1 from PTopoDS);
	---Purpose: Sets the field <myNewShapes>.
    
    NewShapes(me) returns HArray1OfShape1 from PTopoDS;
	---Purpose: Returns the field <myNewShapes>.
    

    ShapeStatus(me : mutable; theShapeStatus : Integer from Standard);
	---Purpose: Sets the field <myShapeStatus>.
    
    ShapeStatus(me) returns Integer from Standard;
	---Purpose: Returns the field <myShapeStatus>.
    
    Version (me : mutable; theVersion : Integer from Standard);
    	---Purpose: Sets the field <myVersion>.
    
    Version (me) returns Integer from Standard;
        ---Purpose: Returns the field <myVersion>.
	    
fields

    myOldShapes    : HArray1OfShape1 from PTopoDS;
    myNewShapes    : HArray1OfShape1 from PTopoDS;
    myShapeStatus  : Integer         from Standard;
    myVersion      : Integer         from Standard;

end NamedShape;
