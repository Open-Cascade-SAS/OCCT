-- Created on: 1994-05-26
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class GeometryData from TopOpeBRepDS 

    ---Purpose: mother-class of SurfaceData, CurveData, PointData 

uses

    Interference from TopOpeBRepDS,
    ListOfInterference from TopOpeBRepDS

is

    Create returns GeometryData from TopOpeBRepDS; 
     
--modified by NIZNHY-PKV Tue Oct 30 09:24:30 2001  f 
    Create  (Other:GeometryData from TopOpeBRepDS) 
    	returns GeometryData from TopOpeBRepDS;  
    
    Assign (me:out; 
    	    Other:GeometryData from TopOpeBRepDS); 
    ---C++: alias operator=	 
--modified by NIZNHY-PKV Tue Oct 30 09:24:33 2001  t

    Interferences(me) returns ListOfInterference from TopOpeBRepDS
    ---C++: return const &
    is static;

    ChangeInterferences(me : in out) 
    returns ListOfInterference from TopOpeBRepDS
    ---C++: return &
    is static;
    
    AddInterference(me : in out; I : Interference from TopOpeBRepDS)
    is static;
    
fields

    myInterferences : ListOfInterference from TopOpeBRepDS;
    
end GeometryData from TopOpeBRepDS;
