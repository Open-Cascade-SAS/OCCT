-- Created on: 1999-11-29
-- Created by: Peter KURNEV
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Tools2d from TopOpeBRepBuild 

	---Purpose: 

uses
    IndexedDataMapOfShapeVertexInfo from TopOpeBRepBuild,
    Wire  from  TopoDS,
    ListOfShape from TopTools 
    
is

   MakeMapOfShapeVertexInfo  (myclass;  
    aWire:Wire  from  TopoDS;
    aMap:out  IndexedDataMapOfShapeVertexInfo  from  TopOpeBRepBuild);

   DumpMapOfShapeVertexInfo   (myclass;   
    aMap: IndexedDataMapOfShapeVertexInfo  from  TopOpeBRepBuild);


   Path  (myclass; aWire:Wire  from  TopoDS; aResList:out  ListOfShape from TopTools);
    
end Tools2d;
