-- Created on: 1993-01-09
-- Created by: CKY / Contract Toubro-Larsen (Arun MENON)
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package IGESBasic


        ---Purpose : This package represents basic entities from IGES

uses

        Standard,
        TCollection,
        gp,
	TColgp,
	TColStd,
	Message,
        Interface,
        IGESData

is

        class SubfigureDef;

        class Group;

        class GroupWithoutBackP;

        class SingleParent;

        class ExternalRefFileIndex;

        class OrderedGroup;

        class OrderedGroupWithoutBackP;

        class Hierarchy;

        class ExternalReferenceFile;

        class Name;

        class AssocGroupType;

        class SingularSubfigure;

        class ExternalRefFileName;

        class ExternalRefFile;

        class ExternalRefName;

        class ExternalRefLibName;

    	--    Tools for Entities    --

        class ToolSubfigureDef;
        class ToolGroup;
        class ToolGroupWithoutBackP;
        class ToolSingleParent;
        class ToolExternalRefFileIndex;
        class ToolOrderedGroup;
        class ToolOrderedGroupWithoutBackP;
        class ToolHierarchy;
        class ToolExternalReferenceFile;
        class ToolName;
        class ToolAssocGroupType;
        class ToolSingularSubfigure;
        class ToolExternalRefFileName;
        class ToolExternalRefFile;
        class ToolExternalRefName;
        class ToolExternalRefLibName;

    -- Definition and Exploitation of Entities defined in this Package

    class Protocol;
    class ReadWriteModule;
    class GeneralModule;
    class SpecificModule;

    -- The class instantiations :

    class Array2OfHArray1OfReal    instantiates 
        Array2 from TCollection (HArray1OfReal from TColStd);
    class Array1OfLineFontEntity instantiates
        Array1 from TCollection (LineFontEntity from IGESData);

    class HArray1OfHArray1OfInteger instantiates
    	JaggedArray from Interface (HArray1OfInteger     from TColStd);
    -- HArray1 from TCollection (HArray1OfInteger from TColStd,Array1OfHArray1OfInteger);
    class HArray1OfHArray1OfReal    instantiates
    	JaggedArray from Interface (HArray1OfReal        from TColStd);
    -- HArray1 from TCollection (HArray1OfReal from TColStd,Array1OfHArray1OfReal);
    class HArray1OfHArray1OfXY      instantiates
    	JaggedArray from Interface (HArray1OfXY          from TColgp);
    -- HArray1 from TCollection (HArray1OfXY   from TColgp, Array1OfHArray1OfXY);
    class HArray1OfHArray1OfXYZ     instantiates
    	JaggedArray from Interface (HArray1OfXYZ         from TColgp);
    -- HArray1 from TCollection (HArray1OfXYZ  from TColgp, Array1OfHArray1OfXYZ);

    class HArray2OfHArray1OfReal    instantiates HArray2 from TCollection
    	 (HArray1OfReal from TColStd,Array2OfHArray1OfReal);

    class HArray1OfHArray1OfIGESEntity instantiates
    	JaggedArray from Interface (HArray1OfIGESEntity  from IGESData);
    -- HArray1 from TCollection (HArray1OfIGESEntity from IGESData,Array1OfHArray1OfIGESEntity);

    class HArray1OfLineFontEntity   instantiates HArray1 from TCollection
    	 (LineFontEntity from IGESData,Array1OfLineFontEntity);

    --  Package methods 

    Init;
    ---Purpose : Prepares dynqmic data (Protocol, Modules) for this package

    Protocol  returns Protocol from IGESBasic;
    ---Purpose : Returns the Protocol for this Package

end IGESBasic;
