-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package PShort 

uses PCollection,
     TCollection,
     TShort

is


--                             Instantiations de PCollection          --
--                             *****************************          --
------------------------------------------------------------------------

--
--       Instantiations HSequence 
--       **************************************************
--       
class HSequenceOfShortReal instantiates 
           HSequence from PCollection(ShortReal);

--
--       Instantiations HArray1
--       ****************************************************
--       
-----

    class HArray1OfShortReal instantiates 
                        HArray1 from PCollection(ShortReal);
--    class Array1FromHArray1OfShortReal instantiates 
--    	  Array1FromHArray1(ShortReal
--                           ,Array1OfShortReal from TShort
--                           ,HArray1OfShortReal from PShort);

--
--       Instantiations HArray2
--       ****************************************************
--       

    class HArray2OfShortReal instantiates 
                        HArray2 from PCollection(ShortReal);
--    class Array2FromHArray2OfShortReal instantiates 
--    	  Array2FromHArray2(ShortReal
--                           ,Array2OfShortReal from TShort
--                           ,HArray2OfShortReal from PShort);


end PShort;
