-- Created on: 1992-08-24
-- Created by: Ramin BARRETO
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class AncestorIterator from Standard
    ---Purpose:
    -- The class <AncestorIterator> is a iterator which provides 
    -- information about inheritance. 
    -- An AncestorIterator object is used to scan sequentially the 
    -- hierarchy of a type object from its direct super-type to the root.
    --
    -- Warning:
    --   The near parents are first.
    --   
uses 
    Boolean from Standard
   ,Integer from Standard
   ,Type from Standard

raises 
    NoMoreObject from Standard
   
is

    ------------------------------------------------------------------------
    ---Category: The Constructur of AncestorIterator.
    ------------------------------------------------------------------------
    Create(anOther: AncestorIterator )  returns AncestorIterator;
    ---Purpose:
    --   The copy constructor for a AncestorIterator . 
    --   
    ---Level: Advanced    
       
    Create(aType: Type) returns AncestorIterator;
    ---Purpose: 
    --   Creates an iterator on the type <aType>.
    --   Set the iterator at the beginning of the ancestors; 
    --   this means near parents are first.
    ---Level: Advanced  
   
    ------------------------------------------------------------------------
    ---Category: Assignation.
    ------------------------------------------------------------------------
    Assign(me: in out; anOther: AncestorIterator); 
    ---Purpose:
    --   Assigns an  AncestorIterator from another AncestorIterator.
    --
    ---C++: alias operator =        
    ---Level: Advanced        
          
    ------------------------------------------------------------------------
    ---Category: The methods for iterating.
    ------------------------------------------------------------------------

    More(me) returns Boolean;
    ---Purpose: 
    -- Returns True if there are other ancestors.
    --
    -- Example:
    --
    -- Handle(Standard_Type) type;
    -- Standard_AncestorIterator super(TYPE(Geom_Circle));
    -- while(super.More()) { type = super.Value();
    --      super.Next();
    -- }  

    Next(me: in out) 
    ---Purpose: 
    -- Moves the position of the iterator to the next super-type. 
    -- If the current position corresponds to a root class, it becomes undefined.
    --
    -- Exceptions:
    -- Standard_NoMoreObject if the position of the iterator is undefined
    raises NoMoreObject; -- If there are no more ancestors.
    ---Level: Advanced  
          
    ------------------------------------------------------------------------
    ---Category: The information of each ancestor.
    ------------------------------------------------------------------------

    Iterator(me) returns AncestorIterator
    ---Purpose: 
    --   Returns an <AncestorIterator> corresponding to the current position 
    --   of the iterator.
    raises NoMoreObject; -- If there are no more Ancestors.
    ---Level: Advanced  

    Value(me) returns Type 
    ---Purpose:
    -- Returns the type corresponding to the current position of 
    -- the iterator.
    --
    -- Example:
    --
    -- Standard_AncestorIterator super(TYPE(Geom_Circle));
    -- assert (super.Value() == TYPE(Geom_Conic));
    --
    -- Exceptions:
    -- Standard_NoSuchObject if the position of the iterator is undefined.
    raises NoMoreObject; -- If there are no more ancestors.
   
fields

    myType  : Type;
    myNbIter: Integer;
   
end AncestorIterator from Standard;
