-- Created on: 1995-12-01
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DrawableC3D from TestTopOpeDraw inherits Curve from DrawTrSurf

    ---Purpose: 

uses  

    Interpretor from Draw,
    Curve from Geom,
    Color from Draw,
    Display from Draw,
    Text3D from Draw,
    CString from Standard,
    Pnt from gp

is

    Create (C : Curve from Geom; CColor : Color from Draw)
    returns mutable DrawableC3D from TestTopOpeDraw;

    Create (C : Curve from Geom; CColor : Color from Draw;
    	    Text : CString; TextColor : Color from Draw)
    returns mutable DrawableC3D from TestTopOpeDraw;

    Create (C : Curve from Geom; CColor : Color from Draw;
    	    Text : CString; TextColor : Color from Draw;
    	    Discret : Integer; Deflection : Real; DrawMode : Integer;
    	    DispOrigin : Boolean from Standard = Standard_True)
    returns mutable DrawableC3D from TestTopOpeDraw;

    Pnt(me) returns Pnt from gp is virtual;
    
    ChangePnt(me : mutable; P : Pnt);
    
    ChangeCurve(me : mutable; C : Curve from Geom);
    
    ChangeText(me : mutable; T : CString from Standard);
    
    Name(me : mutable; N : CString) is redefined;
    
    Whatis(me; I : in out Interpretor from Draw) is redefined;
    ---Purpose: For variable whatis command.

    DrawOn(me; dis : in out Display from Draw) is redefined;
    
fields

    myText3D : Text3D from Draw is protected;
    myText :CString from Standard is protected;
    myTextColor : Color from Draw;

end DrawableC3D;
