-- Created on: 1998-07-22
-- Created by: Christian CAILLET
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Vars  from XSControl    inherits TShared  from MMgt

    ---Purpose : Defines a receptacle for externally defined variables, each
    --           one has a name
    --           
    --           I.E. a WorkSession for XSTEP is generally used inside a
    --           context, which brings variables, especially shapes and
    --           geometries. For instance DRAW or an application engine
    --           
    --           This class provides a common form for this. It also provides
    --           a default implementation (locally recorded variables in a
    --           dictionary), but which is aimed to be redefined

uses CString, Transient, DictionaryOfTransient,
     Pnt from gp, Pnt2d from gp,
     Geometry from Geom, Curve from Geom, Curve from Geom2d, Surface from Geom,
     Shape from TopoDS

is

    Create returns mutable Vars;

    Set (me : mutable; name : CString; val : Transient)  is virtual;

    Get (me; name : in out CString) returns Transient  is virtual;


    GetGeom (me; name : in out CString) returns Geometry  is virtual;

    GetCurve2d (me; name : in out CString) returns Curve from Geom2d  is virtual;

    GetCurve   (me; name : in out CString) returns Curve from Geom  is virtual;

    GetSurface (me; name : in out CString) returns Surface from Geom  is virtual;

    SetPoint   (me : mutable; name : CString; val : Pnt   from gp)  is virtual;

    SetPoint2d (me : mutable; name : CString; val : Pnt2d from gp)  is virtual;

    GetPoint   (me; name : in out CString; pnt : out Pnt   from gp) returns Boolean  is virtual;

    GetPoint2d (me; name : in out CString; pnt : out Pnt2d from gp) returns Boolean  is virtual;


    SetShape   (me : mutable; name : CString; val : Shape from TopoDS)  is virtual;

    GetShape   (me; name : in out CString) returns Shape from TopoDS  is virtual;

fields

    thevars : DictionaryOfTransient;

end Vars;
