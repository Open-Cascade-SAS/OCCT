-- File:	StepAP203_CcDesignSpecificationReference.cdl
-- Created:	Fri Nov 26 16:26:33 1999 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0
-- Copyright:	Matra Datavision 1999

class CcDesignSpecificationReference from StepAP203
inherits DocumentReference from StepBasic

    ---Purpose: Representation of STEP entity CcDesignSpecificationReference

uses
    Document from StepBasic,
    HAsciiString from TCollection,
    HArray1OfSpecifiedItem from StepAP203

is
    Create returns CcDesignSpecificationReference from StepAP203;
	---Purpose: Empty constructor

    Init (me: mutable; aDocumentReference_AssignedDocument: Document from StepBasic;
                       aDocumentReference_Source: HAsciiString from TCollection;
                       aItems: HArray1OfSpecifiedItem from StepAP203);
	---Purpose: Initialize all fields (own and inherited)

    Items (me) returns HArray1OfSpecifiedItem from StepAP203;
	---Purpose: Returns field Items
    SetItems (me: mutable; Items: HArray1OfSpecifiedItem from StepAP203);
	---Purpose: Set field Items

fields
    theItems: HArray1OfSpecifiedItem from StepAP203;

end CcDesignSpecificationReference;
