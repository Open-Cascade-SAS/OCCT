-- Created on: 1999-07-12
-- Created by: Denis PASCAL
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

private class Owner from TDocStd inherits Attribute from TDF

	---Purpose: 

uses Attribute from TDF,
     GUID      from Standard, 
     RelocationTable from TDF, 
     Data      from TDF,
     Label     from TDF,
     Document  from TDocStd

is 

    ---Purpose: class methods
    --          =============

    GetID (myclass)   
    	---C++: return const &  
    returns GUID from Standard;

    SetDocument (myclass; indata : Data from TDF; doc : Document from TDocStd);
    
    GetDocument (myclass; ofdata : Data from TDF)
    returns Document from TDocStd;

    ---Purpose: Owner methods
    --          ===============
    
    Create
    returns Owner from TDocStd;  
    
    SetDocument (me : mutable; document : Document from TDocStd);    

    GetDocument (me)
    returns Document from TDocStd;
    
    ---Category: methodes de TDF_Attribute
    --           =========================
    
    ID (me)
    	---C++: return const & 
    returns GUID from Standard;

    Restore (me: mutable; With : Attribute from TDF);

    NewEmpty (me)
    returns Attribute from TDF;

    Paste (me; Into : Attribute from TDF;
	       RT   : RelocationTable from TDF);    

    Dump(me; anOS : in out OStream from Standard)
    	returns OStream from Standard
    	is redefined;
	---C++: return &

fields

    myDocument : Document from TDocStd;

end Owner;
