-- File:	Dynamic_ObjectParameter.cdl
-- Created:	Fri Dec 24 10:26:25 1993
-- Author:	Gilles DEBARBOUILLE
--		<gde@mastox>
---Copyright:	 Matra Datavision 1993

class ObjectParameter from Dynamic

inherits

    Parameter from Dynamic     
    
	---Purpose: This  inherited class from Parameter describes all
	--          the parameters, which   are characterized   by  an
	--          object value.

    
uses
    OStream from Standard,
    CString from Standard 

is

    Create(aparameter : CString from Standard) returns mutable ObjectParameter from Dynamic;
    
    ---Level: Public 
    
    ---Purpose: Creates an ObjectParameter with <aparameter> as name.
    
    Create(aparameter : CString from Standard; anobject : any Transient)
    
    ---Level: Public 
    
    ---Purpose: With  the name of  the  Parameter <aparameter> and the
    --          object  <anobject>,      creates an   instance      of
    --          ObjectParameter.
    
    returns mutable ObjectParameter from Dynamic;
    
    Value(me) returns any Transient
    
    ---Level: Public 
    
    ---Purpose: Returns the value of the parameter which is an object.
    
    is static;

    Value (me : mutable ; anobject : Transient)
    
    ---Level: Public 
    
    --- Purpose: Sets the object <anobject> in <me>.

    is static;
    
    Dump(me ; astream : in out OStream from Standard)
    
    ---Level: Internal 
    
    ---Purpose: Useful for debugging.
    
    is redefined;
    
fields

    theobject : Transient;

end ObjectParameter;
