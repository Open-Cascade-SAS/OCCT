-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ShellBasedSurfaceModel from StepShape 

inherits GeometricRepresentationItem from StepGeom

uses

	HArray1OfShell from StepShape, 
	Shell from StepShape, 
	HAsciiString from TCollection
is

	Create returns mutable ShellBasedSurfaceModel;
	---Purpose: Returns a ShellBasedSurfaceModel


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aSbsmBoundary : mutable HArray1OfShell from StepShape) is virtual;

	-- Specific Methods for Field Data Access --

	SetSbsmBoundary(me : mutable; aSbsmBoundary : mutable HArray1OfShell);
	SbsmBoundary (me) returns mutable HArray1OfShell;
	SbsmBoundaryValue (me; num : Integer) returns Shell;
	NbSbsmBoundary (me) returns Integer;

fields

	sbsmBoundary : HArray1OfShell from StepShape; -- a SelectType

end ShellBasedSurfaceModel;
