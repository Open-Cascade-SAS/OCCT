-- File:        UniformSurfaceAndRationalBSplineSurface.cdl
-- Created:     Mon Dec  4 12:02:34 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWUniformSurfaceAndRationalBSplineSurface from RWStepGeom

	---Purpose : Read & Write Module for UniformSurfaceAndRationalBSplineSurface

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     UniformSurfaceAndRationalBSplineSurface from StepGeom,
     EntityIterator from Interface

is

	Create returns RWUniformSurfaceAndRationalBSplineSurface;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable UniformSurfaceAndRationalBSplineSurface from StepGeom);

	WriteStep (me; SW : in out StepWriter; ent : UniformSurfaceAndRationalBSplineSurface from StepGeom);

	Share(me; ent : UniformSurfaceAndRationalBSplineSurface from StepGeom; iter : in out EntityIterator);

end RWUniformSurfaceAndRationalBSplineSurface;
