-- Created on: 1993-04-29
-- Created by: Gerard GRAS
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class TextManager from MFT inherits TShared from MMgt

---Purpose: defines the common behaviour of the MFT output driver. 
--  Warning: Permits to receives draw primitives from the FontManager
--	    at DrawText(...) time.
--	    This class must be redefined by the user as an application class
--	    connected to a user driver.

uses
	FontManager	from MFT,
	PlaneAngle      from Quantity,
	Length          from Quantity

is


        -------------------------
        -- Category: Constructors
        -------------------------

	Create returns TextManager from MFT;
        ---Purpose: Does NOTHING 

        -------------------------
	-- Category: Draw methods
        -------------------------

        BeginString (me: mutable;
		X,Y: Length from Quantity;
		anOrientation: PlaneAngle from Quantity;
		aWidth,aHeight: Length from Quantity;
		aSlant: PlaneAngle from Quantity;
		aPaintType: Integer from Standard) is virtual;
        ---Purpose: Calls when string drawing is started.
	--	    with a string aspect <aPaintType> :
	--	      0 for filled string
	--	      1 for stroke string
	--	      2 for outline string 
	--	    The origine of the string <X>,<Y>,
	--	    The orientation of the string <anOrientation>,
	--	    The medium size of the char <aWidth,aHeight>,
	--	    The Slant of the char <aSlant>,

        BeginChar (me: mutable;
		aCharCode: Integer from Standard;
		X,Y: Length from Quantity) 
		returns Boolean from Standard is virtual;
        ---Purpose: Calls when a char drawing is started 
	--	    and give the relative char start position from the beginning
	--	    of the string.
	--	    The application can returns FALSE for skipping the char drawing.

        SetCharBoundingBox (me: mutable;
		X1,Y1,X2,Y2,X3,Y3,X4,Y4: Length from Quantity) 
		returns Boolean from Standard is virtual;
        ---Purpose: Calls to defines the current char bounding-box with :
	--	     X1,Y1 : the lower left corner of the box,
	--	     X2,Y2 : the lower right corner of the box,
	--	     X3,Y3 : the upper right corner of the box,
	--	     X4,Y4 : the upper left corner of the box.
	--  Warning: the char bounding box is not rectangular when the Slant is != 0.
	--	    The application can returns FALSE for skipping the char drawing.

	SetCharEncoding (me: mutable;
		anEncoding: CString from Standard) 
		returns Boolean from Standard is virtual;
        ---Purpose: Calls to defines the current char encoding.
	--  Warning: The application can returns FALSE for skipping the char drawing.

        Moveto (me: mutable;
		X,Y: Length from Quantity) 
		returns Boolean from Standard is virtual;
        ---Purpose: Calls to sets the current string position. 
	--	    The application can returns FALSE for skipping the char drawing.

        Lineto (me: mutable;
		X,Y: Length from Quantity) 
		returns Boolean from Standard is virtual;
        ---Purpose: Calls to drawn to the current string position. 
	--	    The application can returns FALSE for skipping the char drawing.
        Curveto (me: mutable;
		X1,Y1,X2,Y2,X3,Y3,X4,Y4: Length from Quantity) 
		returns Boolean from Standard is virtual;
        ---Purpose: Calls to drawn to the current string position. 
	--	    The application can drawn the curve defined by
	--	    his descriptor P1,P2,P3,P4 or
	--	    returns FALSE to let the interpretor compute the curve
	--	    vectors.

        ClosePath (me: mutable) is virtual;
        ---Purpose: Calls when a char path drawing is ended 

        EndChar (me: mutable;
		X,Y: Length from Quantity) 
		returns Boolean from Standard is virtual;
        ---Purpose: Calls when a char drawing is ended 
	--	    and give the relative char ending position from the 
	--	    beginning of the string.
	--	    The application can returns FALSE for skipping the string 
	--	    drawing.

        EndString (me: mutable ) is virtual;
        ---Purpose: Calls when string drawing is ended (Normally the last call).
 
        -------------------------
	-- Category: Private methods
        -------------------------

	MinMax (myclass;
		Xmin,Ymin,Xmax,Ymax: out Length from Quantity)
		is private;
        ---Purpose: Returns the current drawn string min-max.

	Encoding (myclass)
		returns CString from Standard is private;
        ---Purpose: Returns the current drawn char encoding.

friends
	class FontManager from MFT

end TextManager from MFT;
