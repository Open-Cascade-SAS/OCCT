-- Created on: 1990-12-17
-- Created by: Remi Lequette
-- Copyright (c) 1990-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.





class TWire1 from PTopoDS  inherits TShape1 from PTopoDS

	---Purpose: a Topological  Wire1 is a  structure of Edge1s.  The
	--          Edge1s may have 2D curves stored with them. This is
	--          a curve in the parametric space of a Surface.

uses
    ShapeEnum from TopAbs

is
    Create returns mutable TWire1;
    	---Level: Internal 

    ShapeType(me) returns ShapeEnum from TopAbs;
    	---Level: Internal 

end TWire1;


