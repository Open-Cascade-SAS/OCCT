-- Created on: 1993-01-11
-- Created by: Christophe MARION
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class EdgeIterator from HLRAlgo

uses
    EdgeStatus from HLRAlgo,
    Address    from Standard,
    Integer    from Standard,
    Boolean    from Standard,
    ShortReal  from Standard,
    Real       from Standard

is
    Create returns EdgeIterator from HLRAlgo;
	---Purpose: Iterator  on the  visible or  hidden  parts of  an
	--          edge.
    
    InitHidden(me : in out; status : EdgeStatus from HLRAlgo)
    is static;
    
    MoreHidden(me) returns Boolean from Standard
    	---C++: inline
    is static;
    
    NextHidden(me : in out)
    is static;
    
    Hidden(me; Start    : out Real      from Standard;
               TolStart : out ShortReal from Standard;
               End      : out Real      from Standard;
               TolEnd   : out ShortReal from Standard)
	---C++: inline
	---Purpose: Returns the bounds and the tolerances
	--          of the current Hidden Interval
    is static;
    
    InitVisible(me : in out; status : EdgeStatus from HLRAlgo)
	---C++: inline
    is static;
    
    MoreVisible(me) returns Boolean from Standard
    	---C++: inline
    is static;
    
    NextVisible(me : in out)
	---C++: inline
    is static;
    
    Visible(me : in out;
            Start    : out Real      from Standard;
            TolStart : out ShortReal from Standard;
            End      : out Real      from Standard;
            TolEnd   : out ShortReal from Standard)
	---C++: inline
	---Purpose: Returns the bounds and the tolerances
	--          of the current Visible Interval
    is static;
    
fields
    myNbVis       : Integer   from Standard;
    myNbHid       : Integer   from Standard;
    EVis          : Address   from Standard;
    EHid          : Address   from Standard;
    iVis          : Integer   from Standard;
    iHid          : Integer   from Standard;
    myHidStart    : Real      from Standard;
    myHidEnd      : Real      from Standard;
    myHidTolStart : ShortReal from Standard;
    myHidTolEnd   : ShortReal from Standard;

end EdgeIterator;
