-- Created on: 2003-06-04
-- Created by: Galina KULIKOVA
-- Copyright (c) 2003-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class GeometricToleranceWithDatumReference from StepDimTol
inherits GeometricTolerance from StepDimTol

    ---Purpose: Representation of STEP entity GeometricToleranceWithDatumReference

uses
    HAsciiString from TCollection,
    MeasureWithUnit from StepBasic,
    ShapeAspect from StepRepr,
    HArray1OfDatumReference from StepDimTol

is
    Create returns GeometricToleranceWithDatumReference from StepDimTol;
	---Purpose: Empty constructor

    Init (me: mutable; aGeometricTolerance_Name: HAsciiString from TCollection;
                       aGeometricTolerance_Description: HAsciiString from TCollection;
                       aGeometricTolerance_Magnitude: MeasureWithUnit from StepBasic;
                       aGeometricTolerance_TolerancedShapeAspect: ShapeAspect from StepRepr;
                       aDatumSystem: HArray1OfDatumReference from StepDimTol);
	---Purpose: Initialize all fields (own and inherited)

    DatumSystem (me) returns HArray1OfDatumReference from StepDimTol;
	---Purpose: Returns field DatumSystem
    SetDatumSystem (me: mutable; DatumSystem: HArray1OfDatumReference from StepDimTol);
	---Purpose: Set field DatumSystem

fields
    theDatumSystem: HArray1OfDatumReference from StepDimTol;

end GeometricToleranceWithDatumReference;
