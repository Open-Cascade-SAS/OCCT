-- Created on: 1992-01-21
-- Created by: GG
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Update: 	FDA Oct 15 1994, 
--		ZOV - Mars 30 1998


class AmbientLight from V3d

    	---Purpose: Creation of an ambient light source in a viewer.


inherits Light from V3d

uses 

	Viewer from V3d,
        TypeOfRepresentation from V3d,
	NameOfColor from Quantity,
	View from V3d,
	Coordinate from V3d,
	Structure from Graphic3d,
	Vertex from Graphic3d,
	Group from Graphic3d

is

    	Create ( VM : mutable Viewer ;
		 Color : NameOfColor = Quantity_NOC_WHITE ) 
				returns mutable AmbientLight;
	---Purpose: Constructs an ambient light source in the viewer VM.
    	-- The default Color of this light source is WHITE.

end AmbientLight;
