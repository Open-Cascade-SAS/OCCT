-- File:	StepData_FieldList.cdl
-- Created:	Tue Apr  1 13:11:37 1997
-- Author:	Christian CAILLET
--		<cky@heliox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1997


class FieldList  from StepData

    ---Purpose : Describes a list of fields, in a general way
    --           This basic class is for a null size list
    --           Subclasses are for 1, N (fixed) or Dynamic sizes

uses Field from StepData, EntityIterator from Interface

raises OutOfRange

is

    Create returns FieldList;
    ---Purpose : Creates a FieldList of 0 Field

    NbFields (me) returns Integer  is virtual;
    ---Purpose : Returns the count of fields. Here, returns 0

    Field  (me; num : Integer) returns Field
    ---Purpose : Returns the field n0 <num> between 1 and NbFields (read only)
	raises OutOfRange
    --           Error if <num> out of range
    	is virtual;
    ---C++ : return const &

    CField (me : in out; num : Integer) returns Field
    ---Purpose : Returns the field n0 <num> between 1 and NbFields, in order to
    --           modify its content
	raises OutOfRange
    --           Error if <num> out of range
    	is virtual;
    ---C++ : return &

    FillShared (me; iter : in out EntityIterator);
    ---Purpose : Fills an iterator with the entities shared by <me>

end FieldList;
