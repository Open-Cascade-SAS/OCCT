-- Created on: 1993-06-17
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PointIterator from TopOpeBRepDS 
    inherits InterferenceIterator from TopOpeBRepDS

	---Purpose: 

uses

    State from TopAbs,
    Orientation  from TopAbs,
    Interference from TopOpeBRepDS,
    ListOfInterference from TopOpeBRepDS

is

    Create(L : ListOfInterference from TopOpeBRepDS) returns PointIterator;
    ---Purpose: Creates an  iterator on the  points on curves
    --          described by the interferences in <L>.
    
    MatchInterference(me; I : Interference from TopOpeBRepDS) 
    returns Boolean from Standard
    ---Purpose: Returns  True if the Interference <I>  has a 
    --          GeometryType() TopOpeBRepDS_POINT or TopOpeBRepDS_VERTEX
    --          returns False else.
    is redefined;

    Current(me) returns Integer from Standard
    ---Purpose: Index of the point in the data structure.
    is static;
    
    Orientation(me; S : State from TopAbs) 
    returns Orientation from TopAbs
    is static;
    
    Parameter(me) returns Real from Standard
    	-- Edge/Point Interference
    	-- Curve/Point Interference
    	-- Edge/Vertex Interference
    is static;
    
    IsVertex(me) returns Boolean from Standard
    is static;

    IsPoint(me) returns Boolean from Standard
    is static;
    
    DiffOriented(me) returns Boolean from Standard
    is static;

    SameOriented(me) returns Boolean from Standard
    is static;

    Support(me) returns Integer from Standard
    is static;

end PointIterator from TopOpeBRepDS;
