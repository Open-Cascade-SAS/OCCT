-- Created on: 1999-06-22
-- Created by: data exchange team
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class ApplySequence from ShapeProcessAPI 

    ---Purpose: Applies one of the sequence read from resource file.

uses
    
    ShapeEnum           from TopAbs,
    Shape               from TopoDS,
    DataMapOfShapeShape from TopTools,
    Printer             from Message,
    ShapeContext        from ShapeProcess,
    AsciiString         from TCollection
is

    Create (rscName: CString; seqName: CString = "") returns ApplySequence from ShapeProcessAPI;
    	---Purpose: Creates an object and loads resource file and sequence of
    	--          operators given by their names.
    
    Context (me: in out) returns ShapeContext from ShapeProcess;
    	---C++ : return &
	---Purpose: Returns object for managing resource file and sequence of
    	--          operators.
    
    PrepareShape (me: in out; shape  : Shape from TopoDS;
    	    	    	      fillmap: Boolean = Standard_False;
			      until  : ShapeEnum from TopAbs = TopAbs_SHAPE)
    returns Shape from TopoDS;
    	---Purpose: Performs sequence of operators stored in myRsc.
	--          If <fillmap> is True adds history "shape-shape" into myMap
	--          for shape and its subshapes until level <until> (included).
    	--          If <until> is TopAbs_SHAPE,  all the subshapes are considered.
	
    ClearMap (me: in out);
    	---Purpose: Clears myMap with accumulated history.
	
    Map (me) returns DataMapOfShapeShape from TopTools;
    	---C++: return const &
	---Purpose: Returns myMap with accumulated history.

    PrintPreparationResult (me);
    	---Purpose: Prints result of preparation onto the messenger of the context.
	--          Note that results can be accumulated from previous preparations
	--          it method ClearMap was not called before PrepareShape.
	---Remark: At the moment outputs information only on shells and faces.
    
fields

    myContext: ShapeContext from ShapeProcess;
    myMap    : DataMapOfShapeShape from TopTools;
    mySeq    : AsciiString from TCollection;

end ApplySequence;
