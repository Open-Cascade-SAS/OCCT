-- File:	Transfer_DispatchControl.cdl
-- Created:	Thu Jun 17 15:44:03 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class DispatchControl  from Transfer  inherits CopyControl from Interface

    ---Purpose : This is an auxiliary class for TransferDispatch, which allows
    --           to record simple copies, as CopyControl from Interface, but
    --           based on a TransientProcess. Hence, it allows in addition
    --           more actions (such as recording results of adaptations)

uses Transient, TransientProcess, InterfaceModel

raises InterfaceError

is

    Create (model : InterfaceModel; TP : mutable TransientProcess)
    	returns mutable DispatchControl;
    ---Purpose : Creates the DispatchControl, ready for use

    TransientProcess (me) returns mutable TransientProcess;
    ---Purpose : Returns the content of the DispatchControl : it can be used
    --           for a direct call, if the basic methods do not suffice
    ---C++ : return const &

    StartingModel (me) returns any InterfaceModel;
    ---Purpose : Returns the Model from which the transfer is to be done
    ---C++ : return const &

    	--  Now, inherited methods used for Copy (the minimum set)

    Clear (me : mutable);
    ---Purpose : Clears the List of Copied Results

    Bind (me : mutable; ent : Transient; res : mutable Transient)
    ---Purpose : Binds a (Transient) Result to a (Transient) Starting Entity
    	raises InterfaceError;
    --           Error if <ent> is already bound

    Search (me; ent : Transient; res : out mutable Transient)
    	returns Boolean;
    ---Purpose : Searches for the Result bound to a Starting Entity
    --           If Found, returns True and fills <res>
    --           Else, returns False and nullifies <res>

fields

    theTP    : TransientProcess;
    themodel : InterfaceModel;

end DispatchControl;
