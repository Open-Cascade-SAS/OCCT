-- Created on: 1995-10-24
-- Created by: Mister rmi
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package MgtPoly

	---Purpose: This  package   provides   methods  to   translate
	--          transient objects from Poly to  persistent objects
	--          from PPoly and vice-versa.
	--          As far as objects can be shared (just as Geometry),
	--          a map is given as translate argument.


uses Poly,
     PPoly,
     PTColStd
     
is

    -- Triangle (Storable)

    Translate(POjb: Triangle from PPoly)
    	returns Triangle from Poly;
	---Purpose: translates Transient -> Persistent
    
    Translate(TObj: Triangle from Poly)
    	returns Triangle from PPoly;
	---Purpose: translates Persistent -> Transient

    -- Triangulation

    Translate(PObj : Triangulation from PPoly;
    	      aMap : in out PersistentTransientMap from PTColStd)
    	returns Triangulation from Poly;
	---Purpose: translates Persistent -> Transient

    Translate(TObj : Triangulation from Poly;
    	      aMap : in out TransientPersistentMap from PTColStd)
    	returns Triangulation from PPoly;
	---Purpose: translates Transient -> Persistent
    
    -- Polygon3D

    Translate(PObj : Polygon3D from PPoly;
    	      aMap : in out PersistentTransientMap from PTColStd)
    	returns Polygon3D from Poly;
	---Purpose: translates Persistent -> Transient

    Translate(TObj : Polygon3D from Poly;
    	      aMap : in out TransientPersistentMap from PTColStd)
    	returns Polygon3D from PPoly;
	---Purpose: translates Transient -> Persistent

    -- Polygon2D


    Translate(PObj : Polygon2D from PPoly;
    	      aMap : in out PersistentTransientMap from PTColStd)
    	returns Polygon2D from Poly;
	---Purpose: translates Persistent -> Transient

    Translate(TObj : Polygon2D from Poly;
    	      aMap : in out TransientPersistentMap from PTColStd)
    	returns Polygon2D from PPoly;
	---Purpose: translates Transient -> Persistent

    -- PolygonOnTriangulation

    Translate(PObj : PolygonOnTriangulation from PPoly;
    	      aMap : in out PersistentTransientMap from PTColStd)
    	returns PolygonOnTriangulation from Poly;
	---Purpose: translates Persistent -> Transient

    Translate(TObj : PolygonOnTriangulation from Poly;
    	      aMap : in out TransientPersistentMap from PTColStd)
    	returns PolygonOnTriangulation from PPoly;
	---Purpose: translates Transient -> Persistent

end MgtPoly;
