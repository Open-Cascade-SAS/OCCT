-- Created on: 1994-06-16
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class FileName from HeaderSection 

inherits TShared from MMgt

uses

	HAsciiString from TCollection, 
	HArray1OfHAsciiString from Interface
is

	Create returns FileName;
	---Purpose: Returns a FileName

	Init (me : mutable;
	      aName : HAsciiString from TCollection;
	      aTimeStamp : HAsciiString from TCollection;
	      aAuthor : HArray1OfHAsciiString from Interface;
	      aOrganization : HArray1OfHAsciiString from Interface;
	      aPreprocessorVersion : HAsciiString from TCollection;
	      aOriginatingSystem : HAsciiString from TCollection;
	      aAuthorisation : HAsciiString from TCollection);

	-- Specific Methods for Field Data Access --

	SetName(me : mutable; aName : HAsciiString);
	Name (me) returns HAsciiString;
	SetTimeStamp(me : mutable; aTimeStamp : HAsciiString);
	TimeStamp (me) returns HAsciiString;
	SetAuthor(me : mutable; aAuthor : HArray1OfHAsciiString);
	Author (me) returns HArray1OfHAsciiString;
	AuthorValue (me; num : Integer) returns HAsciiString;
	NbAuthor (me) returns Integer;
	SetOrganization(me : mutable; aOrganization : HArray1OfHAsciiString);
	Organization (me) returns HArray1OfHAsciiString;
	OrganizationValue (me; num : Integer) returns HAsciiString;
	NbOrganization (me) returns Integer;
	SetPreprocessorVersion(me : mutable; aPreprocessorVersion : HAsciiString);
	PreprocessorVersion (me) returns HAsciiString;
	SetOriginatingSystem(me : mutable; aOriginatingSystem : HAsciiString);
	OriginatingSystem (me) returns HAsciiString;
	SetAuthorisation(me : mutable; aAuthorisation : HAsciiString);
	Authorisation (me) returns HAsciiString;

fields

	name : HAsciiString from TCollection;
	timeStamp : HAsciiString from TCollection;
	author : HArray1OfHAsciiString from Interface;
	organization : HArray1OfHAsciiString from Interface;
	preprocessorVersion : HAsciiString from TCollection;
	originatingSystem : HAsciiString from TCollection;
	authorisation : HAsciiString from TCollection;

end FileName;
