-- Created on: 1993-06-14
-- Created by: Martine LANGLOIS
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MakeVector from GeomToStep inherits Root from GeomToStep

    ---Purpose: This class implements the mapping between classes 
    --          Vector from Geom, Geom2d and Vec, Vec2d from gp, and the class
    --          Vector from StepGeom which describes a Vector from
    --          Prostep. 
  
uses Vec from gp,
     Vec2d from gp,
     Vector from Geom,
     Vector from Geom2d,
     Vector from StepGeom
     
raises NotDone from StdFail
     
is 

Create ( V : Vec from gp ) returns MakeVector;

Create ( V : Vec2d from gp ) returns MakeVector;

Create ( V : Vector from Geom ) returns MakeVector;

Create ( V : Vector from Geom2d ) returns MakeVector;

Value (me) returns Vector from StepGeom
    raises NotDone
    is static;
    ---C++: return const&

fields

    theVector : Vector from StepGeom;
    	-- The solution from StepGeom
    	
end MakeVector;


