-- Created by: Peter KURNEV
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class IndexRange from BOPDS 

	---Purpose: 
    	-- The class BOPDS_IndexRange is to store  
    	-- the information about range of two indices 
--uses
--raises

is 
    Create 
    	returns IndexRange from BOPDS; 
    ---C++: alias "Standard_EXPORT virtual ~BOPDS_IndexRange();"   
    ---C++: inline 
    	---Purpose:  
    	--- Empty contructor  
    	--- 
	 
    SetFirst(me:out; 
    	    theI1:Integer from Standard); 
    ---C++: inline		 
     	---Purpose: 
    	--- Modifier   
	--- Sets the first index <theI1>  of the range  
	
    SetLast(me:out; 
    	    theI2:Integer from Standard);	 
    ---C++: inline 
    	---Purpose: 
    	--- Modifier   
	--- Sets the second index <theI2>  of the range   
     
    First(me) 
    	returns Integer from Standard; 
    ---C++: inline
	---Purpose: 
    	--- Selector   
	--- Returns the first index of the range  
	
    Last(me) 
    	returns Integer from Standard; 				     
    ---C++: inline
     	---Purpose: 
    	--- Selector   
	--- Returns the second index of the range  
	 
    SetIndices(me:out; 
    	    theI1:Integer from Standard;
    	    theI2:Integer from Standard); 
    ---C++: inline	  
    	---Purpose:  
    	--- Modifier   
	--- Sets the first index of the range  <theI1>
	--- Sets the second index of the range <theI2> 
	     
    Indices(me; 
    	    theI1:out Integer from Standard;
    	    theI2:out Integer from Standard);  
    ---C++: inline     
     	---Purpose:  
    	--- Selector   
	--- Returns the first index of the range  <theI1>
	--- Returns the second index of the range <theI2>  
	
    Contains(me; 
    	    theIndex:Integer from Standard) 
    	returns Boolean from Standard;  
    ---C++: inline	 
     	---Purpose:   
    	--- Query   
	--- Returns true if the range contains <theIndex>
	
    Dump(me);
    
     
    
fields 
    myFirst  :  Integer from Standard is protected;  
    myLast   :  Integer from Standard is protected;  

end IndexRange;
