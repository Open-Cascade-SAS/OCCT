-- Created on: 2012-06-01
-- Created by: Eugeny MALTCHIKOV
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.
 
class Builder from BRepFeat
    inherits BOP from BOPAlgo 
 
    ---Purpose: Provides a basic tool to implement features topological  
    --          operations. The main goal of the algorithm is to perform
    --          the result of the operation according to the  
    --          kept parts of the tool.
    --          Input data: a) DS;
    --                      b) The kept parts of the tool;
    --                         If the map of the kept parts of the tool 
    --                         is not filled boolean operation of the 
    --                         given type will be performed;
    --                      c) Operation required.
    --          Steps: a) Fill myShapes, myRemoved maps; 
    --                 b) Rebuild edges and faces; 
    --                 c) Build images of the object; 
    --                 d) Build the result of the operation.
    --          Result: Result shape of the operation required.
     
uses 
    Shape from TopoDS,  
    Face from TopoDS,  
    ListOfShape from TopTools, 
    MapOfOrientedShape from BOPCol,  
    MapOfShape from BOPCol,  
    IndexedMapOfShape from BOPCol, 
    DataMapOfShapeListOfShape from BOPCol, 
    DataMapOfShapeShape from BOPCol,  
    BaseAllocator from BOPCol,
    ListOfShape from BOPCol,
    BOP from BOPAlgo
     
is 
    Create 
      returns Builder from BRepFeat;  
    ---C++: alias "Standard_EXPORT virtual ~BRepFeat_Builder();"
 
    Clear(me:out) 
      is redefined;
    ---Purpose:  Clears internal fields and arguments.
 
    Init(me:out; 
        theShape : Shape from TopoDS); 
    ---Purpose: Initialyzes the object of local boolean operation.
    --          
 
    Init(me:out; 
        theShape : Shape from TopoDS; 
        theTool  : Shape from TopoDS);
    ---Purpose: Initialyzes the arguments of local boolean operation.
    --          
  
    SetOperation(me:out; 
        theFuse : Integer from Standard);
    ---Purpose: Sets the operation of local boolean operation.  
    --          If theFuse = 0 than the operation is CUT, otherwise FUSE.
 
    SetOperation(me:out; 
        theFuse : Integer from Standard;
        theFlag : Boolean from Standard);
    ---Purpose: Sets the operation of local boolean operation.
    --          If theFlag = TRUE it means that no selection of parts 
    --          of the tool is needed, t.e. no second part. In that case 
    --          if theFuse = 0 than operation is COMMON, otherwise CUT21. 
    --          If theFlag = FALSE SetOperation(theFuse) function  is called.
    
    Prepare(me:out) 
    is redefined protected;   
    ---Purpose: Prepares builder of local operation.
    --          
    
    PartsOfTool(me:out; 
        theLT  :  out ListOfShape from TopTools); 
    ---Purpose: Collects parts of the tool.
     
    KeepParts(me:out;
        theIm : ListOfShape from TopTools);
    ---Purpose: Initialyzes parts of the tool for second step of algorithm.
    --          Collects shapes and all sub-shapes into myShapes map.
 
    KeepPart(me:out;
        theS : Shape from TopoDS);
    ---Purpose: Adds shape theS and all its sub-shapes into myShapes map.
    --          
 
    PerformResult(me:out);
    ---Purpose: Main function to build the result of the 
    --          local operation required.
    
    RebuildFaces(me:out); 
    ---Purpose: Rebuilds faces in accordance with the kept parts of the tool.
    --          
     
    RebuildEdge(me:out; 
        theE:Shape from TopoDS; 
        theF:Face from TopoDS; 
        theME:MapOfShape from BOPCol; 
        aLEIm:out ListOfShape from BOPCol); 
    ---Purpose: Rebuilds edges in accordance with the kept parts of the tool.
    --          
    
    CheckSolidImages(me:out);
    ---Purpose: Collects the images of the object, that contains in 
    --          the images of the tool.
        
    FillRemoved(me:out); 
    ---Purpose: Collects the removed parts of the tool into myRemoved map.
    --          
    
    FillRemoved(me:out; 
        theS : Shape from TopoDS;
        theM : in out MapOfShape from BOPCol);  
    ---Purpose: Adds the shape S and its sub-shapes into myRemoved map.
    --          
         
    FillIn3DParts(me:out; 
        theInParts:out DataMapOfShapeListOfShape from BOPCol; 
        theDraftSolids:out DataMapOfShapeShape from BOPCol; 
        theAllocator:BaseAllocator from BOPCol)  
    is redefined protected;   
    ---Purpose: Function is redefined to avoid the usage of removed faces.
    --          

fields 
    myShapes : MapOfShape from BOPCol is protected;
    myRemoved : MapOfShape from BOPCol is protected; 
    myFuse : Integer from Standard is protected; 
 
end Builder;
