-- Created on: 1993-08-10
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PointOnCurve from BRep inherits PointRepresentation from BRep

	---Purpose: 

uses
    Curve    from Geom,
    Location from TopLoc
    
is

    Create(P : Real;
    	   C : Curve    from Geom;
	   L : Location from TopLoc)
    returns mutable PointOnCurve from BRep;
    
    
    IsPointOnCurve(me)          returns Boolean
	---Purpose: Returns True
    is redefined;
	
    IsPointOnCurve(me; C : Curve    from Geom;
    	    	       L : Location from TopLoc)   returns Boolean
    is redefined;
	

    Curve(me) returns any Curve from Geom
	---C++: return const &
    is redefined;
	
    Curve(me : mutable; C : Curve from Geom)
    is redefined;
	

fields
    
    myCurve : Curve from Geom;

end PointOnCurve;
