-- File:        FacetedBrepAndBrepWithVoids.cdl
-- Created:     Fri Jun 17 11:43:49 1994
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class FacetedBrepAndBrepWithVoids from StepShape 

inherits ManifoldSolidBrep from StepShape 


	--- This class is an implementation of EXPRESS
	--  ANDOR Subtype Declaration.
uses

	FacetedBrep from StepShape, 
	BrepWithVoids from StepShape, 
	ClosedShell from StepShape, 
	HArray1OfOrientedClosedShell from StepShape, 
	OrientedClosedShell from StepShape,
	HAsciiString from TCollection
is

	Create returns mutable FacetedBrepAndBrepWithVoids;
	---Purpose: Returns a FacetedBrepAndBrepWithVoids


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aOuter : mutable ClosedShell from StepShape) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aOuter : mutable ClosedShell from StepShape;
	      aFacetedBrep : mutable FacetedBrep from StepShape;
	      aBrepWithVoids : mutable BrepWithVoids from StepShape);

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aOuter : mutable ClosedShell from StepShape;
	      aVoids : mutable HArray1OfOrientedClosedShell from StepShape);

	-- Specific Methods for Field Data Access --

	SetFacetedBrep(me : mutable; aFacetedBrep : mutable FacetedBrep);
	FacetedBrep (me) returns mutable FacetedBrep;
	SetBrepWithVoids(me : mutable; aBrepWithVoids : mutable BrepWithVoids);
	BrepWithVoids (me) returns mutable BrepWithVoids;

	-- Specific Methods for ANDOR Field Data Access --

	SetVoids(me : mutable; aVoids : mutable HArray1OfOrientedClosedShell);
	Voids (me) returns mutable HArray1OfOrientedClosedShell;
	VoidsValue (me; num : Integer) returns mutable OrientedClosedShell;
	NbVoids (me) returns Integer;

	-- Specific Methods for ANDOR Field Data Access --


fields

	facetedBrep : FacetedBrep from StepShape;
	brepWithVoids : BrepWithVoids from StepShape;

end FacetedBrepAndBrepWithVoids;
