-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class RectangularTrimmedSurface from StepGeom 

inherits BoundedSurface from StepGeom 

uses

	Surface from StepGeom, 
	Real from Standard, 
	Boolean from Standard, 
	HAsciiString from TCollection
is

	Create returns mutable RectangularTrimmedSurface;
	---Purpose: Returns a RectangularTrimmedSurface


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aBasisSurface : mutable Surface from StepGeom;
	      aU1 : Real from Standard;
	      aU2 : Real from Standard;
	      aV1 : Real from Standard;
	      aV2 : Real from Standard;
	      aUsense : Boolean from Standard;
	      aVsense : Boolean from Standard) is virtual;

	-- Specific Methods for Field Data Access --

	SetBasisSurface(me : mutable; aBasisSurface : mutable Surface);
	BasisSurface (me) returns mutable Surface;
	SetU1(me : mutable; aU1 : Real);
	U1 (me) returns Real;
	SetU2(me : mutable; aU2 : Real);
	U2 (me) returns Real;
	SetV1(me : mutable; aV1 : Real);
	V1 (me) returns Real;
	SetV2(me : mutable; aV2 : Real);
	V2 (me) returns Real;
	SetUsense(me : mutable; aUsense : Boolean);
	Usense (me) returns Boolean;
	SetVsense(me : mutable; aVsense : Boolean);
	Vsense (me) returns Boolean;

fields

	basisSurface : Surface from StepGeom;
	u1 : Real from Standard;
	u2 : Real from Standard;
	v1 : Real from Standard;
	v2 : Real from Standard;
	usense : Boolean from Standard;
	vsense : Boolean from Standard;

end RectangularTrimmedSurface;
