-- Created on: 1991-04-04
-- Created by: Remi GILET
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package GccGeo


    ---Purpose :
    -- This package provides an implementation of analytic algorithms
    -- (using only non-persistant entities) used to create 2d lines or
    -- circles with geometric constraints.

uses GccEnt,
     GccInt,
     IntCurve,
     GeomAbs,
     TColStd,
     Standard,
     StdFail,
     TColgp,
     gp

is

generic class CurvePGTool;

generic class ParGenCurve;

generic class Circ2dTanCen;
    -- Create a 2d circle TANgent to a 2d entity and CENtered on a 2d point.

generic class Circ2d2TanRad;
    -- Create a 2d circle TANgent to 2 2d entities with the given RADius.

generic class Circ2dTanOnRad;
    -- Create a 2d circle TANgent to a 2d entity and centered ON a 2d 
    -- entity (not a point) with the given radius.

generic class Circ2d2TanOn;
    -- Create a 2d circle TANgent to 2 2d entities (circle, line or point) 
    -- and centered ON a 2d curve.

end GccGeo;
