-- File:	StepData_DescrProtocol.cdl
-- Created:	Wed May 21 15:00:44 1997
-- Author:	Christian CAILLET
--		<cky@heliox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1997


class DescrProtocol  from StepData    inherits FileProtocol  from StepData

    ---Purpose : A DescrProtocol is a protocol dynamically (at execution time)
    --           defined with :
    --           - a list of resources (inherits FileProtocol)
    --           - a list of entity descriptions
    --           i.e. it can be defined with only C++ writing to initialize it
    --           Its initialization must :
    --           - set its schema name
    --           - define its resources (which can also be other DescrProtocol)
    --           - define its entity descriptions
    --           - record it in the system by calling RecordLib

uses CString, AsciiString from TCollection

is

    Create returns mutable DescrProtocol;

    SetSchemaName (me : mutable; name : CString);
    ---Purpose : Defines a specific Schema Name for this Protocol

    LibRecord     (me);
    ---Purpose : Records this Protocol in the service libraries, with a
    --           DescrGeneral and a DescrReadWrite
    --           Does nothing if the Protocol brings no proper description

    SchemaName (me) returns CString  is redefined;
    ---Purpose : Returns the Schema Name attached to each class of Protocol
    --           here, returns the SchemaName set by SetSchemaName
    -- was C++ : return const

fields

    thename : AsciiString;

end DescrProtocol;
