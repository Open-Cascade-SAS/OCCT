-- Created on: 2002-12-12
-- Created by: data exchange team
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class FeaShellMembraneBendingCouplingStiffness from StepFEA
inherits FeaMaterialPropertyRepresentationItem from StepFEA

    ---Purpose: Representation of STEP entity FeaShellMembraneBendingCouplingStiffness

uses
    HAsciiString from TCollection,
    SymmetricTensor42d from StepFEA

is
    Create returns FeaShellMembraneBendingCouplingStiffness from StepFEA;
	---Purpose: Empty constructor

    Init (me: mutable; aRepresentationItem_Name: HAsciiString from TCollection;
                       aFeaConstants: SymmetricTensor42d from StepFEA);
	---Purpose: Initialize all fields (own and inherited)

    FeaConstants (me) returns SymmetricTensor42d from StepFEA;
	---Purpose: Returns field FeaConstants
    SetFeaConstants (me: mutable; FeaConstants: SymmetricTensor42d from StepFEA);
	---Purpose: Set field FeaConstants

fields
    theFeaConstants: SymmetricTensor42d from StepFEA;

end FeaShellMembraneBendingCouplingStiffness;
