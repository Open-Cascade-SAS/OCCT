-- Created on: 1994-11-03
-- Created by: Marie Jose MARTZ
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Actor from IGESToBRep
    inherits ActorOfTransientProcess  from Transfer

    ---Purpose : This class performs the transfer of an Entity from
    --           IGESToBRep
    --           
    --           I.E. for each type of Entity, it invokes the appropriate Tool
    --           then returns the Binder which contains the Result

uses TransientProcess, Binder, InterfaceModel from Interface

is

    Create  returns mutable Actor from IGESToBRep;

    SetModel (me : mutable; model : InterfaceModel from Interface);
    
    SetContinuity (me : mutable; continuity : Integer from Standard = 0);
    ---Purpose   By default continuity = 0
    --           if continuity = 1 : try C1
    --           if continuity = 2 : try C2
    
    GetContinuity (me) returns Integer from Standard;
    ---Purpose : Return "thecontinuity"

    Recognize (me : mutable; start : Transient) returns Boolean  is redefined;

    Transfer (me : mutable; start : Transient; TP : mutable TransientProcess)
    	returns mutable Binder  is redefined;

    UsedTolerance (me) returns Real;
    ---Purpose : Returns the tolerance which was actually used, either from
    --           the file or from statics

fields

    themodel      : InterfaceModel from Interface;
    thecontinuity : Integer;
    theeps        : Real;

end Actor;
