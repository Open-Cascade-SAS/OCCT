-- Created on: 2002-12-15
-- Created by: data exchange team
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class RWSiUnitAndMassUnit from RWStepBasic

	---Purpose : Read & Write Module for SiUnitAndMassUnit

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     SiUnitAndMassUnit from StepBasic

is

	Create returns RWSiUnitAndMassUnit;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : SiUnitAndMassUnit from StepBasic);

	WriteStep (me; SW : in out StepWriter; ent : SiUnitAndMassUnit from StepBasic);

end RWSiUnitAndMassUnit;
