-- Created on: 1992-04-06
-- Created by: Christian CAILLET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class IGESReaderTool  from IGESData  inherits FileReaderTool

    ---Purpose : specific FileReaderTool for IGES
    --           Parameters are accessed through specific objects, ParamReaders

uses Integer, Boolean,  Transient,
     Check,  InterfaceModel, GeneralLib,  ReaderLib,  ParamList,
     IGESReaderData,  Protocol from IGESData, FileRecognizer,
     IGESType,        IGESEntity,   DirPart,  ReadStage,   ParamReader

is

    Create (reader : IGESReaderData; protocol : Protocol from IGESData)
    	returns IGESReaderTool;
    ---Purpose : creates IGESReaderTool to work with an IGESReaderData and an
    --           IGES Protocol.
    --           Actually, no Lib is used

    	-- --   General   -- --

    Prepare (me : in out; reco : FileRecognizer);
    ---Purpose : binds empty entities to records, works with the Protocol
    --           (from IGESData) stored and later used
    --           RQ : Actually, sets DNum into IGES Entities
    --           Also loads the list of parameters for ParamReader

    Recognize (me : in out; num : Integer;
    	       ach : in out Check; ent : out Transient)
    	returns Boolean;
    ---Purpose : recognizes records by asking Protocol (on data of DirType)

    	--    Loading the IGESModel    --

    BeginRead (me : in out; amodel : InterfaceModel);
    ---Purpose : fills model's header, that is, its GlobalSection

    AnalyseRecord (me : in out;
    	num : Integer; anent : Transient; acheck : in out Check)
	    returns Boolean;
    ---Purpose : fills an entity, given record no; works by calling ReadDirPart
    --           then ReadParams (with help of a ParamReader), then if required
    --           ReadProps and ReadAssocs, from IGESEntity
    --           Returns True if no fail has been recorded

    EndRead (me : in out; amodel : InterfaceModel) is redefined;
    ---Purpose : after reading entities, true line weights can be computed

    	--    For each IGESEntity    --

    ReadDir       (me; ent : IGESEntity; IR : IGESReaderData;
    	           DP : DirPart; ach : in out Check);
    ---Purpose : Reads directory part componants from file; DP is the litteral
    --           directory part, IR detains entities referenced by DP

    ReadOwnParams (me; ent : IGESEntity;
    	    	   IR : IGESReaderData; PR : in out ParamReader);
    ---Purpose : Performs Reading of own Parameters for each IGESEntity
    --           Works with the ReaderLib loaded with ReadWriteModules for IGES
    --           In case of failure, tries UndefinedEntity from IGES

    ReadProps     (me; ent : IGESEntity; IR : IGESReaderData;
    	    	   PR : in out ParamReader);
    ---Purpose : Reads Property List, if there is (if not, does nothing)
    --           criterium is : current parameter of PR remains inside params
    --           list, and Stage is "Own"
    --           Current parameter must be a positive integer, which value
    --           gives the length of the list; else, a Fail is produced (into
    --           Check of PR) and reading process is stopped

    ReadAssocs    (me; ent : IGESEntity; IR : IGESReaderData;
    	    	   PR : in out ParamReader);
    ---Purpose : Reads Associativity List, if there is (if not, does nothing)
    --           criterium is : current parameter of PR remains inside params
    --           list, and Stage is "Own"
    --           Same conditions as above; in addition, no parameter must be
    --           let after the list once read
    --           Note that "Associated" entities are not declared "Shared"

fields

    thelist : ParamList;         -- (loaded once, allows optimization)
    thereco : FileRecognizer;
    theglib : GeneralLib;
    therlib : ReaderLib;
    thecnum : Integer;           -- current entity number for recognize
    thectyp : IGESType;          -- its IGESType (for purpose of optimization)
    thestep : ReadStage;         -- to continue an interrupted party
    thechk  : Check;             -- check on header (kept by IGESModel)
    thegradweight : Integer;
    themaxweight  : Real;
    thedefweight  : Real;

end IGESReaderTool;
