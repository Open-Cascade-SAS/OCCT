-- Created on: 2002-04-18
-- Created by: Michael KLOKOV
-- Copyright (c) 2002-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class TopolTool from IntTools inherits TopolTool from Adaptor3d

    	---Purpose: Class redefine methods of TopolTool from Adaptor3d
	---         concerning sample points
	---
uses
    Pnt   from gp,
    Pnt2d from gp,
    HSurface from Adaptor3d, 
    HArray1OfReal  from  TColStd

raises DomainError from Standard

is
    Create returns mutable TopolTool from IntTools;
    	---Purpose:
	--- Empty constructor
	---

    Create(theSurface: HSurface from Adaptor3d)
    	returns mutable TopolTool from IntTools;
	---Purpose:
	--- Initializes me by surface
	---

    Initialize(me: mutable)
    	is redefined;
	---Purpose:
	--- Redefined empty initializer
	---
	--  Warning:
	--- Raises the exception NotImplemented
	---
    
    Initialize(me: mutable; theSurface: HSurface from Adaptor3d)
	is redefined;
	---Purpose:
	--- Initializes me by surface
	---

    --- sample points  tools

    ComputeSamplePoints(me: mutable)
    	is redefined;
	---Purpose:
	--- 
	---
    
    NbSamplesU(me: mutable) 
    	returns Integer from Standard
    	is redefined;
    	---Purpose: 
    	--- Computes the sample-points for the intersections algorithms
	---
    
    NbSamplesV(me: mutable) 
    	returns Integer from Standard
    	is redefined;
    	---Purpose: 
    	--- Computes the sample-points for the intersections algorithms
	---
    
    NbSamples(me: mutable)
    	returns Integer from Standard
    	is redefined;
        ---Purpose: 
    	--- Computes the sample-points for the intersections algorithms
	---

    SamplePoint(me: mutable; Index: Integer from Standard;
                             P2d  : out Pnt2d   from gp;
                             P3d  : out Pnt     from gp)
    	is redefined;
	---Purpose:
	--- Returns a 2d point from surface myS
	--- and a corresponded 3d point
	--- for given index.
	--- The index should be from 1 to NbSamples()
	---

    --modified by NIZNHY-IFV Sep 28 16:01:38 2005 f
    SamplePnts(me: mutable; theDefl:  Real  from  Standard; theNUmin, theNVmin: Integer from Standard)
        ---Purpose: compute the sample-points for the intersections algorithms
	-- by adaptive algorithm for BSpline surfaces. For other surfaces algorithm
	-- is the same as in method ComputeSamplePoints(), but only fill arrays of U
	-- and V sample parameters;
	-- theDefl is a requred deflection
	-- theNUmin, theNVmin are minimal nb points for U and V.
    is redefined;
    
fields
    --myS         : HSurface from Adaptor3d;  now inherits myS from Adaptor3d_TopolTool
    myNbSmplU   : Integer  from Standard;
    myNbSmplV   : Integer  from Standard;
    myU0        : Real     from Standard;
    myV0        : Real     from Standard;
    myDU        : Real     from Standard;
    myDV        : Real     from Standard;
     
end TopolTool from IntTools;
