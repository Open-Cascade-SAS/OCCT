-- Created on: 1993-04-15
-- Created by: Philippe DAUTRY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package TColGeom2d


        ---Purpose : 
-- The package TColGeom2d provides standard and
-- frequently used instantiations of generic classes from
-- the TCollection package with geometric objects from the Geom2d package.

uses TCollection, Geom2d

is


    class Array1OfGeometry 
    	instantiates Array1 from TCollection (Geometry from Geom2d);
    class Array1OfCurve 
    	instantiates Array1 from TCollection (Curve from Geom2d);
    class Array1OfBoundedCurve 
    	instantiates Array1 from TCollection (BoundedCurve from Geom2d);
    class Array1OfBezierCurve 
    	instantiates Array1 from TCollection (BezierCurve from Geom2d);
    class Array1OfBSplineCurve 
    	instantiates Array1 from TCollection (BSplineCurve from Geom2d);

    class HArray1OfGeometry
    	instantiates HArray1 from TCollection (Geometry from Geom2d,
    	    	    	    	Array1OfGeometry from TColGeom2d);
    class HArray1OfCurve
    	instantiates HArray1 from TCollection (Curve from Geom2d,
    	    	    	    	Array1OfCurve from TColGeom2d);
    class HArray1OfBoundedCurve 
    	instantiates HArray1 from TCollection (BoundedCurve from Geom2d,
    	    	    	    	Array1OfBoundedCurve from TColGeom2d);
    class HArray1OfBezierCurve  
    	instantiates HArray1 from TCollection (BezierCurve from Geom2d,
    	    	    	    	Array1OfBezierCurve from TColGeom2d);
    class HArray1OfBSplineCurve 
    	instantiates HArray1 from TCollection (BSplineCurve from Geom2d,
    	    	    	    	Array1OfBSplineCurve from TColGeom2d);


    class SequenceOfGeometry  
    	instantiates Sequence from TCollection (Geometry from Geom2d);
    class SequenceOfCurve  
    	instantiates Sequence from TCollection (Curve from Geom2d);
    class SequenceOfBoundedCurve  
    	instantiates Sequence from TCollection (BoundedCurve from Geom2d);

    class HSequenceOfGeometry  
    	instantiates HSequence from TCollection (Geometry from Geom2d,
    	    	    	    	SequenceOfGeometry from TColGeom2d);
    class HSequenceOfCurve  
    	instantiates HSequence from TCollection (Curve from Geom2d,
    	    	    	    	SequenceOfCurve from TColGeom2d);
    class HSequenceOfBoundedCurve  
    	instantiates HSequence from TCollection (BoundedCurve from Geom2d,
    	    	    	    	SequenceOfBoundedCurve from TColGeom2d);


end TColGeom2d;
