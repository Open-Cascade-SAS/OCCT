-- Created on: 1994-11-14
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Pave from TopOpeBRepBuild 
    inherits Loop from TopOpeBRepBuild

uses
    
    ShapeEnum from TopAbs,
    Shape from TopoDS, 
    --modified by NIZHNY-MZV  Mon Feb 21 14:29:26 2000
    Kind  from  TopOpeBRepDS
is

    Create(V : Shape from TopoDS; P : Real; bound : Boolean) returns mutable Pave;
    ---Purpose: V = vertex, P = parameter of vertex <V>
    --          bound = True if <V> is an old vertex
    --          bound = False if <V> is a new vertex
    
    HasSameDomain(me : mutable; b : Boolean);
    SameDomain(me : mutable; VSD : Shape from TopoDS);

    HasSameDomain(me) returns Boolean from Standard;
    SameDomain(me) returns Shape from TopoDS;
    ---C++: return const &

    Vertex(me) returns Shape from TopoDS is static;
    ---C++: return const &

    ChangeVertex(me : mutable) returns Shape from TopoDS is static;
    ---C++: return &
    -- used only by PaveSet
    Parameter(me) returns Real from Standard is static;
 
    --modified by NIZHNY-MZV  Mon Feb 21 14:09:47 2000 
    Parameter(me:  mutable;  Par:  Real  from  Standard)  is static;
    --modified by NIZHNY-MZV  Mon Feb 21 14:25:58 2000 
    InterferenceType(me:  mutable)  returns  Kind  from  TopOpeBRepDS; 
    ---C++: return &
	  
    IsShape(me) returns Boolean from Standard is redefined;
    Shape(me) returns Shape from TopoDS is redefined;
    ---C++: return const &

    Dump(me) is redefined;
    
fields

    myVertex  : Shape from TopoDS;
    myParam   : Real from Standard;
    myIsShape : Boolean from Standard;
    myHasSameDomain : Boolean from Standard;
    mySameDomain : Shape from TopoDS;

    --modified by NIZHNY-MZV  Mon Feb 21 14:26:58 2000 
    myIntType  :  Kind  from  TopOpeBRepDS; 

end Pave from TopOpeBRepBuild;
