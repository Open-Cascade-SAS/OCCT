-- Created on: 1997-02-12
-- Created by: Alexander BRIVIN
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class MatrixTransform from Vrml 

	---Purpose: defines a MatrixTransform node of VRML specifying matrix and transform
	--          properties. 
    	--  This  node  defines  3D  transformation  with  a  4  by  4  matrix.
    	--  By  default  :   
    	--  a11=1  a12=0  a13=0  a14=0
    	--  a21=0  a22=1  a23=0  a24=0
    	--  a31=0  a32=0  a33=1  a34=0
    	--  a41=0  a42=0  a43=0  a44=1	
	--  It  is  written  to  the  file  in  row-major  order  as  16  Real numbers 
	--  separated  by  whitespace.  For  example ,  matrix  expressing  a  translation 
	--  of  7.3  units  along  the  X  axis  is  written  as: 
	--  1  0  0  0   0  1  0  0   0  0  1  0   7.3 0  0  1
uses
 
   Trsf   from   gp

is
 
    Create returns  MatrixTransform from Vrml;
 
    Create  ( aMatrix  :  Trsf    from  gp )
        returns  MatrixTransform from Vrml;
   
    SetMatrix ( me : in out;  aMatrix  :  Trsf    from  gp );
    Matrix ( me )  returns  Trsf    from  gp;

    Print  ( me;  anOStream: in out OStream from Standard) returns OStream from Standard;
    ---C++:  return  & 

fields
 
    myMatrix  :  Trsf    from  gp; -- Transformation matrix

end MatrixTransform;

