-- Created on: 1995-02-07
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class LineConstructor from GeomInt

        ---Purpose: Splits given Line.

uses Line           from IntPatch,
     TopolTool      from Adaptor3d,
     HSurface        from GeomAdaptor,
     SequenceOfReal from TColStd

raises NotDone    from StdFail,
       OutOfRange from Standard

is

    Create
    	returns LineConstructor from GeomInt;
        ---C++: inline
	---Purpose: 
	--- Empty constructor
	---

    Load(me: in out; D1,D2: TopolTool from Adaptor3d;
                     S1,S2: HSurface  from GeomAdaptor)
    	is static;
        ---C++: inline
	---Purpose:
	--- Initializes me by two surfaces and corresponding
	--- tools which represent boundaries of surfaces
	---

    Perform(me: in out; L: Line from IntPatch)
    	is static;
	---Purpose:
	--- Splits line
	---

    IsDone(me)
    	returns Boolean from Standard
	is static;
	---C++: inline
	---Purpose:
	--- Returns True if splitting was successful
	---

    NbParts(me)
    	returns Integer from Standard
	raises NotDone from StdFail
	is static;
	---C++: inline
	---Purpose:
	--- Returns number of splits
	---

    Part(me; I: Integer from Standard; WFirst,WLast: out Real from Standard) 
    	raises NotDone    from StdFail,
               OutOfRange from Standard
	is static;
	---C++: inline
	---Purpose:
	--- Return first and last parameters 
    	--- for given index of split
	---

    PeriodicLine(me; L: Line from IntPatch)
    	is static private;

fields

    done  : Boolean        from Standard;
    seqp  : SequenceOfReal from TColStd;
    myDom1: TopolTool      from Adaptor3d;
    myDom2: TopolTool      from Adaptor3d;
    myHS1 : HSurface       from GeomAdaptor;
    myHS2 : HSurface       from GeomAdaptor;

end LineConstructor;
