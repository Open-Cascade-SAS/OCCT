-- Created on: 1991-07-19
-- Created by: Isabelle GRIGNON
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

private class MyGaussFunction from CPnts 
inherits Function from math

uses
    RealFunction from CPnts

is

    Create returns MyGaussFunction;
	---C++: inline

    Init(me : in out;
    	   F : RealFunction from CPnts;
           D : Address from Standard);
	---Purpose: F  is a pointer on a  function  D is a client data
	--          
	--          Each value is computed with F(D)
    
    Value(me: in out; X : Real; F : out Real)
    returns Boolean
    is static;

fields

    myFunction : RealFunction from CPnts;
    myData     : Address      from Standard;

end MyGaussFunction;
