-- Created on: 1993-12-13
-- Created by: Christophe MARION
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class   ExtPElC2d from Extrema 
    	---Purpose: It calculates all the distances between a point
    	--          and an elementary curve.
    	--          These distances can be minimum or maximum.

uses    POnCurv2d from Extrema,
        Lin2d     from gp,
    	Circ2d    from gp,
    	Elips2d   from gp,
    	Hypr2d    from gp,
    	Parab2d   from gp,
    	Pnt2d     from gp

raises  NotDone     from StdFail,
    	OutOfRange  from Standard

is
    Create returns ExtPElC2d;

    Create (P: Pnt2d; C: Lin2d; Tol: Real;
            Uinf: Real; Usup: Real)
    	returns ExtPElC2d;
    	---Purpose: Calculates the extremum distance between the
    	--          point P and the segment [Uinf,Usup] of the line L.


    Perform(me: in out; P: Pnt2d; L: Lin2d; Tol: Real; Uinf,Usup: Real)
    is static;

    Create (P: Pnt2d; C: Circ2d; Tol: Real;
            Uinf: Real; Usup: Real)
    	returns ExtPElC2d;
    	---Purpose: Calculates the 2 extremum distances between the
    	--          point P and the segment [Uinf,Usup] of the circle C.
    	--          Tol is used to determine
    	--          if P is on the axis of the circle or
    	--          if an extremum is on an endpoint of the segment.
    	--          If P is on the axis of the circle,
    	--          there are infinite solution then IsDone(me)=False.
    	--          The conditions on the Uinf and Usup are:
    	--            0. <= Uinf <= 2.*PI and Usup > Uinf.
    	--          If Usup > Uinf + 2.*PI, then only the solutions in
    	--          the range [Uinf,Uinf+2.*PI[ are computed.


    Perform(me: in out; P: Pnt2d; C: Circ2d; Tol: Real; Uinf,Usup: Real)
    is static;

    Create (P: Pnt2d; C: Elips2d; Tol: Real;
            Uinf: Real; Usup: Real)
    returns ExtPElC2d;
    	---Purpose: Calculates the 4 extremum distances between the
    	--          point P and the segment [Uinf,Usup] of the elipse C.
     	--          Tol is used to determine
     	--          if the point is on the axis of the elipse and
     	--          if the major radius is equal to the minor radius or
     	--          if an extremum is on an endpoint of the segment.
    	--          If P is on the axis of the elipse,
    	--          there are infinite solution then IsDone(me)=False.
    	--          The conditions on the Uinf and Usup are:
    	--            0. <= Uinf <= 2.*PI and Usup > Uinf.
    	--          If Usup > Uinf + 2.*PI, then only the solutions in
    	--          the range [Uinf,Uinf+2.*PI[ are computed.


    Perform(me: in out; P: Pnt2d; C: Elips2d; Tol: Real; Uinf,Usup: Real)
    is static;

    Create (P: Pnt2d; C: Hypr2d; Tol: Real; Uinf: Real;
            Usup: Real)
    returns ExtPElC2d;
    	---Purpose: Calculates the extremum distances between the
    	--          point P and the segment [Uinf,Usup] of the hyperbola
    	--          C.
    	--          Tol is used to determine if two solutions u and v
    	--          are identical; the condition is:
    	--          dist(C(u),C(v)) < Tol.

    Perform(me: in out; P: Pnt2d; C: Hypr2d; Tol: Real; Uinf,Usup: Real)
    is static;

    Create (P: Pnt2d; C: Parab2d; Tol: Real; Uinf: Real;
            Usup: Real)
    returns ExtPElC2d;
    	---Purpose: Calculates the 4 extremum distances between the
    	--          point P and the segment [Uinf,Usup] of the parabola
    	--          C.
    	--          Tol is used to determine if two solutions u and v
    	--          are identical; the condition is:
    	--          dist(C(u),C(v)) < Tol.

    Perform(me: in out; P: Pnt2d; C: Parab2d; Tol: Real; Uinf,Usup: Real)
    is static;
    

    IsDone (me) returns Boolean
    	---Purpose: True if the distances are found.
    	is static;

    NbExt (me) returns Integer
    	---Purpose: Returns the number of extremum distances.
	raises  NotDone from StdFail
	    	-- if IsDone(me)=False.
    	is static;
    
    SquareDistance (me; N: Integer) returns Real
    	---Purpose: Returns the value of the Nth extremum square distance.
    	raises  NotDone from StdFail,
	    	-- if IsDone(me)=False.
    	    	OutOfRange
	    	-- if N < 1 or N > NbPoints(me).
    	is static;

    IsMin (me; N: Integer) returns Boolean
    	---Purpose: Returns True if the Nth extremum distance is a
    	--          minimum.
    	raises  NotDone from StdFail,
	    	-- if IsDone(me)=False.
    	    	OutOfRange
	    	-- if N < 1 or N > NbPoints(me).
    	is static;

    Point (me; N: Integer) returns POnCurv2d
        ---C++: return const &
    	---Purpose: Returns the point of the Nth extremum distance.
    	raises  NotDone from StdFail,
	    	-- if IsDone(me)=False.
    	    	OutOfRange
	    	-- if N < 1 or N > NbPoints(me).
    	is static;

fields
    myDone : Boolean;
    myNbExt: Integer;
    mySqDist: Real [4];
    myIsMin: Boolean [4];
    myPoint: POnCurv2d from Extrema [4];

end ExtPElC2d;
