-- File:        FileName.cdl
-- Created:     Thu Jun 16 18:05:53 1994
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class FileName from HeaderSection 

inherits TShared from MMgt

uses

	HAsciiString from TCollection, 
	HArray1OfHAsciiString from Interface
is

	Create returns mutable FileName;
	---Purpose: Returns a FileName

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aTimeStamp : mutable HAsciiString from TCollection;
	      aAuthor : mutable HArray1OfHAsciiString from Interface;
	      aOrganization : mutable HArray1OfHAsciiString from Interface;
	      aPreprocessorVersion : mutable HAsciiString from TCollection;
	      aOriginatingSystem : mutable HAsciiString from TCollection;
	      aAuthorisation : mutable HAsciiString from TCollection);

	-- Specific Methods for Field Data Access --

	SetName(me : mutable; aName : mutable HAsciiString);
	Name (me) returns mutable HAsciiString;
	SetTimeStamp(me : mutable; aTimeStamp : mutable HAsciiString);
	TimeStamp (me) returns mutable HAsciiString;
	SetAuthor(me : mutable; aAuthor : mutable HArray1OfHAsciiString);
	Author (me) returns mutable HArray1OfHAsciiString;
	AuthorValue (me; num : Integer) returns mutable HAsciiString;
	NbAuthor (me) returns Integer;
	SetOrganization(me : mutable; aOrganization : mutable HArray1OfHAsciiString);
	Organization (me) returns mutable HArray1OfHAsciiString;
	OrganizationValue (me; num : Integer) returns mutable HAsciiString;
	NbOrganization (me) returns Integer;
	SetPreprocessorVersion(me : mutable; aPreprocessorVersion : mutable HAsciiString);
	PreprocessorVersion (me) returns mutable HAsciiString;
	SetOriginatingSystem(me : mutable; aOriginatingSystem : mutable HAsciiString);
	OriginatingSystem (me) returns mutable HAsciiString;
	SetAuthorisation(me : mutable; aAuthorisation : mutable HAsciiString);
	Authorisation (me) returns mutable HAsciiString;

fields

	name : HAsciiString from TCollection;
	timeStamp : HAsciiString from TCollection;
	author : HArray1OfHAsciiString from Interface;
	organization : HArray1OfHAsciiString from Interface;
	preprocessorVersion : HAsciiString from TCollection;
	originatingSystem : HAsciiString from TCollection;
	authorisation : HAsciiString from TCollection;

end FileName;
