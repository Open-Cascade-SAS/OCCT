-- Created on: 1992-11-05
-- Created by: Remi LEQUETTE
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Sphere from BRepPrim inherits Revolution from BRepPrim

	---Purpose: Implements the sphere primitive

uses
    Face from TopoDS,
    
    Pnt from gp,
    Ax2 from gp    

raises
    DomainError

is

    Create(Radius : Real)
    returns Sphere from BRepPrim
	---Purpose: Creates a Sphere at  origin with  Radius. The axes
	--          of the sphere are the  reference axes. An error is
	--          raised if the radius is < Resolution.
    raises DomainError;
    
    Create(Center : Pnt from gp; Radius : Real)
    returns Sphere from BRepPrim
	---Purpose: Creates a Sphere with Center and Radius.  Axes are
	--          the   referrence    axes.   This    is the    STEP
	--          constructor.
    raises DomainError;
    
    Create(Axes : Ax2 from gp; Radius : Real)
    returns Sphere from BRepPrim
	---Purpose: Creates a sphere with given axes system.
    raises DomainError;
    
    MakeEmptyLateralFace(me) returns Face from TopoDS
	---Purpose: The surface normal should be directed  towards the
	--          outside.
    is redefined;
    
    SetMeridian(me : in out)
    is static private;
    
fields
    myRadius : Real;

end Sphere;
