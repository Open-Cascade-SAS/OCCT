-- Created on: 1999-06-24
-- Created by: Sergey ZARITCHNY
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class CopyLabel from TDF 

	---Purpose: 

uses
 
    Boolean             from Standard,
    Label               from TDF,
    Attribute           from TDF,
    DataSet             from TDF,
    RelocationTable     from TDF,
    AttributeMap        from TDF,
    LabelMap            from TDF,
    IDFilter            from TDF


is
 
    Create  returns  CopyLabel  from TDF; 
    ---Purpose: Empty  constructor  
    
    Create(aSource,  aTarget  :  Label  from  TDF) 
      returns  CopyLabel  from TDF;  
    ---Purpose: CopyTool  
    
    Load(me  :  in  out;  aSource,  aTarget  :  Label  from  TDF);  
    ---Purpose: Loads  src  and  tgt  labels 
     
    UseFilter(me  :  in  out;  aFilter : IDFilter from TDF); 
    ---Purpose:  Sets  filter

    ExternalReferences(myclass;  Lab  :  Label  from  TDF; 
    	    	    	    	 aExternals:in  out  AttributeMap  from  TDF; 
    	    	    	    	 aFilter   :  IDFilter  from  TDF) 
      returns  Boolean  from  Standard; 
    ---Purpose: Check  external  references and  if  exist  fills  the  aExternals  Map 
     
    ExternalReferences(myclass;  aRefLab, Lab  :  Label  from  TDF; 
    	    	    	   aExternals    :  in  out  AttributeMap  from  TDF; 
			   aFilter       :  IDFilter  from  TDF;
    	    	    	   aDataSet      :  in  out  DataSet  from  TDF) ;
    ---Purpose: Check  external  references and  if  exist  fills  the  aExternals  Map 
     
    Perform(me:in  out);  
    ---Purpose:  performs  algorithm  of  selfcontained  copy 
     
    IsDone(me) 
      returns  Boolean  from  Standard;  
    ---C++:  inline      
	 
    RelocationTable(me)     	 
      returns  RelocationTable  from  TDF;  
    ---Purpose: returns  relocation  table 
    ---C++: return const&
    
fields
 
    myRT        :  RelocationTable  from  TDF;
    mySL        :  Label            from  TDF; --  source  label
    myTL        :  Label            from  TDF; --  target  label 
    myFilter    :  IDFilter         from  TDF;
    myMapOfExt  :  AttributeMap     from  TDF; --  map  of  attribute  with  external  reference
    myIsDone    :  Boolean          from  Standard;

end CopyLabel;
