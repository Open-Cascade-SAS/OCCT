-- Created on: 1992-04-07
-- Created by: Christian CAILLET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class LevelListEntity  from IGESData  inherits IGESEntity

    ---Purpose : defines required type for LevelList in directory part
    --           an effective LevelList entity must inherits it

uses Boolean, Integer

raises OutOfRange

is

    NbLevelNumbers (me) returns Integer  is deferred;
    ---Purpose : Must return the count of levels

    LevelNumber (me; num : Integer) returns Integer
        raises OutOfRange  is deferred;
    ---Purpose : returns the Level Number of <me>, indicated by <num>
    -- raises an exception if num is out of range

    HasLevelNumber (me; level : Integer) returns Boolean;
    ---Purpose : returns True if <level> is in the list

end LevelListEntity;
