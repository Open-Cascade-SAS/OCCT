-- Created on: 1992-02-17
-- Created by: Christian CAILLET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



generic class SimpleBinder  from Transfer

    	  (TheResult as any;  -- any : avoid Transient classes
	   TheInfo   as any)  -- template : DataInfo

        inherits Binder

    ---Purpose : Allows direct binding between a starting Object and the Result
    --           of its transfer when it is Unique.
    --           The Result itself is defined as a formal parameter <TheResult>           
    --  Warning : While it is possible to instantiate SimpleBinder with any Type
    --           for the Result, it is not advisable to instantiate it with
    --           Transient Classes, because such Results are directly known and
    --           managed by TransferProcess & Co, through
    --           SimpleBinderOfTransient : this class looks like instantiation
    --           of SimpleBinder, but its method ResultType
    --           is adapted (reads DynamicType of the Result)

uses CString, Type

raises TransferFailure

is

    Create returns mutable SimpleBinder;
    ---Purpose : normal standard constructor, creates an empty SimpleBinder

    Create (res : any TheResult) returns mutable SimpleBinder;
    ---Purpose : constructor which in the same time defines the result

--    IsMultiple (me) returns Boolean;
    ---Purpose : Returns True if a starting object is bound with SEVERAL
    --           results : Here, returns allways False
    --           But it can have next results

    ResultType (me) returns Type;
    ---Purpose : Returns the Type permitted for the Result, i.e. the Type
    --           of the Parameter Class <TheResult> (statically defined)

    ResultTypeName (me) returns CString;
    ---Purpose : Returns the Type Name computed for the Result (dynamic)

    SetResult (me : mutable; res : any TheResult)
    ---Purpose : Defines the Result
    	raises TransferFailure;
    --           Error if the Result is already used (see class Binder)

    Result (me) returns any TheResult
    ---Purpose : Returns the defined Result, if there is one
    	raises TransferFailure;
    --           Error if the Result is not defined (see class Binder)
    ---C++ : return const &

    CResult (me : mutable) returns any TheResult;
    ---Purpose : Returns the defined Result, if there is one, and allows to
    --           change it (avoids Result + SetResult).
    --           Admits that Result can be not yet defined
    --  Warning : a call to CResult causes Result to be known as defined
    ---C++ : return &

fields

    theres : TheResult;

end SimpleBinder;
