-- Created on: 1992-09-23
-- Created by: Christian CAILLET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Cycles  from IFGraph  inherits SubPartsIterator

    	---Purpose : determines strong componants in a graph which are Cycles

uses Graph, StrongComponants

is

    Create (agraph : Graph; whole : Boolean) returns Cycles;
    ---Purpose : creates with a Graph, and will analyse :
    --           whole True  : all the contents of the Model
    --           whole False : sub-parts which will be given later

    Create (subparts : in out StrongComponants);
    ---Purpose : creates from a StrongComponants which was already computed

    Evaluate (me : in out) is redefined;
    ---Purpose : does the computation. Cycles are StrongComponants which are
    --           not Single

    	-- --   Iteration : More-Next-etc... will give Cycles

end Cycles;
