-- Created on: 1998-07-17
-- Created by: Jean-Louis Frenkel
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

private class Timer from CDF
uses Timer from OSD
is
    Create returns Timer from CDF;

     
    ShowAndRestart(me: in out; aMessage: CString from Standard);
    
    ShowAndStop(me: in out; aMessage: CString from Standard);
   

    Show(me: in out; aMessage: CString from Standard)
    is private;

    MustShow(me: in out)  returns Boolean from Standard;
    
fields
    myTimer: Timer from OSD;
end Timer from OSD;
