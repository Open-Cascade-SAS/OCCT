-- Created on: 2000-09-08
-- Created by: data exchange team
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Centroid from XCAFDoc inherits Attribute from TDF

	---Purpose: attribute to store centroid

uses
    Pnt from gp,
    Label from TDF,
    RelocationTable from TDF
    
is
    Create returns Centroid from XCAFDoc;
  	---Purpose: class methods
    	--          =============

    GetID (myclass)   
    	---C++: return const &  
    returns GUID from Standard;

    Set (myclass; label : Label from TDF; pnt : Pnt from gp)
    	---Purpose: Find, or create, a Location attribute and set it's value
    	--          the Location attribute is returned.
    returns Centroid from XCAFDoc;

    	---Purpose: Location methods
    	--          ===============
    
    Set (me : mutable; pnt : Pnt from gp);
    
    Get (me)
    returns Pnt from gp;

    Get (myclass ; label : Label from TDF; pnt: in out Pnt from gp)
    returns Boolean from Standard;
        ---Purpose: Returns point as argument
	--          returns false if no such attribute at the <label>

    	---Category: methodes de TDF_Attribute
    	--           =========================
    
    ID (me)
    	---C++: return const & 
    returns GUID from Standard;

    Restore (me: mutable; With : Attribute from TDF);

    NewEmpty (me)
    returns Attribute from TDF;

    Paste (me; Into : Attribute from TDF;
	       RT   : RelocationTable from TDF);    

    Dump(me; anOS : in out OStream from Standard)
    	returns OStream from Standard
    	is redefined;
	---C++: return &

fields

    myCentroid : Pnt from gp;
    
end Centroid;
