-- Created on: 2000-08-16
-- Created by: data exchange team
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Color from XCAFDoc inherits     Attribute from TDF

	---Purpose: attribute to store color

uses
    Color from Quantity,
    NameOfColor from Quantity,
    Label from TDF,
    RelocationTable from TDF

is
    Create returns Color from XCAFDoc;
    
    ---Category: class methods
    --           =============

    GetID (myclass)   
    	---C++: return const &  
    returns GUID from Standard;
    
    
    Set (myclass; label : Label from TDF; C : Color from Quantity)
    returns Color from XCAFDoc;

    Set (myclass; label : Label from TDF; C : NameOfColor from Quantity)
    returns Color from XCAFDoc;

    Set (myclass; label : Label from TDF; R,G,B : Real from Standard)
    returns Color from XCAFDoc;

    ---Purpose: Find, or create, a Color attribute and set it's value
    --          the Color attribute is returned.

    
    
    ---Category: Color methods
    --           ===============
    
    Set (me : mutable;  C : Color from Quantity);
	     
    Set (me : mutable;  C : NameOfColor from Quantity);
	     
    Set (me : mutable;  R,G,B : Real from Standard);
		    
    GetColor (me) returns Color from Quantity;
        ---C++: return const & 

    GetNOC (me) returns NameOfColor from Quantity;
	     
    GetRGB (me;  R,G,B : out Real from Standard);
    
    --IsCaptured(me) returns Boolean;
	---Purpose: Returns True if there is a reference on the same label

    ---Category: methodes de TDF_Attribute
    --           =========================
    
    ID (me)
    	---C++: return const & 
    returns GUID from Standard;

    Restore (me: mutable; With : Attribute from TDF);

    NewEmpty (me)
    returns Attribute from TDF;

    Paste (me; Into : Attribute from TDF;
	       RT   : RelocationTable from TDF);    

--    Dump(me; anOS : in out OStream from Standard)
--    	returns OStream from Standard
--    	is redefined;
--	-C++: return &

fields
    myColor   : Color from Quantity;
    
end Color;
