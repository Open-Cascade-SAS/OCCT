-- File:	XDEDRAW_Layers.cdl
-- Created:	Fri Aug  4 14:39:39 2000
-- Author:	Pavel TELKOV
--		<ptv@zamox.nnov.matra-dtv.fr>
---Copyright:	 Matra Datavision 2000

class Layers from XDEDRAW 

    ---Purpose: Contains commands to work with layers

uses
    Interpretor from Draw
    
is

    InitCommands (myclass; theCommands: in out Interpretor from Draw);
	
end Layers;
