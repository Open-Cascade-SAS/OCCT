-- Created on: 1993-08-10
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PointOnCurveOnSurface from BRep inherits  PointsOnSurface from  BRep

uses

    Curve    from Geom2d,
    Surface  from Geom,
    Location from TopLoc

is

    Create(P : Real;
    	   C : Curve from Geom2d;
	   S : Surface from Geom;
	   L : Location from TopLoc)
    returns PointOnCurveOnSurface from BRep;
    
    IsPointOnCurveOnSurface(me) returns Boolean
	---Purpose: Returns True
    is redefined;

    IsPointOnCurveOnSurface(me; PC : Curve     from Geom2d;
    	    	    	    	S  : Surface  from Geom;
    	    	                L  : Location from TopLoc)
    returns Boolean
    is redefined;
    

    PCurve(me) returns any Curve from Geom2d
	---C++: return const &
    is redefined;
    
    PCurve(me : mutable; C : Curve from Geom2d)
    is redefined;
    
fields

    myPCurve : Curve from Geom2d;

end PointOnCurveOnSurface;
