-- Created on: 1993-02-05
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Contour from Contap

uses PathPoint               from IntSurf,
     PathPointTool           from IntSurf,
     SequenceOfPathPoint     from IntSurf,
     InteriorPoint           from IntSurf,
     InteriorPointTool       from IntSurf,
     SequenceOfInteriorPoint from IntSurf,
     Pnt                     from gp,
     Vec                     from gp,
     Point                   from Contap,
     Line                    from Contap,
     SurfFunction            from Contap,
     ArcFunction             from Contap,
     TheSequenceOfLine       from Contap,
     TheSearch               from Contap,
     TheSearchInside         from Contap,
     HSurface                from Adaptor3d,
     TopolTool               from Adaptor3d


raises NotDone           from StdFail,
       OutOfRange        from Standard,
       ConstructionError from Standard


is

    Create
    
    	returns Contour from Contap;


    Create(Direction: Vec from gp)
    
    	returns Contour from Contap;


    Create(Direction: Vec from gp; Angle: Real from Standard)
    
    	returns Contour from Contap;


    Create(Eye: Pnt from gp)
    
    	returns Contour from Contap;


    Create(Surf: HSurface from Adaptor3d; Domain: TopolTool from Adaptor3d; 
           Direction: Vec from gp)

	---Purpose: Creates the contour in a given direction.

    	returns Contour from Contap;


    Create(Surf: HSurface from Adaptor3d; Domain: TopolTool from Adaptor3d; 
           Direction: Vec from gp; Angle: Real from Standard)

	---Purpose: Creates the contour in a given direction.

    	returns Contour from Contap;


    Create(Surf: HSurface from Adaptor3d; Domain: TopolTool from Adaptor3d; 
           Eye: Pnt from gp)

	---Purpose: Creates the contour for a perspective view.

    	returns Contour from Contap;


    Perform(me: in out; Surf: HSurface from Adaptor3d; Domain: TopolTool from Adaptor3d)

	---Purpose: Creates the contour in a given direction.

    	raises ConstructionError from Standard
    	is static;


    Perform(me: in out; Surf: HSurface from Adaptor3d; Domain: TopolTool from Adaptor3d; 
                        Direction: Vec from gp)

	---Purpose: Creates the contour in a given direction.

    	is static;


    Perform(me: in out; Surf: HSurface from Adaptor3d; Domain: TopolTool from Adaptor3d; 
                        Direction: Vec from gp; Angle: Real from Standard)

	---Purpose: Creates the contour in a given direction.

    	is static;


    Perform(me: in out; Surf: HSurface from Adaptor3d; Domain: TopolTool from Adaptor3d; 
                        Eye: Pnt from gp)

	---Purpose: Creates the contour for a perspective view.

    	is static;


    Init(me: in out; Direction: Vec from gp)
    
    	is static;


    Init(me: in out; Direction: Vec from gp; Angle: Real from Standard)
    
    	is static;


    Init(me: in out; Eye: Pnt from gp)
    
    	is static;


    IsDone(me)
    
    	returns Boolean from Standard
	---C++: inline
	
	is static;


    IsEmpty(me)
    
    	---Purpose: Returns true if the is no line.

    	returns Boolean from Standard
	---C++: inline

    	raises NotDone from StdFail

    	is static;


    NbLines(me)
    
    	returns Integer from Standard
	---C++: inline
	
	raises NotDone from StdFail
	
	is static;
	
	
    Line(me; Index: Integer from Standard)
    
    	returns Line from Contap
	---C++: return const& 
	---C++: inline

	raises NotDone    from StdFail,
	       OutOfRange from Standard
	
	is static;


    SurfaceFunction(me : in out)
    returns SurfFunction
	---Purpose: Returns    a     reference   on     the   internal
	--          SurfaceFunction.  This is used to compute tangents
	--          on the lines.
        ---C++: return &
	---C++: inline
    is static;


    Perform(me: in out; Domain: TopolTool from Adaptor3d)
			   
	is static private;


    PerformAna(me: in out; Domain: TopolTool from Adaptor3d)
			   
	is static private;


fields

    done     : Boolean           from Standard;
    slin     : TheSequenceOfLine from Contap;
    solrst   : TheSearch         from Contap;
    solins   : TheSearchInside   from Contap;
    mySFunc  : SurfFunction      from Contap;
    myAFunc  : ArcFunction       from Contap;
    modeset  : Boolean           from Standard;

end Contour;
