-- Created on: 1997-09-18
-- Created by: Philippe MANGIN
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class LinearTension from FEmTool inherits ElementaryCriterion from FEmTool

	---Purpose: Criterium of LinearTension To Hermit-Jacobi  elements      

uses
   Vector  from  math, 
   Matrix  from  math,  
   Shape   from GeomAbs,
   HArray2OfReal  from  TColStd, 
   HArray2OfInteger  from TColStd   
    
raises 
  NotImplemented,   
  DomainError   
    
is
    Create(WorkDegree      : Integer ; 
           ConstraintOrder : Shape from GeomAbs)   
    returns LinearTension from FEmTool;        
     
    DependenceTable(me)  
    returns  HArray2OfInteger  from TColStd   
    is  redefined;  
    
    Value  (me  : mutable)  
    returns  Real  is  redefined; 
     
    Hessian(me  :  mutable ;  
	    Dimension1  :  Integer; 
	    Dimension2  :  Integer;
            H  :  out  Matrix  from  math)
     raises  DomainError -- If DependenceTable(Dimension1,Dimension2) is False 
     is  redefined;  
   
    Gradient(me  : mutable;   
	     Dimension  :  Integer;
             G  :  out  Vector  from  math) 
    is redefined;

fields 
RefMatrix  :  Matrix  from  math;  
myOrder    :  Integer; 
end LinearTension;
