-- Created on: 1996-02-15
-- Created by: PLOTNIKOV Eugeny
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class WNTGraphicDevice from Graphic3d inherits GraphicDevice from WNT

      	---Purpose: This class initializes a Windows NT Graphic Device.
        
uses

	Color		from Quantity,
	ColorRef	from WNT,
	Long		from WNT,
	SharedLibrary	from OSD,
	GraphicDriver	from Aspect,
	GraphicDriver	from Graphic3d

raises
 
	GraphicDeviceDefinitionError	from Aspect
  
is
 
	Create
		returns mutable WNTGraphicDevice from Graphic3d
	---Purpose: Creates a class instance and provide initialization
	--	    of the graphic library.
	--  Warning: Raises if something wrong.
	raises GraphicDeviceDefinitionError from Aspect;
 
	Create ( graphicLib : CString from Standard )
		returns mutable WNTGraphicDevice from Graphic3d
	---Purpose: Creates a class instance and provide initialization
	--	    of the graphic library defined by "graphicLib".
	--  Warning: Raises if something wrong.
	raises GraphicDeviceDefinitionError from Aspect;
   
	Destroy ( me : mutable )
		is redefined static;
	---Purpose: Destroys all resources attached to the graphic device.
	---C++:     alias~

	GraphicDriver ( me )
		returns GraphicDriver from Aspect
		is redefined static;
	---Level: Public
	---Purpose: Returns the GraphicDriver.

	SetGraphicDriver ( me	: mutable )
		is private;
	---Level: Internal
	---Purpose: Sets the GraphicDriver.

	SetGraphicDriver ( me	: mutable;
					   graphicLib : CString from Standard )
		is private;
	---Level: Internal
	---Purpose: Sets the GraphicDriver defined by "graphicLib".

fields

	MyGraphicDriver	:	GraphicDriver from Graphic3d;
	MySharedLibrary	:	SharedLibrary from OSD;

end WNTGraphicDevice;
