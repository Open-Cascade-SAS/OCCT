-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class OrientedFace from StepShape 

inherits Face from StepShape 

uses

	Boolean from Standard, 
	HArray1OfFaceBound from StepShape, 
	FaceBound from StepShape, 
	HAsciiString from TCollection
is

	Create returns mutable OrientedFace;
	---Purpose: Returns a OrientedFace


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aBounds : mutable HArray1OfFaceBound from StepShape) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aFaceElement : mutable Face from StepShape;
	      aOrientation : Boolean from Standard) is virtual;

	-- Specific Methods for Field Data Access --

	SetFaceElement(me : mutable; aFaceElement : mutable Face);
	FaceElement (me) returns mutable Face;
	SetOrientation(me : mutable; aOrientation : Boolean);
	Orientation (me) returns Boolean;
	SetBounds(me : mutable; aBounds : mutable HArray1OfFaceBound) is redefined;
	Bounds (me) returns mutable HArray1OfFaceBound is redefined;
	BoundsValue (me; num : Integer) returns mutable FaceBound is redefined;
	NbBounds (me) returns Integer is redefined;

fields

	faceElement : Face from StepShape;
	orientation : Boolean from Standard;

 -- 
 -- NB : field <bounds> inherited from classe <face> is redeclared.
 --      it shall appears in a physical file as a *.
 --

end OrientedFace;
