-- Created on: 1993-07-30
-- Created by: Jean-Louis FRENKEL
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class DatumAspect from Prs3d inherits CompositeAspect from Prs3d
    	---Purpose: A framework to define the display of datums.
uses

    LineAspect from Prs3d,
    Length from Quantity    
is

    Create returns mutable DatumAspect from Prs3d;
    	---Purpose: An empty framework to define the display of datums.
      
    FirstAxisAspect(me) returns mutable LineAspect from Prs3d;
    	---Purpose: Returns the attributes for display of the first axis.    
    SecondAxisAspect(me) returns mutable LineAspect from Prs3d;
    	---Purpose: Returns the attributes for display of the second axis.    
    ThirdAxisAspect(me) returns mutable LineAspect from Prs3d;
    	---Purpose: Returns the attributes for display of the third axis.    
    SetDrawFirstAndSecondAxis(me:mutable ; draw: Boolean from Standard);
    	---Purpose: Sets the DrawFirstAndSecondAxis attributes to active.    
    
    DrawFirstAndSecondAxis(me) returns Boolean from Standard; 
    	---Purpose: Returns true if the first and second axes can be drawn. 
    
    SetDrawThirdAxis(me:mutable; draw: Boolean from Standard);
    	---Purpose: Sets the DrawThirdAxis attributes to active.
    
    DrawThirdAxis(me) returns Boolean from Standard;
    	---Purpose: Returns true if the third axis can be drawn.    
    SetAxisLength(me:mutable; L1,L2,L3: Real from Standard);
    	---Purpose: Sets the lengths L1, L2 and L3 of the three axes. 
        
    FirstAxisLength(me) returns Length from Quantity;
    	--- Purpose: Returns the length of the displayed first axis.   
    
    SecondAxisLength(me) returns Length from Quantity;
    	---Purpose: Returns the length of the displayed second axis.    
    
    ThirdAxisLength(me) returns Length from Quantity;
    	---Purpose: Returns the length of the displayed third axis.
    
fields

    myFirstAxisAspect: LineAspect from Prs3d;
    mySecondAxisAspect: LineAspect from Prs3d;
    myThirdAxisAspect: LineAspect from Prs3d;
    myDrawFirstAndSecondAxis: Boolean from Standard;
    myDrawThirdAxis: Boolean from Standard;
    myFirstAxisLength: Length from Quantity;    
    mySecondAxisLength: Length from Quantity;    
    myThirdAxisLength: Length from Quantity;    
end DatumAspect from Prs3d;

