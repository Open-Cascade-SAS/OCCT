-- Created on: 1997-09-11
-- Created by: Philippe MANGIN
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



deferred class ElementaryCriterion from FEmTool inherits  TShared  from  MMgt

	---Purpose:  defined J Criteria to used in minimisation 

uses
   Vector  from  math, 
   Matrix  from  math,  
   HArray2OfReal  from  TColStd, 
   HArray2OfInteger  from TColStd 
    
raises 
  NotImplemented,   
  DomainError

is
    Set(me  :  mutable;   
        Coeff : HArray2OfReal) 
	 ---Purpose: Set the coefficient of the Element (the  Curve)
    is  static;
     
    Set(me : mutable; 
        FirstKnot  :  Real; 
        LastKnot   :  Real) 
	---Purpose: Set the definition interval of the Element         
    is virtual;  
     
    DependenceTable(me)  
    returns  HArray2OfInteger  from TColStd 
	---Purpose: To know if two dimension are independent.        
    is  deferred;  
    
    Value  (me  : mutable) 
    	---Purpose: To Compute J(E) where E  is the current Element        
    returns  Real  is  deferred;
     
    Hessian(me  :  mutable ;
	    Dim1  :  Integer; 
	    Dim2  :  Integer;
            H  :  out  Matrix  from  math) 
    ---Purpose: To Compute J(E)  the coefficients of Hessian matrix of
    --          J(E) wich are crossed derivatives in dimensions <Dim1>
    --          and  <Dim2>.          
     raises  DomainError -- If DependenceTable(Dimension1,Dimension2) is False 
     is  deferred;  
   
    Gradient(me   : mutable; 
	     Dim  :  Integer;
             G    :  out  Vector  from  math)     	 
    ---Purpose: To Compute the  coefficients in the dimension <dim> 
    --          of  the  J(E)'s  Gradient where E  is  the current  Element
    is  deferred;

fields 
  myCoeff           :  HArray2OfReal  is  protected; 
  myFirst,  myLast  :  Real is  protected;
end ElementaryCriterion;



