-- Created on: 1994-03-30
-- Created by: Laurent BUCHARD
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




generic class Classifier3d from TopClass 
    	(TheIntersector as any)  -- as Intersection3d from TopClass

	---Purpose: 

uses
    Lin             from gp,
    CurveTransition from TopTrans,
    Orientation     from TopAbs,
    State           from TopAbs,
    Face            from TopoDS

raises
    DomainError from Standard
    
is
    Create returns Classifier3d from TopClass;
	---Purpose: Creates an undefined classifier.
	
    Reset(me : in out; L   : Lin  from gp;
                       P   : Real from Standard; 
                       Tol : Real from Standard)
	---Purpose: Starts  a  classification process.   The  point to
	--          classify is the origin of  the  line <L>.  <P>  is
	--          the original length of the segment on <L>  used to
	--          compute  intersections.   <Tol> is the   tolerance
	--          attached to the intersections.
    is static;
    
    Compare(me : in out; F   : Face        from TopoDS;
                         Or  : Orientation from TopAbs)
	---Purpose: Updates  the classification process with  the face
	--          <F> from the boundary. 
    raises
    	DomainError  -- The classifier has not been set
    is static;

    Parameter(me) returns Real
	---Purpose: Returns the current value of the parameter.
	---C++: inline
    is static;

    HasIntersection(me) returns Boolean from Standard
    	---Purpose: Returns True if an intersection is computed.
    is static;

    Intersector(me : in out) returns TheIntersector
	---Purpose: Returns the intersecting algorithm.
	--          
	---C++: inline
	---C++: return &
    is static;
    
    State(me) returns State from TopAbs
	---Purpose: Returns the current state of the point.
	--          
	---C++: inline
    is static;
    

fields
    isSet          : Boolean          from Standard;
    myFace         : Face             from TopoDS;
    myLin          : Lin              from gp;
    myParam        : Real             from Standard;
    myTolerance    : Real             from Standard;
    myState        : State            from TopAbs;
    hasIntersect   : Boolean          from Standard;
    myIntersector  : TheIntersector;
    
end Classifier3d;

