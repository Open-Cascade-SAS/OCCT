-- Created on: 1995-10-23
-- Created by: Mister rmi
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Polygon3D from PBRep inherits CurveRepresentation from PBRep

	---Purpose: 

uses
    Polygon3D           from PPoly,
    CurveRepresentation from PBRep,
    Location            from PTopLoc

is

    Create(P: Polygon3D from PPoly;
    	   L: Location  from PTopLoc) 
    	---Purpose:
    returns mutable Polygon3D from PBRep;
        
    IsPolygon3D(me) returns Boolean
    	---Purpose: Returns True.
    is redefined;
    
    Polygon3D(me) returns any Polygon3D from PPoly;

fields

    myPolygon3D: Polygon3D from PPoly;

end Polygon3D;
