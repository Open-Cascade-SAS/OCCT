-- Created on: 1997-12-24
-- Created by: Xuan PHAM PHU
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Edge3dInterferenceTool from TopOpeBRepDS

---Purpose: a tool computing edge / face complex transition,
--          Interferences of edge reference are given by
--          I = (T on face, G = point or vertex, S = edge)

uses
    Pnt2d from gp,
    Pnt from gp,
    Dir from gp,
    Shape from TopoDS, 
    SurfaceTransition from TopTrans,
    Interference from TopOpeBRepDS
is
	  
    Create returns Edge3dInterferenceTool from TopOpeBRepDS;

    InitPointVertex(me : in out; 
            	    IsVertex : Integer;
    	    	    VonOO    : Shape from TopoDS);
	
    Init(me : in out; 
         Eref : Shape from TopoDS; 
	 E : Shape from TopoDS;   
	 F : Shape from TopoDS;
         I : Interference from TopOpeBRepDS);
    
    Add(me : in out; 
        Eref : Shape from TopoDS; 
	E : Shape from TopoDS;   
	F : Shape from TopoDS;
        I : Interference from TopOpeBRepDS);

    Transition(me; I : mutable Interference from TopOpeBRepDS)
    is static;

fields
    
    myFaceOriented : Integer;
    myTool         : SurfaceTransition from TopTrans;
    myTole         : Real; 
    myrefdef       : Boolean;

    myIsVertex     : Integer; -- 0 : geometry is a point
                              -- 1 : geometry is a vertex of reference
                              -- 2 : geometry is a vertex of the other shape
                              -- 3 : geometry is a vertex on the 2 shapes
    myVonOO        : Shape; -- only if myisvertex = 2,3
    myP3d          : Pnt from gp;
    myTgtref       : Dir from gp;

end Edge3dInterferenceTool from TopOpeBRepDS;
