-- Created on: 1995-07-17
-- Created by: Modelistation
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class BCurveTool from HLRBRep

uses 
     Array1OfReal from TColStd,
     Array1OfPnt  from TColgp,     
     Shape        from GeomAbs,
     CurveType    from GeomAbs,
     Vec          from gp,
     Pnt          from gp,
     Circ         from gp,
     Elips        from gp,
     Hypr         from gp,
     Parab        from gp,
     Lin          from gp,
     BezierCurve  from Geom,
     BSplineCurve from Geom,
     Curve        from BRepAdaptor
     
raises
    OutOfRange   from Standard,
    NoSuchObject from Standard,
    DomainError  from Standard
 
is
    --
    --     Global methods - Apply to the whole curve.
    --     
    
    FirstParameter(myclass; C: Curve from BRepAdaptor)
    returns Real from Standard;
    	---C++: inline
    

    LastParameter(myclass; C: Curve from BRepAdaptor)
    returns Real from Standard;
   	---C++: inline    

    --
    -- Services to break the curves to the expected continuity
    -- 
    --  If  for example you  need the  curve to  be C2  and the method
    --  Continuity   returns you something lower than   C2 (say C1 for
    --  example).
    --  
    --  First  compute the   number  of intervals  with  the requested
    --  continuity with the method  NbIntervals().   Note that if  the
    --  continuity  is higher than the one   you need NbIntervals will
    --  return 1.
    --  
    --  Then you get the parameters  bounding  the intervals with  the
    --  method  Intervals,   using   an array    of  length  at  least
    --  NbIntervals()+1.
    -- 
    -- If you need  to create a curve  with a restricted span you  can
    -- use the method Trim().

    
    Continuity(myclass; C: Curve from BRepAdaptor)
    returns Shape from GeomAbs;
	---Purpose: 
	---C++: inline
    
    NbIntervals(myclass; C : in out Curve from BRepAdaptor;
                         S : Shape from GeomAbs)
    returns Integer from Standard;
	---Purpose: Returns  the number  of  intervals for  continuity
	--          <S>. May be one if Continuity(myclass) >= <S>
	---C++: inline
    
    Intervals(myclass; C : in out Curve        from BRepAdaptor;
                       T : in out Array1OfReal from TColStd; 
    	               S :        Shape        from GeomAbs)
	---Purpose: Stores in <T> the  parameters bounding the intervals
	--          of continuity <S>.
	--          
	--          The array must provide  enough room to  accomodate
	--          for the parameters. i.e. T.Length() > NbIntervals()
    raises OutOfRange from Standard;
    	---C++: inline
    
    IsClosed(myclass; C: Curve from BRepAdaptor)
    returns Boolean from Standard;
    	---C++: inline    
     
    IsPeriodic(myclass; C: Curve from BRepAdaptor)
    returns Boolean from Standard;
    	---C++: inline
    
    Period(myclass; C: Curve from BRepAdaptor)
    returns Real from Standard
    raises DomainError from Standard;
    	---C++: inline	
     
    Value(myclass; C : Curve from BRepAdaptor;
                   U : Real  from Standard)
    returns Pnt from gp;
    	--- Purpose : Computes the point of parameter U on the curve.
    	---C++: inline
    
    D0 (myclass; C :     Curve from BRepAdaptor;
                 U :     Real  from Standard;
                 P : out Pnt   from gp);
        --- Purpose : Computes the point of parameter U on the curve.
    	---C++: inline
    
    D1 (myclass; C :     Curve from BRepAdaptor;
                 U :     Real  from Standard;
                 P : out Pnt   from gp ;
                 V : out Vec   from gp)
        --- Purpose : Computes the point of parameter U on the curve with its
        --  first derivative.
     raises DomainError from Standard;
        --- Purpose : Raised if the continuity of the current interval
        --  is not C1.
    	---C++: inline
    
    D2 (myclass; C      :     Curve from BRepAdaptor;
                 U      :     Real  from Standard;
                 P      : out Pnt   from gp;
                 V1, V2 : out Vec   from gp)
        --- Purpose :
        --  Returns the point P of parameter U, the first and second
        --  derivatives V1 and V2.
     raises DomainError from Standard;
        --- Purpose : Raised if the continuity of the current interval
        --  is not C2.
    	---C++: inline

    D3 (myclass; C          :     Curve from BRepAdaptor;
                 U          :     Real  from Standard;
                 P          : out Pnt   from gp;
                 V1, V2, V3 : out Vec   from gp)
        --- Purpose :
        --  Returns the point P of parameter U, the first, the second 
        --  and the third derivative.
     raises DomainError from Standard;
        --- Purpose : Raised if the continuity of the current interval
        --  is not C3.
    	---C++: inline
        
    DN (myclass; C : Curve   from BRepAdaptor;
                 U : Real    from Standard;
                 N : Integer from Standard)
    returns Vec from gp
        --- Purpose :
        --  The returned vector gives the value of the derivative for the 
        --  order of derivation N.
    raises  
    	DomainError from Standard,
        --- Purpose : Raised if the continuity of the current interval
        --  is not CN.
        OutOfRange from Standard;
        --- Purpose : Raised if N < 1.            
	---C++: inline

    Resolution(myclass; C   : Curve from BRepAdaptor;
                        R3d : Real  from Standard)
    returns Real from Standard;
        ---Purpose :  Returns the parametric  resolution corresponding
        --         to the real space resolution <R3d>.
	---C++: inline
        
    GetType(myclass; C: Curve from BRepAdaptor)
    returns CurveType from GeomAbs;
    	---Purpose: Returns  the  type of the   curve  in the  current
	--          interval :   Line,   Circle,   Ellipse, Hyperbola,
	--          Parabola, BezierCurve, BSplineCurve, OtherCurve.
	---C++: inline

    --
    --     The following methods must  be called when GetType returned
    --     the corresponding type.
    --     

    Line(myclass; C: Curve from BRepAdaptor)
    returns Lin from gp
    raises NoSuchObject from Standard;
	---C++: inline
     
    Circle(myclass; C: Curve from BRepAdaptor)
    returns Circ from gp
    raises NoSuchObject from Standard;
    	---C++: inline
     
    Ellipse(myclass; C: Curve from BRepAdaptor)
    returns Elips from gp
    raises NoSuchObject from Standard;
    	---C++: inline
     
    Hyperbola(myclass; C: Curve from BRepAdaptor)
    returns Hypr from gp
    raises NoSuchObject from Standard;
    	---C++: inline
     
    Parabola(myclass; C: Curve from BRepAdaptor)
    returns Parab from gp
    raises NoSuchObject from Standard;
    	---C++: inline
     
    Bezier(myclass; C: Curve from BRepAdaptor)
    returns BezierCurve from Geom
    raises NoSuchObject from Standard;
    
    BSpline(myclass; C: Curve from BRepAdaptor)
    returns BSplineCurve from Geom
    raises NoSuchObject from Standard;

    Degree(myclass; C: Curve from BRepAdaptor)
    returns Integer from Standard;
    	---C++: inline
    
    IsRational(myclass; C: Curve from BRepAdaptor)
    returns Boolean from Standard;
    	---C++: inline
    
    NbPoles(myclass; C: Curve from BRepAdaptor)
    returns Integer from Standard;
	---C++: inline

    NbKnots(myclass; C: Curve from BRepAdaptor)
    returns Integer from Standard;
    	---C++: inline

    Poles(myclass; C :        Curve       from BRepAdaptor;
                   T : in out Array1OfPnt from TColgp);

    PolesAndWeights(myclass; C :        Curve        from BRepAdaptor;
                             T : in out Array1OfPnt  from TColgp; 
                             W : in out Array1OfReal from TColStd);

    NbSamples(myclass; C     : Curve from BRepAdaptor;
                       U0,U1 : Real  from Standard) 
    returns Integer from Standard;

end BCurveTool;
