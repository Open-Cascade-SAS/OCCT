-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class PresentationStyleSelect from StepVisual inherits SelectType from StepData

	-- <PresentationStyleSelect> is an EXPRESS Select Type construct translation.
	-- it gathers : PointStyle, CurveStyle, SurfaceStyleUsage, SymbolStyle, FillAreaStyle, TextStyle
	-- Rev4 : only remain PointStyle, CurveStyle, SurfaceStyleUsage

uses

	PointStyle,
	CurveStyle,
	SurfaceStyleUsage
--	SymbolStyle,
--	FillAreaStyle,
--	TextStyle
is

	Create returns PresentationStyleSelect;
	---Purpose : Returns a PresentationStyleSelect SelectType

	CaseNum (me; ent : Transient) returns Integer;
	---Purpose: Recognizes a PresentationStyleSelect Kind Entity that is :
	--        1 -> PointStyle
	--        2 -> CurveStyle
	--        3 -> SurfaceStyleUsage
	--        4 -> SymbolStyle
	--        5 -> FillAreaStyle
	--        6 -> TextStyle
	--        0 else

	PointStyle (me) returns any PointStyle;
	---Purpose : returns Value as a PointStyle (Null if another type)

	CurveStyle (me) returns any CurveStyle;
	---Purpose : returns Value as a CurveStyle (Null if another type)

	SurfaceStyleUsage (me) returns any SurfaceStyleUsage;
	---Purpose : returns Value as a SurfaceStyleUsage (Null if another type)

end PresentationStyleSelect;

