-- Created on: 1996-09-04
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class DPrism from LocOpe 

	---Purpose: Defines a  pipe  (near from   Pipe from BRepFill),
	--          with modifications provided for the Pipe feature.

uses Evolved from BRepFill,
     DataMapOfShapeListOfShape    from TopTools,
     ListOfShape  from TopTools,
     
     Shape from TopoDS,
     Wire  from TopoDS,
     Edge  from TopoDS, 
     Face  from TopoDS,
     Curve from Geom,
     SequenceOfPnt   from TColgp,
     SequenceOfCurve from TColGeom
     

raises NoSuchObject from Standard,
       DomainError  from Standard,
       NotDone      from StdFail

is

    Create (Spine     : Face from TopoDS;
            Height1   : Real from Standard;
	    Height2   : Real from Standard;
	    Angle     : Real from Standard)
	    
	returns DPrism from LocOpe;     

    Create (Spine     : Face from TopoDS;
    	    Height    : Real from Standard;
	    Angle     : Real from Standard)

    	returns DPrism from LocOpe;


    IsDone(me)
    
    	returns Boolean from Standard
	is static;


    Spine(me)
    
    	returns Shape from TopoDS
	---C++: return const &
	is static;


    Profile(me)
    
    	returns Shape from TopoDS
	---C++: return const &
	is static;


    FirstShape(me)
    
    	returns Shape from TopoDS
	---C++: return const &
	is static;


    LastShape(me)
    
    	returns Shape from TopoDS
	---C++: return const &
	is static;


    Shape(me)
    
    	returns Shape from TopoDS
	---C++: return const &
    	raises NotDone from StdFail
	is static;


    Shapes(me; S: Shape from TopoDS)
    
    	returns ListOfShape from TopTools
	---C++: return const &
    	raises NoSuchObject from Standard,
	       -- The exception is raised if S is not a subshape of the profile
               DomainError  from Standard,
	       -- The exception is raised if S is neither a vertex nor
	       -- an edge
    	       NotDone from StdFail
	is static;


    Curves(me;  SCurves:  in  out  SequenceOfCurve  from  TColGeom)
    
	is static;
 
    BarycCurve(me) 
     
    	returns  Curve  from  Geom 
	is  static;

    IntPerf(me:  in  out) 
     
    	is  static  private;
  
fields

    myDPrism     : Evolved         from BRepFill;
    myRes        : Shape           from TopoDS;
    mySpine      : Face            from TopoDS; 
    myProfile    : Wire            from TopoDS;
    myProfile1   : Edge            from TopoDS;
    myProfile2   : Edge            from TopoDS;
    myProfile3   : Edge            from TopoDS;
    myHeight     : Real            from Standard;
    myFirstShape : Shape           from TopoDS;
    myLastShape  : Shape           from TopoDS;
    myCurvs      : SequenceOfCurve from TColGeom;
    myMap        : DataMapOfShapeListOfShape    from TopTools;
    
end DPrism;     
