-- Created on: 1993-06-21
-- Created by: Martine LANGLOIS
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class MakeBoundedCurve from GeomToStep inherits Root from GeomToStep

    ---Purpose: This class implements the mapping between classes 
    --          BoundedCurve from Geom, Geom2d and the class BoundedCurve from 
    --          StepGeom which describes a BoundedCurve from prostep.
    --          As BoundedCurve is an abstract BoundedCurve this class 
    --          is an access to the sub-class required.
  
uses BoundedCurve from Geom,
     BoundedCurve from Geom2d,
     BoundedCurve from StepGeom
     
raises NotDone from StdFail
     
is 

Create ( C : BoundedCurve from Geom ) returns MakeBoundedCurve;

Create ( C : BoundedCurve from Geom2d ) returns MakeBoundedCurve;

Value (me) returns BoundedCurve from StepGeom
    raises NotDone
    is static;
    ---C++: return const&
 
fields

    theBoundedCurve : BoundedCurve from StepGeom;
    	-- The solution from StepGeom
    	
end MakeBoundedCurve;



