-- Created on: 1992-08-18
-- Created by: Modelistation
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

private class Line from Hatch

	---Purpose: Stores a Line in the Hatcher. Represented by :
	--          
	--          * A Lin2d from gp, the geometry of the line.
	--          
	--          * Bounding parameters for the line.
	--          
	--          * A sorted List  of Parameters, the  intersections
	--          on the line.

uses
    Real                from Standard,
    Integer             from Standard,
    Boolean             from Standard,
    Lin2d               from gp,
    LineForm            from Hatch,
    SequenceOfParameter from Hatch

is

    Create;
    
    Create(L : Lin2d from gp; T : LineForm from Hatch)
    returns Line from Hatch;
    
    AddIntersection(me       : in out; 
                    Par1     : Real    from Standard;
		    Start    : Boolean from Standard;
                    Index    : Integer from Standard;
                    Par2     : Real    from Standard;
    	    	    theToler : Real    from Standard)
	---Purpose: Insert a new intersection in the sorted list.
    is static;
    
fields

    myLin    : Lin2d               from gp;
    myForm   : LineForm            from Hatch;
    myInters : SequenceOfParameter from Hatch;

friends
    class Hatcher from Hatch

end Line;
