-- Created on: 1993-03-23
-- Created by: BBL
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Modified:	02-06-98 : FMN ; Suppression appel Clear (deja fait dans ALienData)

class SunRFAlienImage from AlienImage inherits AlienUserImage from AlienImage

	
	---Purpose: Defines a SunRF Alien image, i.e. an image using the
-- image format for SUN workstations.

uses
	File 			from OSD,
	AsciiString 		from TCollection,
	ColorImage 		from Image,
	PseudoColorImage 	from Image,
	Image			from Image,
	SunRFAlienData 		from AlienImage,
	SUNRFFormat	 	from AlienImage

is
	Create returns mutable SunRFAlienImage from AlienImage;
---Purpose: Constructs an empty SunRF alien image.
    
	Clear( me : in out mutable) ;
	---Level: Public
	---Purpose: Frees memory allocated by SunRFAlienImage

	ToImage( me : in immutable ) 
	  returns mutable Image from Image ;
	---Level: Public
	  ---Purpose : Converts a SunRFAlienImage object to a Image object.

	FromImage( me : in out mutable ; anImage : in Image from Image ) ;
	---Level: Public
	  ---Purpose : Converts an Image object to a SunRFAlienImage object.

	Read ( me : in out mutable; afile : in out File from OSD )
	  returns Boolean from Standard ;
	---Level: Public
	  ---Purpose: Reads the content of a  SunRFAlienImage object from a file
	  --          Returns True if file is a XWD file .

	Write( me : in immutable; afile : in out File from OSD )
	  returns Boolean from Standard ;
	  ---Purpose: Writes content of a  SunRFAlienImage object to a file

	SetFormat( me : in out mutable ;
		   aFormat : SUNRFFormat from AlienImage);
	  ---Purpose: Sets the  SUN Raster File Format for Write method.

	Format( me : in  immutable )
	    returns SUNRFFormat from AlienImage ;
	  ---Purpose: Returns the SUN Raster File Format .

fields
	myData : SunRFAlienData from AlienImage ;

end ;
 
