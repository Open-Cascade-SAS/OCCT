-- Created on: 1993-01-11
-- Created by: CKY / Contract Toubro-Larsen ( Anand NATRAJAN )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class FlowLineSpec from IGESAppli  inherits IGESEntity

        ---Purpose: defines FlowLineSpec, Type <406> Form <14>
        --          in package IGESAppli
        --          Attaches one or more text strings to entities being
        --          used to represent a flow line

uses

        HAsciiString          from TCollection,
        HArray1OfHAsciiString from Interface

raises OutOfRange

is

        Create returns mutable FlowLineSpec;

        -- Specific Methods pertaining to the class

        Init (me : mutable; allProperties : HArray1OfHAsciiString);
        ---Purpose : This method is used to set the fields of the class
        --           FlowLineSpec
        --       - allProperties : primary flow line specification and modifiers

        NbPropertyValues (me) returns Integer;
        ---Purpose : returns the number of property values

        FlowLineName (me) returns HAsciiString from TCollection;
        ---Purpose : returns primary flow line specification name

        Modifier (me; Index : Integer) returns HAsciiString from TCollection
        raises OutOfRange;
        ---Purpose : returns specified modifier element
        -- raises exception if Index <= 1 or Index > NbPropertyValues

fields

--
-- Class    : IGESAppli_FlowLineSpec
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class FlowLineSpec.
--
-- Reminder : A FlowLineSpec instance is defined by :
--            - primary flow line specification name and modifiers

        theNameAndModifiers : HArray1OfHAsciiString;

end FlowLineSpec;
