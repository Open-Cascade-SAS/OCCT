-- Created on: 1997-08-07
-- Created by: Jean-Louis Frenkel
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Directory from CDF inherits Transient from Standard


---Purpose: A directory is a collection of documents. There is only one instance
--          of a given document in a directory.
--          put.

uses Document from CDM, ListOfDocument from CDM

raises  NoSuchObject
    
is
    Create 
    returns Directory from CDF;
    ---Purpose: Creates an empty directory.
    
    
    Add(me:mutable; aDocument: Document from CDM);
    ---Purpose: adds a document into the directory.
    
    Remove(me: mutable; aDocument: Document from CDM);
    ---Purpose: removes the document.
    
    
---Category: Inquire Methods
--           

    Contains(me; aDocument: Document from CDM) 
    ---Purpose: Returns true if the document aDocument is in the directory
    returns Boolean from Standard
    is static;

    Last(me:mutable) returns Document from CDM
    ---Purpose: returns the last document (if any) which has been added
    --          in the directory.
    raises NoSuchObject from Standard
    ---Warning: if the directory is empty.
    is static;

    Length(me) returns Integer from Standard
    ---Purpose: returns the number of documents of the directory.
    is static;

    IsEmpty(me) returns Boolean from Standard
    ---Purpose: returns true if the directory is empty.
    is static;
    
---Category: Private methods
   
   List(me) returns ListOfDocument from CDM
   is static private;
   ---C++: return const &
   --      
   
fields

    myDocuments: ListOfDocument from CDM;

friends    
    class DirectoryIterator from CDF

end Directory from CDF;
