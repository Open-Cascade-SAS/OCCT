-- Created on: 1996-04-03
-- Created by: Stagiaire Frederic CALOONE
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Modified:	Wed Mar  5 09:45:42 1997
--    by:	Joelle CHAUVET
--              G1134 : New methods EcartContraintes, EcartContour,
--                      Disc2dContour, Disc3dContour,
--                      Surface, Sense, Curves2d,
--                      for using of GeomPlate_MakeApprox
--              + no more reference to TopoDS (suppression of method Face)
-- Modified:
--              New fields myTolCurv, myAnisotropie
--              and new method ComputeAnisotropie
--              New methods G0Eror( Index ), G1Error( Index ), G2Error( Index )

class BuildPlateSurface from GeomPlate
    	---Purpose:
    	-- This class provides an algorithm for constructing such a plate surface that
    	-- it conforms to given curve and/or point constraints.
    	-- The algorithm accepts or constructs an initial surface
    	-- and looks for a deformation of it satisfying the
    	-- constraints and minimizing energy input.
    	-- A BuildPlateSurface object provides a framework for:
    	-- -   defining or setting constraints
    	-- -   implementing the construction algorithm
    	-- -   consulting the result.


uses Pnt from gp,
     Plate from Plate,
     Surface from GeomPlate,
     Surface from Geom,
     HArray1OfInteger from TColStd,
     Array1OfInteger from TColStd,
     HArray1OfReal from TColStd,
     HArray2OfReal from TColStd,
     HArray1OfCurve from TColGeom2d,
     SequenceOfXY from TColgp,
     SequenceOfXYZ from TColgp,
     HArray1OfHCurveOnSurface from GeomPlate,
     Array1OfHCurveOnSurface from GeomPlate,
     CurveConstraint  from  GeomPlate, 
     PointConstraint  from  GeomPlate, 
     HSequenceOfCurveConstraint from GeomPlate, 
     HSequenceOfPointConstraint  from  GeomPlate, 
     HArray1OfPnt2d  from  TColgp, 
     HArray1OfSequenceOfReal from GeomPlate, 
     ExtPS  from Extrema, 
     Pnt2d  from  gp, 
     HCurve  from  Adaptor3d, 
     HCurve2d  from  Adaptor2d,
     Curve  from  Geom2d
      
raises   
     ConstructionError  from  Standard, 
     RangeError  from  Standard      
     
is
  Create(  NPoints : HArray1OfInteger from TColStd;
    	   TabCurve : HArray1OfHCurveOnSurface from GeomPlate;
	   Tang : HArray1OfInteger from TColStd;
    	   Degree : Integer from Standard;  
	   NbIter  :  Integer  from  Standard  =  3;
	   Tol2d  :  Real  from  Standard  =  0.00001;
	   Tol3d  :  Real  from  Standard  =  0.0001; 
	   TolAng  :  Real  from  Standard  =  0.01; 
	   TolCurv : Real  from  Standard  =  0.1;
	   Anisotropie : Boolean from Standard = Standard_False )
           returns BuildPlateSurface from  GeomPlate 
	   raises  ConstructionError;
	   
    	--- Purpose : Constructor  compatible  with  the  old  version
    	-- with this constructor the constraint are given in a Array of Curve on Surface
    	-- The array NbPoints  contains the number of points for each constraint.
    	-- The Array Tang contains the order of constraint for each Constraint: The possible values for this
    	-- order has to be -1 , 0 , 1 , 2 . Order i means constraint Gi.
    	-- NbIter is the maximum number of iteration to optimise the number of points for resolution
    	-- Degree is the degree of resolution for Plate
    	-- Tol2d is the tolerance used to test if two points of different constraint are identical in the 
    	-- parametric space of the initial surface
    	-- Tol3d is used to test if two identical points in the 2d space are identical in 3d space
    	-- TolAng is used to compare the angle between normal of two identical points in the 2d space
    	-- Raises  ConstructionError;
       	--if NbIter<1 or length of TabCurve is <1 or Degree <  2 
    
    Create  ( Surf  :  Surface  from  Geom;   
    	      Degree  :  Integer  from  Standard  =  3;   
    	      NbPtsOnCur  :  Integer  from  Standard  =  10 ; 
	      NbIter  :  Integer  from  Standard  =  3;
	      Tol2d  :  Real  from  Standard  =  0.00001;
	      Tol3d  :  Real  from  Standard  =  0.0001; 
	   TolAng  :  Real  from  Standard  =  0.01;
	   TolCurv : Real  from  Standard  =  0.1;
           Anisotropie : Boolean from Standard = Standard_False )
            returns  BuildPlateSurface  from  GeomPlate
 	   raises  ConstructionError;
	   --if NbIter<1 or Degree <  2
    
    Create  (Degree  :  Integer  from  Standard =  3;   
             NbPtsOnCur  :  Integer  from  Standard  =  10; 
	     NbIter  :  Integer  from  Standard  =  3;
	     Tol2d  :  Real  from  Standard  =  0.00001;
	     Tol3d  :  Real  from  Standard  =  0.0001; 
	   TolAng  :  Real  from  Standard  =  0.01;
	   TolCurv : Real  from  Standard  =  0.1;
	   Anisotropie : Boolean from Standard = Standard_False )
            returns  BuildPlateSurface  from  GeomPlate 
 	   raises  ConstructionError;
    	---Purpose: Initializes the BuildPlateSurface framework for
    	-- deforming plate surfaces using curve and point
    	-- constraints. You use the first constructor if you have
    	-- an initial surface to work with at construction time. If
    	-- not, you use the second. You can add one later by
    	-- using the method LoadInitSurface. If no initial
    	-- surface is loaded, one will automatically be computed.
    	-- The curve and point constraints will be defined by
    	-- using the method Add.
    	-- Before the call to the algorithm, the curve constraints
    	-- will be transformed into sequences of discrete points.
    	-- Each curve defined as a constraint will be given the
    	-- value of NbPtsOnCur as the average number of points on it.
    	-- Several arguments serve to improve performance of
    	-- the algorithm. NbIter, for example, expresses the
    	-- number of iterations allowed and is used to control the
    	-- duration of computation. To optimize resolution,
    	-- Degree will have the default value of 3.
    	-- The surface generated must respect several tolerance values:
    	-- -   2d tolerance given by Tol2d, with a default value of 0.00001
    	-- -   3d tolerance expressed by Tol3d, with a default value of 0.0001
    	-- -   angular tolerance given by TolAng, with a default
    	--   value of 0.01, defining the greatest angle allowed
    	--   between the constraint and the target surface.
    	-- Exceptions
    	-- Standard_ConstructionError if NbIter is less than 1 or Degree is less than 3.
    
    Init  (me:  in  out);
    	--- Purpose:  Resets all constraints

    LoadInitSurface  (me  :  in  out;  Surf  :  Surface  from  Geom);
    	--- Purpose: Loads the initial Surface
    
    Add  (me  :  in  out;Cont  :  CurveConstraint  from  GeomPlate); 
    	---Purpose: Adds the linear constraint cont.  
    SetNbBounds (me : in out; NbBounds : Integer from Standard);
         
    Add  (me  :  in  out;Cont  :  PointConstraint  from  GeomPlate); 
    	---Purpose: Adds the point constraint cont. 
    Perform ( me: in out ) 
    raises RangeError; 
    	---Purpose:
    	-- Calls the algorithm and computes the plate surface using
    	-- the loaded constraints. If no initial surface is given, the
    	-- algorithm automatically computes one.
    	-- Exceptions
    	-- Standard_RangeError if the value of the constraint is
    	-- null or if plate is not done.
     
    CurveConstraint(me  ;  order  :  Integer  from  Standard)   
    returns  CurveConstraint  from  GeomPlate; 
    	--- Purpose : returns the CurveConstraints of order order
    	--  

    PointConstraint(me  ;  order  :  Integer  from  Standard)   
    returns  PointConstraint  from  GeomPlate ;
    	---Purpose : returns the PointConstraint of order order
    	--         
         

    Disc2dContour (me :in  out; nbp : Integer from Standard; 
                        Seq2d : out SequenceOfXY from TColgp);  
    --   for the moment, nbp can be equal to 1, 2 or 4 if nbp = 1, the
    --   evaluation takes place only on constraints points (*)
    --   
    --   --*-------*---------------*-------------------*---------------*--
    --   
    --   if nbp = 2, middle points (+) are added to constraints points
    --   
    --   --*---+---*-------+-------*---------+---------*-------+-------*--
    --   
    --   if nbp = 4, quarter points (o) and middle points (+) are added to constraints points
    --   
    --   --*-o-+-o-*---o---+---o---*----o----+----o----*---o---+---o---*--
    --   computes 2d constraints on Frontiere
    --   see EcartContraintes for nbp
    
    Disc3dContour (me :in  out; nbp : Integer from Standard;
                        iordre : Integer from Standard; 
                    	Seq3d : out SequenceOfXYZ from TColgp);  
    --   computes 3d G0 constraints on Frontiere if iordre = 0
    --   computes 3d G1 constraints on Frontiere if iordre = 1
-- see Disc2dContour for nbp
	    
    IsDone ( me ) returns Boolean;
    	--- Purpose:
    	-- Tests whether computation of the plate has been completed.
    Surface ( me ) returns Surface from GeomPlate;  
    	---Purpose:
    	-- Returns the result of the computation. This surface can
    	-- then be used by GeomPlate_MakeApprox for
    	-- converting the resulting surface into a BSpline.
     
    SurfInit  (me)  returns  Surface  from  Geom;
    	---Purpose: Returns the initial surface
	    
    Sense ( me ) returns HArray1OfInteger from TColStd;
    	---Purpose:
    	-- Allows you to ensure that the array of curves returned by
    	-- Curves2d has the correct orientation. Returns the
    	-- orientation of the curves in the the array returned by
    	-- Curves2d. Computation changes the orientation of
    	-- these curves. Consequently, this method returns the
    	-- orientation prior to computation.    
    Curves2d ( me ) returns HArray1OfCurve from TColGeom2d; 
    	--- Purpose:
    	-- Extracts the array of curves on the plate surface which
    	-- correspond to the curve constraints set in Add.    
    Order ( me ) returns HArray1OfInteger from TColStd; 
    	---Purpose:
    	-- Returns the order of the curves in the array returned by
    	-- Curves2d. Computation changes this order.
    	-- Consequently, this method returns the order of the
    	-- curves prior to computation.     
    G0Error  (me)  returns  Real  from  Standard; 
    	---Purpose: Returns the max distance betwen the result and the constraints

    G1Error  (me)  returns  Real  from  Standard; 
     	---Purpose: Returns  the max angle betwen the result and the constraints

    G2Error  (me)  returns  Real  from  Standard; 
    	---Purpose: Returns  the max difference of curvature betwen the result and the constraints
    -- 
    G0Error( me : in out; Index : Integer from Standard ) returns Real from Standard;
    	---Purpose: Returns   the max distance between the result and the constraint Index
    
    G1Error( me : in out; Index : Integer from Standard ) returns Real from Standard;
    	---Purpose: Returns the max angle between the result and the constraint Index
    
    G2Error( me : in out; Index : Integer from Standard ) returns Real from Standard;
     	---Purpose: Returns the max difference of curvature between the result and the constraint Index
    --
    EcartContraintesMil (me : in out; c : Integer from Standard; 
                    	    	   d,an,courb : out HArray1OfReal from TColStd )  is  private;  
    
    	--- Purpose: Evaluates the distance, the angle between normals, and the "courbure"
   	--   on middle points of contraints an corresponding points on the GeomPlate_Surface
    	--   the results are given for a curve c
   
    ----Private methods 

    ProjectPoint  (me :in  out  ;  P  :  Pnt  from  gp)   
                    returns  Pnt2d  from  gp  is  private; 
		    
    ProjectCurve  (me :in  out  ;  Curv  :  HCurve  from  Adaptor3d)   
                    returns  Curve  from  Geom2d  is  private;
 
    ProjectedCurve  (me :in  out  ;  Curv  :  in  out  HCurve  from  Adaptor3d)   
                    returns  HCurve2d  from  Adaptor2d  is  private;                                                                                 
									  
    ComputeSurfInit (me : in out)
    is  private;
     
    Intersect  (me  :  in  out;   
                PntInter  : out HArray1OfSequenceOfReal from  GeomPlate; 
                PntG1G1   : out HArray1OfSequenceOfReal from  GeomPlate )   
    is  private; 
    
    Discretise  (me  :  in  out; 
    	    	PntInter  : HArray1OfSequenceOfReal from  GeomPlate; 
                PntG1G1   : HArray1OfSequenceOfReal from  GeomPlate )   
    is  private; 
        
    LoadCurve  (me  :  in  out; NbBoucle : Integer from Standard;
                    	    	OrderMax : Integer = 2)
    is  private;  
     
    LoadPoint  (me  :  in  out; NbBoucle : Integer from Standard;
                    	    	OrderMax : Integer = 2)
    is  private;    

    CalculNbPtsInit  (me  :  in  out)  is  private;  
     
    VerifSurface (me  :  in  out  ;  NbLoop  :  Integer)    
    returns Boolean  from  Standard  
    is  private; 

    VerifPoints (me;  dist,ang,curv  :  out  Real  from  Standard)  is  private; 
   
    CourbeJointive (me : in out; tolerance : Real from Standard)  
    returns Boolean  from  Standard  is  private;

    ComputeAnisotropie(me) returns Real from Standard
    is private;
    
    IsOrderG1(me) returns Boolean from Standard
    is private;
    
fields
    myLinCont : HSequenceOfCurveConstraint from GeomPlate;  
    myParCont  :  HArray1OfSequenceOfReal from GeomPlate;
    myPlateCont  :  HArray1OfSequenceOfReal from GeomPlate;
    myPntCont  :  HSequenceOfPointConstraint  from  GeomPlate;
    mySurfInit : Surface from Geom; 
    myPlanarSurfInit : Surface from Geom;
    myGeomPlateSurface : Surface from GeomPlate;
    myPlate : Plate from Plate;
    myPrevPlate : Plate from Plate;
    myAnisotropie : Boolean from Standard;
    mySense : HArray1OfInteger from TColStd;
    myDegree : Integer from Standard;
    myInitOrder :  HArray1OfInteger from TColStd;  
    myG0Error  :  Real  from  Standard; 
    myG1Error  :  Real  from  Standard; 
    myG2Error  :  Real  from  Standard; 
    myNbPtsOnCur  :  Integer  from  Standard;  
    mySurfInitIsGive  :  Boolean  from  Standard;
    myNbIter  :  Integer  from  Standard; 
    myProj  :  ExtPS  from Extrema;
    --   TOLERANCE
     
    myTol2d  :   Real  from  Standard; 
    myTol3d  :   Real  from  Standard; 
    myTolAng  :   Real  from  Standard;  
    myTolU  :  Real  from  Standard;  
    myTolV  :  Real  from  Standard;
    
    myNbBounds : Integer from Standard;
     
    myIsLinear : Boolean from Standard;
    myFree     : Boolean from Standard;

end;
