-- Created on: 1998-07-16
-- Created by: CAL
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Updated:     GG IMP230300 The color fields are moved in Aspect_Grid

private class CircularGrid from V3d inherits CircularGrid from Aspect

uses
	Ax3			from gp,
	Color			from Quantity,
	Group			from Graphic3d,
	Structure		from Graphic3d,
	GridDrawMode		from Aspect,
	ViewerPointer		from V3d

is
	Create ( aViewer	: ViewerPointer from V3d;
		 aColor		: Color from Quantity;
		 aTenthColor	: Color from Quantity )
	returns CircularGrid from V3d;

	SetColors ( me	: mutable;
		    aColor	: Color from Quantity;
		    aTenthColor	: Color from Quantity )
	is redefined static;

	Display ( me	: mutable )
	is redefined static;
   
	Erase ( me )
	is redefined static;

	IsDisplayed ( me )
	returns Boolean from Standard
	is redefined static;

	GraphicValues ( me; 
			Radius	: out Real from Standard;
			OffSet	: out Real from Standard )
	is static;

	SetGraphicValues ( me	: mutable; 
			   Radius	: Real from Standard;
			   OffSet	: Real from Standard )
	is static;

	DefineLines ( me : mutable )
	is static private;

	DefinePoints ( me : mutable )
	is static private;

	UpdateDisplay ( me	: mutable )
	is redefined static protected;

fields
	myStructure		: Structure from Graphic3d;
	myGroup	        : Group from Graphic3d;
	myCurViewPlane	: Ax3 from gp;
	myViewer		: ViewerPointer from V3d;
	myCurAreDefined		: Boolean from Standard;
	myCurDrawMode		: GridDrawMode from Aspect;
	myCurXo, myCurYo	: Real from Standard;
	myCurAngle		: Real from Standard;
	myCurStep		: Real from Standard;
	myCurDivi		: Integer from Standard;
	myRadius		: Real from Standard;
	myOffSet		: Real from Standard;

end CircularGrid from V3d;
