-- Created on: 1993-10-14
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class Cut from BRepAlgoAPI inherits BooleanOperation from BRepAlgoAPI
	---Purpose:  The class Cut provides a Boolean
    	-- cut operation on a pair of arguments (Boolean Subtraction).
    	-- The class Cut provides a framework for:
    	--   -      Defining the construction of a cut shape
    	--   -      Implementing the building algorithm
    	--   -      Consulting the result

uses
    Shape from TopoDS,
    PaveFiller from BOPAlgo

is
    Create (S1,S2 : Shape from TopoDS)  
    	returns Cut from BRepAlgoAPI;  
	---Purpose: Shape aS2 cuts shape aS1. The
    	-- resulting shape is a new shape produced by the cut operation.
	

    Create (S1,S2 : Shape from TopoDS; 
    	    aDSF  : PaveFiller  from BOPAlgo; 
    	    bFWD  : Boolean from Standard=Standard_True)  
    	returns Cut from BRepAlgoAPI;	 
    	--- Purpose: Constructs a new shape cut from
    	-- shape aS1 by shape aS2 using aDSFiller (see
    	-- BRepAlgoAPI_BooleanOperation Constructor).
        
end Cut;
