-- File:        ManifoldSolidBrep.cdl
-- Created:     Mon Dec  4 12:02:27 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWManifoldSolidBrep from RWStepShape

	---Purpose : Read & Write Module for ManifoldSolidBrep

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     ManifoldSolidBrep from StepShape,
     EntityIterator from Interface

is

	Create returns RWManifoldSolidBrep;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable ManifoldSolidBrep from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : ManifoldSolidBrep from StepShape);

	Share(me; ent : ManifoldSolidBrep from StepShape; iter : in out EntityIterator);

end RWManifoldSolidBrep;
