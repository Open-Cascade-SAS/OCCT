-- Created on: 2005-12-15
-- Created by: Julia GERASIMOVA
-- Copyright (c) 2005-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class EigenValuesSearcher from math
        ---Purpose: This class finds eigen values and vectors of
        --          real symmetric tridiagonal matrix

uses 
     
    Array1OfReal  from TColStd, 
    HArray1OfReal from TColStd, 
    HArray2OfReal from TColStd, 
    Vector        from math
    
raises 
 
    NotDone from StdFail

is 
    Create(Diagonal    : Array1OfReal from TColStd; 
    	   Subdiagonal : Array1OfReal from TColStd)
    returns EigenValuesSearcher
    raises NotDone;  -- if length(Subdiagonal) != length(Diagonal)-1 
    
    IsDone(me)
     	---Purpose: Returns Standard_True if computation is performed 
        --          successfully.
    returns Boolean from Standard;

    Dimension(me)
     	---Purpose: Returns the dimension of matrix
    returns Integer from Standard;

    EigenValue(me; Index : Integer from Standard)
     	---Purpose: Returns the Index_th eigen value of matrix
        --          Index must be in [1, Dimension()]
    returns Real from Standard;

    EigenVector(me; Index : Integer from Standard)
     	---Purpose: Returns the Index_th eigen vector of matrix
        --          Index must be in [1, Dimension()]
    returns Vector from math;
     
fields 

    myDiagonal    : HArray1OfReal from TColStd;
    mySubdiagonal : HArray1OfReal from TColStd;  
    
    myIsDone       : Boolean from Standard; 
    myN            : Integer from Standard;
    myEigenValues  : HArray1OfReal from TColStd; 
    myEigenVectors : HArray2OfReal from TColStd;

end EigenValuesSearcher;
