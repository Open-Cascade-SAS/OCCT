-- File:	IGESDimen_ToolSectionedArea.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolSectionedArea  from IGESDimen

    ---Purpose : Tool to work on a SectionedArea. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses SectionedArea from IGESDimen,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolSectionedArea;
    ---Purpose : Returns a ToolSectionedArea, ready to work


    ReadOwnParams (me; ent : mutable SectionedArea;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : SectionedArea;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : SectionedArea;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a SectionedArea <ent>, from
    --           its specific (own) parameters

    DirChecker (me; ent : SectionedArea) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : SectionedArea;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : SectionedArea; entto : mutable SectionedArea;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : SectionedArea;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolSectionedArea;
