-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

package PShort 

uses PCollection,
     TCollection,
     TShort

is


--                             Instantiations de PCollection          --
--                             *****************************          --
------------------------------------------------------------------------

--
--       Instantiations HSequence 
--       **************************************************
--       
class HSequenceOfShortReal instantiates 
           HSequence from PCollection(ShortReal);

--
--       Instantiations HArray1
--       ****************************************************
--       
-----

    class HArray1OfShortReal instantiates 
                        HArray1 from PCollection(ShortReal);
--    class Array1FromHArray1OfShortReal instantiates 
--    	  Array1FromHArray1(ShortReal
--                           ,Array1OfShortReal from TShort
--                           ,HArray1OfShortReal from PShort);

--
--       Instantiations HArray2
--       ****************************************************
--       

    class HArray2OfShortReal instantiates 
                        HArray2 from PCollection(ShortReal);
--    class Array2FromHArray2OfShortReal instantiates 
--    	  Array2FromHArray2(ShortReal
--                           ,Array2OfShortReal from TShort
--                           ,HArray2OfShortReal from PShort);


end PShort;
