-- Created on: 1995-12-04
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package RWStepAP214 

uses

	StepData, Interface, TCollection, TColStd, StepAP214

is


class ReadWriteModule;

class GeneralModule;

class RWAutoDesignActualDateAndTimeAssignment;
class RWAutoDesignActualDateAssignment;
class RWAutoDesignApprovalAssignment;
class RWAutoDesignDateAndPersonAssignment;
class RWAutoDesignGroupAssignment;
class RWAutoDesignNominalDateAndTimeAssignment;
class RWAutoDesignNominalDateAssignment;
class RWAutoDesignOrganizationAssignment;
class RWAutoDesignPersonAndOrganizationAssignment;
class RWAutoDesignPresentedItem;
class RWAutoDesignSecurityClassificationAssignment;
-- Removed from Rev2 to Rev4 : class RWAutoDesignViewArea;

-- Added from STEP214-CC1 to CC2
class RWAutoDesignDocumentReference;
--Added from CC2 to DIS

class RWAppliedDateAndTimeAssignment;
class RWAppliedDateAssignment;
class RWAppliedApprovalAssignment;
class RWAppliedGroupAssignment;
class RWAppliedOrganizationAssignment;
class RWAppliedPersonAndOrganizationAssignment;
class RWAppliedPresentedItem;
class RWAppliedSecurityClassificationAssignment;
class RWAppliedDocumentReference;

-- added for external references (CAX-IF TRJ4)
class RWAppliedExternalIdentificationAssignment;
class RWClass;
class RWExternallyDefinedClass;
class RWExternallyDefinedGeneralProperty;
class RWRepItemGroup;

	Init;
	---Purpose: enforced the initialisation of the  libraries

end RWStepAP214;
