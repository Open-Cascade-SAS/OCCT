-- Created on: 1991-05-16
-- Created by: Isabelle GRIGNON
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class Int3Pln from IntAna 

	---Purpose: Intersection between 3 planes. The algorithm searches
	--          for an intersection point. If two of the planes are
	--          parallel or identical, IsEmpty returns TRUE.

uses Pln from gp,
     Pnt from gp

raises NotDone     from StdFail,
       DomainError from Standard

is

    Create
    
    	returns Int3Pln from IntAna;


    Create(P1,P2,P3 : Pln from gp)
    
    	---Purpose: Determination of the intersection point between
    	--          3 planes.

    	returns Int3Pln from IntAna;


    Perform(me: in out; P1,P2,P3 : Pln from gp)
    
    	---Purpose: Determination of the intersection point between
    	--          3 planes.

    	is static;


    IsDone(me)
    
	---Purpose: Returns True if the computation was successful.

    	returns Boolean from Standard
	---C++: inline
	is static;


    IsEmpty(me)
    
    	---Purpose: Returns TRUE if there is no intersection POINT.
    	--          If 2 planes are identical or parallel, IsEmpty
    	--          will return TRUE.

    	returns Boolean from Standard
	---C++: inline

	raises NotDone from StdFail
	--- The exception NotDone is raised when IsDone() returns False.
	is static;


    Value(me)
    
    	---Purpose: Returns the intersection point.

    	returns Pnt from gp
	---C++: inline
	---C++: return const&

   	raises NotDone     from StdFail,
               DomainError from Standard
	--- The exception NotDone is raised when IsDone() returns False.
	--- The exception Domain is raised when IsEmpty() returns False.
	
	is static;


fields

    done: Boolean from Standard;
    empt: Boolean from Standard;
    pnt : Pnt     from gp;

end Int3Pln;
