-- Created on: 1997-04-22
-- Created by: Guest Design
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MultipleConnectedInteractive from AIS inherits InteractiveObject from AIS

    
    ---Purpose: Defines an Interactive Object by gathering together
    -- several object presentations. This is done through a
    -- list of interactive objects. These can also be
    -- Connected objects. That way memory-costly
    -- calculations of presentation are avoided.
        
        
uses


    TypeOfPresentation3d   from PrsMgr,
    InteractiveObject      from AIS,
    Boolean                from Standard,
    SequenceOfInteractive  from AIS,
    KindOfInteractive      from AIS,
    PresentationManager3d  from PrsMgr,
    Presentation           from Prs3d,
    Projector             from Prs3d,
    Transformation        from Geom,
    Integer                from Standard,
    Selection              from SelectMgr,
    Trsf                  from gp

is 
    

    Create
    returns  MultipleConnectedInteractive  from  AIS;
    ---Purpose: Initializes the Interactive Object with multiple
    -- connections to AIS_Interactive objects.
    
    Connect(me             : mutable; 
    	    theInteractive : InteractiveObject from AIS);
    ---Purpose: Adds instance of theInteractive to child list.

    Connect(me:mutable;
            anotherIobj: InteractiveObject from AIS;
            aLocation : Trsf from gp) is virtual;
        ---Purpose: Establishes the connection between the Connected
        -- Interactive Object, anotherIobj, and its reference.
        -- Locates instance in aLocation.

    Type(me) returns KindOfInteractive from AIS
    is redefined virtual;	  

    Signature(me) returns Integer from Standard
    is redefined virtual;

    HasConnection(me) returns Boolean from Standard;
    ---Purpose: Returns true if the object is connected to others.
   
    Disconnect(me             : mutable;
    	       theInteractive : InteractiveObject from AIS);
    ---Purpose:  Removes the connection with theInteractive.

    DisconnectAll(me:mutable);
    ---Purpose: Clears all the connections to objects.
    
    Compute(me:mutable;
            aPresentationManager :         PresentationManager3d from PrsMgr;
            aPresentation        : Presentation          from Prs3d;
            aMode                :         Integer               from Standard = 0)
    ---Level: Internal 
    ---Purpose: this method is redefined virtual;
    --          when the instance is connected to another
    --          InteractiveObject,this method doesn't
    --          compute anything, but just uses the 
    --          presentation of this last object, with
    --          a transformation if there's one stored. 
    is redefined virtual protected; 

    Compute(me            : mutable;
    	    aProjector    : Projector from Prs3d;
    	    aTrsf         : Transformation from Geom;
	    aPresentation : Presentation from Prs3d)
    is redefined;
    ---Purpose: computes the presentation according to a point of view
    --          given by <aProjector>. 
    --          To be Used when the associated degenerated Presentations 
    --          have been transformed by <aTrsf> which is not a Pure
    --          Translation. The HLR Prs can't be deducted automatically
    --          WARNING :<aTrsf> must be applied
    --           to the object to display before computation  !!!

    Compute(me:mutable;
    	        aProjector: Projector from Prs3d;
                aPresentation: Presentation from Prs3d)
    is redefined ;

    AcceptShapeDecomposition(me) returns Boolean from Standard is redefined virtual;
        ---Purpose:  Informs the graphic context that the interactive Object
        -- may be decomposed into sub-shapes for dynamic selection.


    ComputeSelection(me:mutable; aSelection : Selection from SelectMgr;
                                 aMode      :        Integer   from Standard)
    is redefined virtual private;
        ---Purpose:  Computes the selection for whole subtree in scene hierarchy.



    
end MultipleConnectedInteractive;
