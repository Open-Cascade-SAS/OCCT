-- Created on: 1993-08-09
-- Created by: Didier PIFFAULT
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Circ from BRepMesh 

  ---Purpose: Describes  a  2d circle  with  a   size of  only 3
  --          Standard Real  numbers instead  of gp who  needs 7
  --          Standard Real numbers.

  uses    Real from Standard,
          XY from gp


  is      Create returns Circ from BRepMesh;

          Create (loc : XY from gp; rad : Real from Standard)
          returns Circ from BRepMesh;

          SetLocation(me : in out; loc : XY from gp)
          is static;

          SetRadius  (me : in out; rad : Real from Standard)
          is static;

          Location   (me)
          ---C++: return const &
          ---C++: inline
          returns XY from gp
          is static;

          Radius     (me)
          ---C++: return const &
          ---C++: inline
          returns Real from Standard
          is static;


fields  location : XY from gp;
        radius   : Real from Standard;

end Circ;
