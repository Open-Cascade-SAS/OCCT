-- Created by: Eugeny MALTCHIKOV
-- Copyright (c) 2013-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class EdgeEdge from IntTools 
    ---Purpose:   
    -- The class provides Edge/Edge intersection algorithm 
    -- based on the intersection between edges bounding boxes.

uses  
    Real  from Standard, 
    Box   from Bnd, 
    Range from IntTools, 
    Edge  from TopoDS,
    Curve from Geom,
    Curve from BRepAdaptor,
    ShapeEnum from TopAbs,  
    SequenceOfRanges from IntTools,
    SequenceOfCommonPrts from IntTools 
    
is  

    Create 
    returns EdgeEdge from IntTools; 
    ---C++: alias "~IntTools_EdgeEdge();"
    ---C++: inline 
    ---Purpose:  
    -- Empty contructor  
    
    Create ( 
        theEdge1 : Edge from TopoDS;  
        theEdge2 : Edge from TopoDS)  
    returns EdgeEdge from IntTools; 
    ---C++: inline 
    ---Purpose:  
    -- Contructor    
 
    Create ( 
        theEdge1   : Edge from TopoDS;  
        aT11, aT12 : Real from Standard;
        theEdge2   : Edge from TopoDS;  
        aT21, aT22 : Real from Standard)
    returns EdgeEdge from IntTools; 
    ---C++: inline
    ---Purpose:  
    -- Contructor    
    
    SetEdge1(me:out;  
        theEdge : Edge from TopoDS);
    ---C++: inline
    ---Purpose:  
    -- Sets the first edge
 
    SetEdge1(me:out;  
        theEdge : Edge from TopoDS; 
        aT1, aT2 : Real from Standard);
    ---C++: inline
    ---Purpose:  
    -- Sets the first edge and its range
    
    SetRange1(me:out;
        theRange1 : Range from IntTools);
    ---C++: inline
    ---Purpose:  
    -- Sets the range for the first edge
    
    SetRange1(me:out;
        aT1, aT2 : Real from Standard);
    ---C++: inline
    ---Purpose:  
    -- Sets the range for the first edge
    
    SetEdge2(me:out;  
        theEdge : Edge from TopoDS);
    ---C++: inline
    ---Purpose:  
    -- Sets the second edge 
     
    SetEdge2(me:out;  
        theEdge : Edge from TopoDS; 
        aT1, aT2 : Real from Standard);
    ---C++: inline
    ---Purpose:  
    -- Sets the first edge and its range
    
    SetRange2(me:out;
        theRange : Range from IntTools);
    ---C++: inline
    ---Purpose:  
    -- Sets the range for the second edge
    
    SetRange2(me:out;
        aT1, aT2 : Real from Standard);
    ---C++: inline
    ---Purpose:  
    -- Sets the range for the second edge  

    CheckData(me:out) 
    is protected; 
    ---C++: inline
    ---Purpose:  
    -- Checks the data

    Prepare(me:out) 
    is protected; 
    ---Purpose:  
    -- Prepares the data

    Perform(me:out); 
    ---Purpose:  
    -- Performs the intersection between edges
    
    ComputeLineLine(me:out)
    is protected;
    ---Purpose:
    -- Computes Line/Line intersection.  
 
    FindRoughRanges(me:out;
        theR1, theR2 : Range from IntTools; 
        theSegments1 : out SequenceOfRanges from IntTools)
    returns Integer from Standard 
    is protected; 
    ---Purpose: 
    -- Looking for the rough intersection ranges
 
    FindSolutions(me:out;  
        theRanges1 : out SequenceOfRanges from IntTools;
        theRanges2 : out SequenceOfRanges from IntTools)
    is protected; 
    ---Purpose:
    -- Looking for solutions

    FindSolutions(me:out;  
        theR1, theR2 : Range from IntTools;
        theBC        : Box from Bnd;
        theRanges1   : out SequenceOfRanges from IntTools;
        theRanges2   : out SequenceOfRanges from IntTools)
    is protected; 
    ---Purpose:
    -- Looking for the exact intersection ranges
    
    MergeSolutions(me:out; 
        theRanges1, theRanges2 : SequenceOfRanges from IntTools)
    is protected; 
    ---Purpose:
    -- Merges found solutions

    FindParameters(myclass; 
        theBAC  : Curve from BRepAdaptor;  
        aT1,aT2 : Real from Standard;  
        theRes  : Real from Standard;
        theCBox : Box from Bnd; 
        aTB1,aTB2 : out Real from Standard)
    returns Boolean from Standard 
    is protected; 
    ---Purpose:
    -- Looking for the range of the edge whick is in the box
     
    CheckCoincidence(me:out; 
        aT11, aT12  : Real from Standard; 
        aT21, aT22  : Real from Standard;  
        theCriteria : Real from Standard; 
        theCurveRes1: Real from Standard)
    returns Integer from Standard
    is protected;
    ---Purpose:  
    -- Checks if edges coincide on the ranges
     
    AddSolution(me:out; 
        aT11, aT12, aT21, aT22 : Real from Standard; 
        theType : ShapeEnum from TopAbs)
    is protected;
    ---Purpose:
    -- Adds common part of the given type to myCommonParts
     
    FindBestSolution(me:out; 
        aT11, aT12, aT21, aT22 : Real from Standard;  
        aT1, aT2 : out Real from Standard) 
    is protected;
    ---Purpose:
    -- Looking for the minimal distance between edges on the ranges
      
    IsIntersection(me:out; 
        aT11, aT12 : Real from Standard; 
        aT21, aT22 : Real from Standard)
    returns Boolean from Standard
    is protected;
    ---Purpose:  
    -- Checks is there an intersection between edges on the given ranges  
    -- (for nearly conicident edges)
    
    IsDone(me) 
    returns Boolean from Standard;
    ---C++: inline 
    ---Purpose: 
    -- Returns TRUE if common part(s) is(are) found
    
    CommonParts(me) 
    returns SequenceOfCommonPrts from IntTools;
    ---C++: inline 
    ---C++: return  const&   
    ---Purpose: 
    -- Returns common parts
    
fields  
    -- source data
    myEdge1  : Edge  from TopoDS is protected; 
    myEdge2  : Edge  from TopoDS is protected;  
    
    myGeom1  : Curve from Geom   is protected; 
    myGeom2  : Curve from Geom   is protected;  
    
    myCurve1 : Curve from BRepAdaptor is protected; 
    myCurve2 : Curve from BRepAdaptor is protected;  
    
    myTol1   : Real  from Standard is protected; 
    myTol2   : Real  from Standard is protected; 
    myTol    : Real  from Standard is protected;   
    
    myRes1   : Real  from Standard is protected;  
    myRes2   : Real  from Standard is protected; 
    
    myRange1 : Range from IntTools is protected; 
    myRange2 : Range from IntTools is protected;  
    
    -- results
    mySwap        : Boolean from Standard is protected; 
    myErrorStatus : Integer from Standard is protected; 
    myCommonParts : SequenceOfCommonPrts from IntTools is protected;
    
end EdgeEdge;
