-- Created on: 1997-08-04
-- Created by: Jean-Louis Frenkel
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ReferenceIterator from CDM

uses Document from CDM, ListIteratorOfListOfReferences from CDM
is

    Create(aDocument: Document from CDM);
    
    
    More(me) returns Boolean from Standard;
    
    
    Next(me: in out);
    
    
    Document(me) returns Document from CDM;
    
    ReferenceIdentifier(me) returns Integer from Standard;
    
    
    DocumentVersion(me) returns Integer from Standard;
    ---Purpose: returns the Document Version in the reference.
    
fields 
    myIterator: ListIteratorOfListOfReferences from CDM;
end ReferenceIterator from CDM;
    
    
