-- File:	QANewBRepNaming_BooleanOperation.cdl
-- Created:	Thu Nov 11 14:07:06 1999
-- Author:	Vladislav ROMASHKO
--		<vro@flox.nnov.matra-dtv.fr>
---Copyright:	 Matra Datavision 1999

 
class BooleanOperation from QANewBRepNaming inherits TopNaming from QANewBRepNaming

    ---Purpose: To load the BooleanOperation results
	
uses 
 
--modified by NIZNHY-PKV Wed Jun 19 09:06:12 2002  f  
    BooleanOperation from BRepAlgo,
    --BooleanOperation from BRepAlgoAPI, 
--modified by NIZNHY-PKV Wed Jun 19 09:06:16 2002  t    
    Shape            from TopoDS,
    Label            from TDF,
    ListOfShape      from TopTools

is
 
    Create returns BooleanOperation from QANewBRepNaming;

    Create(ResultLabel : Label from TDF) 
    returns BooleanOperation from QANewBRepNaming;

    Init(me : in out; ResultLabel :  Label from TDF);
	 
--modified by NIZNHY-PKV Wed Jun 19 09:06:46 2002  f	
    Load (me; mkBoolOp : in out BooleanOperation from BRepAlgo);
--    Load (me; mkBoolOp : in out BooleanOperation from BRepAlgoAPI); 
--modified by NIZNHY-PKV Wed Jun 19 09:06:53 2002  t 

    ---Purpose : Load the boolean operation.
    --           Makes a new part attached to the ResultLabel.

    FirstModified (me)
    ---Purpose: Returns the label of the modified faces
    --          of the first shape (S1).
    returns Label from TDF;  
    
    FirstDeleted (me)
    ---Purpose: Returns the label of the deleted faces
    --          of the first shape (S1).
    returns Label from TDF; 

    SecondModified (me)
    ---Purpose: Returns the label of the modified faces
    --          of the second shape (S2).
    returns Label from TDF;  
    
    SecondDeleted (me)
    ---Purpose: Returns the label of the deleted faces
    --          of the second shape (S2).
    returns Label from TDF; 
          
    Intersections (me)
    ---Purpose: Returns the label of intersections
    returns Label from TDF; 
     
end BooleanOperation;
