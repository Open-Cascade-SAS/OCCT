-- Created on: 1993-07-06
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class CurveOn2Surfaces from BRep inherits CurveRepresentation from BRep

	---Purpose: Defines a continuity between two surfaces.

uses
    Pnt      from gp,
    Surface  from Geom,
    Location from TopLoc,
    Shape    from GeomAbs,
    CurveRepresentation from BRep
    
raises
    NullObject from Standard
    
is

    Create(S1 , S2  : Surface  from Geom;
	   L1 , L2  : Location from TopLoc;
	   C        : Shape    from GeomAbs)
    returns mutable CurveOn2Surfaces from BRep;

    IsRegularity(me) returns Boolean
	---Purpose: Returns True.
    is redefined;
    
    IsRegularity(me; S1,S2 : Surface from Geom; 
                     L1,L2 : Location from TopLoc)  
    returns Boolean
	---Purpose: A curve on two surfaces (continuity). 
    is redefined;

    D0(me; U : Real; P : out Pnt from gp);
	---Purpose: Raises an error.
    
    Surface(me) returns any Surface from Geom
	---C++: return const &
    is redefined;

    Surface2(me) returns any Surface from Geom
	---C++: return const &
    is redefined;

    Location2(me) returns Location from TopLoc
	---C++: return const &
    is redefined;

    Continuity(me) returns Shape from GeomAbs
	---C++: return const &
    is redefined;
    
    Continuity(me : mutable; C : Shape from GeomAbs)
    is redefined;
    
    Copy(me) returns mutable CurveRepresentation from BRep;
	---Purpose: Return a copy of this representation.

fields
    mySurface    : Surface from Geom;
    mySurface2   : Surface from Geom;
    myLocation2  : Location from TopLoc;
    myContinuity : Shape from GeomAbs;

end CurveOn2Surfaces;
