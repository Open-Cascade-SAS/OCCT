-- Created on: 1993-01-11
-- Created by: CKY / Contract Toubro-Larsen (Niraj RANGWALA)
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package IGESDraw


        ---Purpose : This package contains the group of classes necessary for
        --           Structure Entities implied in Drawings and Structured
        --           Graphics (Sets for drawing, Drawings and Views).

uses

        Standard,
        TCollection,
        gp,
	TColgp,
	TColStd,
	Message,
        Interface,
        IGESData,
        IGESDimen,
        IGESBasic,
        IGESGraph,
        IGESGeom

is

     class ConnectPoint;

     class NetworkSubfigureDef;

     class ViewsVisible;

     class ViewsVisibleWithAttr;

     class LabelDisplay;

     class Planar;

     class SegmentedViewsVisible;

     class Drawing;

     class DrawingWithRotation;

     class View;

     class RectArraySubfigure;

     class CircArraySubfigure;

     class NetworkSubfigure;

     class PerspectiveView;

    	--    Tools for Entities    --

     class ToolConnectPoint;
     class ToolNetworkSubfigureDef;
     class ToolViewsVisible;
     class ToolViewsVisibleWithAttr;
     class ToolLabelDisplay;
     class ToolPlanar;
     class ToolSegmentedViewsVisible;
     class ToolDrawing;
     class ToolDrawingWithRotation;
     class ToolView;
     class ToolRectArraySubfigure;
     class ToolCircArraySubfigure;
     class ToolNetworkSubfigure;
     class ToolPerspectiveView;

     -- Definition and Exploitation of Entities defined in this Package

     class Protocol;
     class ReadWriteModule;
     class GeneralModule;
     class SpecificModule;

     -- The class instantiations :

     class  Array1OfConnectPoint   instantiates
    	  Array1 from TCollection (ConnectPoint);
     class  Array1OfViewKindEntity instantiates
          Array1 from TCollection (ViewKindEntity from IGESData);

     class HArray1OfConnectPoint   instantiates  HArray1 from TCollection
    	 (ConnectPoint,Array1OfConnectPoint);
     class HArray1OfViewKindEntity instantiates  HArray1 from TCollection
    	 (ViewKindEntity from IGESData,Array1OfViewKindEntity);

     -- Package Methods :

    Init;
    ---Purpose : Prepares dynamic data (Protocol, Modules) for this package

    Protocol  returns Protocol from IGESDraw;
    ---Purpose : Returns the Protocol for this Package

end IGESDraw;
