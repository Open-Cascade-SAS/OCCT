-- Created on: 1992-11-25
-- Created by: Jean Pierre TIRAULT
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


deferred class Array2Descriptor from TCollection

uses 
    Integer from Standard,
    Address from Standard

is
    Initialize (aLowerRow: Integer; aUpperRow: Integer; 
    	    	aLowerCol: Integer; aUpperCol: Integer;
    	    	anAddress: Address);

    UpperRow (me) returns Integer;
    ---Level: Advanced
    
    LowerRow (me) returns Integer;
    ---Level: Advanced

    UpperCol (me) returns Integer;
    ---Level: Advanced
    
    LowerCol (me) returns Integer;
    ---Level: Advanced

    Address(me) returns Address;
    ---Level: Advanced

fields
    myAddress     : Address;
    myLowerRow    : Integer;
    myLowerCol    : Integer;
    myUpperRow    : Integer;
    myUpperCol    : Integer;

    
end;    
