-- Created on: 2009-04-06
-- Created by: Sergey ZARITCHNY
-- Copyright (c) 2009-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Placement from TDataXtd inherits Attribute from TDF

	---Purpose: 

uses Attribute         from TDF,
     Label             from TDF,
     GUID              from Standard,
     Integer           from Standard,
     DataSet           from TDF,
     RelocationTable   from TDF,
     Constraint        from TDataXtd

is

    ---Purpose: class methods
    --          =============


    GetID (myclass)   
    	---C++: return const &  
    returns GUID from Standard;


    Set (myclass; label : Label from TDF)  
    ---Purpose: Find, or    create,   an Placement  attribute.     the
    --          Placement attribute is returned.
    returns Placement from TDataXtd;  
    

    ---Purpose: Placement methods
    --          =================


    Create
    returns mutable  Placement from TDataXtd;

    ---Category: TDF_Attribute methods
    --           =====================

    ID (me)
    	---C++: return const & 
    returns GUID from Standard;

    Restore (me: mutable; With : Attribute from TDF);

    NewEmpty (me)
    returns mutable Attribute from TDF;

    Paste (me; Into : mutable Attribute from TDF;
	       RT   : mutable RelocationTable from TDF);    

    Dump (me; anOS : in out OStream from Standard)
    	returns OStream from Standard
    	is redefined;
	---C++: return &

end Placement;

