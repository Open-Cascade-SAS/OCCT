-- Created on: 1993-02-22
-- Created by: Philippe DAUTRY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Hyperbola from PGeom inherits Conic from PGeom

        ---Purpose :Defines the main branch of an hyperbola.
        --         
	---See Also : Hyperbola from Geom.

uses Ax2 from gp

is


  Create returns mutable Hyperbola from PGeom;
        ---Purpose :Creates an Hyperbola with default values.
    	---Level: Internal 


  Create (aPosition : Ax2 from gp;
    	  aMajorRadius, aMinorRadius : Real from Standard)
     returns mutable Hyperbola from PGeom;
	---Purpose :  Creates an   Hyperbola    with      <aPosition>,
	--         <aMajorRadius> and  <aMinorRadius> as field values.
	--         The major  radius of the hyperbola is  on the XAxis
	--         and   the minor  radius is  on    the YAxis of  the
	--         hyperbola.
    	---Level: Internal 


  MajorRadius (me : mutable; aMajorRadius : Real from Standard);
	---Purpose: Set the value of the field majorRadius with <aMajorRadius>.
    	---Level: Internal 


  MajorRadius (me)  returns Real from Standard;
	---Purpose: Returns the value of the field majorRadius.
    	---Level: Internal 


  MinorRadius (me : mutable; aMinorRadius : Real from Standard);
	---Purpose: Set the value of the field minorRadius with <aMinorRadius>.
    	---Level: Internal 


  MinorRadius (me)  returns Real from Standard;
	---Purpose: Returns the value of the field minorRadius.
    	---Level: Internal 


fields

     majorRadius : Real from Standard;
     minorRadius : Real from Standard;

end;

