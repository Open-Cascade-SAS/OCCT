-- File:	StepBasic_ProductConceptContext.cdl
-- Created:	Fri Nov 26 16:26:39 1999 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0
-- Copyright:	Matra Datavision 1999

class ProductConceptContext from StepBasic
inherits ApplicationContextElement from StepBasic

    ---Purpose: Representation of STEP entity ProductConceptContext

uses
    HAsciiString from TCollection,
    ApplicationContext from StepBasic

is
    Create returns ProductConceptContext from StepBasic;
	---Purpose: Empty constructor

    Init (me: mutable; aApplicationContextElement_Name: HAsciiString from TCollection;
                       aApplicationContextElement_FrameOfReference: ApplicationContext from StepBasic;
                       aMarketSegmentType: HAsciiString from TCollection);
	---Purpose: Initialize all fields (own and inherited)

    MarketSegmentType (me) returns HAsciiString from TCollection;
	---Purpose: Returns field MarketSegmentType
    SetMarketSegmentType (me: mutable; MarketSegmentType: HAsciiString from TCollection);
	---Purpose: Set field MarketSegmentType

fields
    theMarketSegmentType: HAsciiString from TCollection;

end ProductConceptContext;
