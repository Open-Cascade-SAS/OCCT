-- Created on: 1997-12-09
-- Created by: Jean-Louis Frenkel
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

private class Reference from PCDM
uses ExtendedString from TCollection
is
    Create returns Reference from PCDM;
    
    Create(aReferenceIdentifier: Integer from Standard; aFileName: ExtendedString from TCollection; aDocumentVersion: Integer from Standard)
     returns Reference from PCDM;
    
    ReferenceIdentifier(me) returns Integer from Standard;
    
    FileName(me) returns ExtendedString from TCollection;
    
    DocumentVersion(me) returns Integer from Standard;
    
    
fields
    myReferenceIdentifier: Integer from Standard;
    myFileName: ExtendedString from TCollection;
    myDocumentVersion: Integer from Standard;
end Reference from PCDM;
