-- Created on: 1999-06-11
-- Created by: Vladislav ROMASHKO
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DriverTable from TFunction inherits TShared from MMgt
    	---Purpose: A container for instances of drivers.
    	-- You create a new instance of TFunction_Driver
    	-- and use the method AddDriver to load it into the driver table.
uses 
 
    DataMapOfGUIDDriver from TFunction, 
    Driver              from TFunction, 
    GUID                from Standard, 
    OStream             from Standard,
    DataMapOfGUIDDriver from TFunction,
    HArray1OfDataMapOfGUIDDriver from TFunction
    
is 

    Get (myclass)
    ---Purpose: Returns the driver table. If a driver does not exist, creates it.
    returns DriverTable from TFunction;

    Create returns DriverTable from TFunction; 
    ---Purpose: Default constructor

    AddDriver(me : mutable; guid   : GUID    from Standard;
    	    	    	    driver : Driver  from TFunction;
    	    	    	    thread : Integer from Standard = 0)
    ---Purpose: Returns true if the driver has been added successfully to the driver table.
    returns Boolean from Standard;

    HasDriver (me; guid   : GUID    from Standard;
    	    	   thread : Integer from Standard = 0)
    ---Purpose: Returns true if the driver exists in the driver table.
    returns Boolean from Standard;

    FindDriver(me; guid   :     GUID   from Standard; 
	 	   driver : out Driver from TFunction;
    	    	   thread :     Integer from Standard = 0)  
    ---Purpose: Returns true if the driver was found.
    returns Boolean from Standard;

    Dump(me; anOS : in out OStream from Standard) 
    ---C++: alias operator << 
    ---C++: return &
    returns OStream from Standard;

    RemoveDriver (me : mutable; guid   : GUID    from Standard;
    	    	    	    	thread : Integer from Standard = 0)
    ---Purpose: Removes a driver with the given GUID.
    --     Returns true if the driver has been removed successfully.
    returns Boolean from Standard;

    Clear (me : mutable);
    ---Purpose: Removes all drivers. Returns true if the driver has been removed successfully.

fields

    myDrivers       : DataMapOfGUIDDriver          from TFunction;
    myThreadDrivers : HArray1OfDataMapOfGUIDDriver from TFunction;

end DriverTable;   
