-- Created on: 1991-06-24
-- Created by: Christophe MARION
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- modified by mps (dec 96)  add of  ContinuityCommands



package GeometryTest 

	---Purpose: this  package  provides  commands for  curves  and
	--          surface.
uses
    Draw,
    Standard, 
    GeomliteTest

is

    AllCommands(I : in out Interpretor from Draw);
	---Purpose: defines all geometric commands.
    
    CurveCommands(I : in out Interpretor from Draw);
	---Purpose: defines curve commands.
    
    FairCurveCommands(I : in out Interpretor from Draw);
	---Purpose: defines fair curve commands.
    
    SurfaceCommands(I : in out Interpretor from Draw);
	---Purpose: defines surface commands.

    ConstraintCommands(I : in out Interpretor from Draw);
	---Purpose: defines cosntrained curves commands.
    
    API2dCommands(I : in out Interpretor from Draw);
	---Purpose: defines commands to test the Geom2dAPI
	--          - Intersection
	--          - Extrema
	--          - Projection
	--          - Approximation, interpolation
    
    APICommands(I : in out Interpretor from Draw);
	---Purpose: defines commands to test the Geom2dAPI
	--          - Intersection
	--          - Extrema
	--          - Projection
	--          - Approximation, interpolation
 
    ContinuityCommands(I : in out Interpretor from Draw);
        --- Purpose: defines commands to check local
        --          continuity between curves or surfaces

    PolyCommands(I : in out Interpretor from Draw);
	---Purpose: defines     command  to    test  the    polyhedral
	--          triangulations and the polygons from the Poly package.
    
    TestProjCommands(I : in out Interpretor from Draw);
	---Purpose: defines commands to test projection of geometric objects
    
end GeometryTest;
