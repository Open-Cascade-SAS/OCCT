-- Created on: 1993-01-09
-- Created by: CKY / Contract Toubro-Larsen ( Arun MENON )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class BasicDimension from IGESDimen   inherits IGESEntity
     
    ---Purpose: Defines IGES Basic Dimension, Type 406, Form 31,
    --          in package IGESDimen
    --          The basic Dimension Property indicates that the referencing 
    --          dimension entity is to be displayed with a box around text. 

uses

        Pnt2d       from gp,
        XY          from gp

is

        Create returns mutable BasicDimension;

            -- --specific-- --

        Init(me                    : mutable; 
             nbPropVal             : Integer;
             lowerLeft, lowerRight : XY;
             upperRight, upperLeft : XY); 
        -- This method is used to set the fields of the
        -- class BasicDimension
        --       - nbPropVal  : Number of property values
        --       - lowerLeft  : Coordinates of lower left corner
        --       - lowerRight : Coordinates of lower right corner
        --       - upperRight : Coordinates of upper right corner
        --       - upperLeft  : Coordinates of upper left corner

        NbPropertyValues(me) returns Integer;
        ---Purpose : returns the number of properties = 8

        LowerLeft(me) returns Pnt2d;
        ---Purpose : returns coordinates of lower left corner

        LowerRight(me) returns Pnt2d;
        ---Purpose : returns coordinates of lower right corner

        UpperRight(me) returns Pnt2d;
        ---Purpose : returns coordinates of upper right corner

        UpperLeft(me) returns Pnt2d;
        ---Purpose : returns coordinates of upper left corner

fields

--
-- Class    : IGESDimen_BasicDimension
-- 
-- Purpose  : Declaration of variables specific to the definition
--            of the Class BasicDimension.
--
-- Reminder : A BasicDimension instance is defined by :
--                - The number of property values, always 8
--                - Coordinates of lower left corner
--                - Coordinates of lower right corner
--                - Coordinates of upper right corner
--                - Coordinates of upper left corner
--
--

        theNbPropertyValues : Integer;
        theLowerLeft        : XY;
        theLowerRight       : XY;
        theUpperRight       : XY;
        theUpperLeft        : XY;

end BasicDimension;
