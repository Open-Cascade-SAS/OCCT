-- Created on: 2005-10-05
-- Created by: Mikhail KLOKOV
-- Copyright (c) 2005-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class CurveRangeSample from IntTools inherits BaseRangeSample from IntTools
    ---Purpose: class for range index management of curve

uses
    Range from IntTools
is

    Create
    	returns CurveRangeSample from IntTools;

    Create(theIndex: Integer from Standard)
    	returns CurveRangeSample from IntTools;

    SetRangeIndex(me: in out; theIndex: Integer from Standard);
	---C++: inline

    GetRangeIndex(me)
    	returns Integer from Standard;
	---C++: inline
	
    IsEqual(me; Other: CurveRangeSample from IntTools)
    	returns Boolean from Standard;
	---C++: inline

    GetRange(me; theFirst, theLast: Real from Standard; 
    	    	 theNbSample: Integer from Standard)
    	returns Range from IntTools;

    GetRangeIndexDeeper(me; theNbSample: Integer from Standard)
    	returns Integer from Standard;
	---C++: inline

fields
    myIndex: Integer from Standard;

end CurveRangeSample from IntTools;
