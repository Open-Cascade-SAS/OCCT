-- Created on: 1996-09-10
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class DrawableSUR from TestTopOpeDraw inherits Surface from DrawTrSurf

uses 
    
    Surface     from Geom,
    Color           from Draw,
    Display         from Draw,
    Text3D          from Draw,
    CString         from Standard,
    Pnt             from gp,
    Pnt2d           from gp

is 

    Create (S : Surface from Geom; IsoColor : Color from Draw)
    returns mutable DrawableSUR from TestTopOpeDraw;

    Create (S : Surface from Geom; IsoColor : Color from Draw;
    	    Text : CString from Standard; TextColor : Color from Draw)
    returns mutable DrawableSUR from TestTopOpeDraw;

    Create (S : Surface from Geom; IsoColor : Color from Draw;
            BoundColor,NormalColor : Color from Draw;
    	    Text : CString from Standard; TextColor : Color from Draw;
	    Nu,Nv : Integer;
    	    Discret : Integer; Deflection : Real; DrawMode : Integer;
    	    DispOrigin : Boolean from Standard = Standard_True)
    returns mutable DrawableSUR from TestTopOpeDraw;

    Pnt(me) returns Pnt from gp
    is static;

    Pnt2d(me) returns Pnt2d from gp
    is static;
    
    DrawOn(me; dis : in out Display from Draw)
    is redefined;

    NormalColor(me : mutable; NormalColor : Color from Draw)
    is static;

    DrawNormale(me; dis : in out Display from Draw)
    is static;
    
fields

    myText : Text3D from Draw;
    myNormalColor : Color from Draw;
    
end DrawableSUR;
