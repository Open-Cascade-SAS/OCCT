-- Created on: 1993-08-05
-- Created by: Martine LANGLOIS
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MakeBSplineSurfaceWithKnots from GeomToStep  
    inherits Root from GeomToStep
    
    ---Purpose: This class implements the mapping between class
    --          BSplineSurface from Geom and the class
    --          BSplineSurfaceWithKnots from  
    --          StepGeom which describes a 
    --          bspline_Surface_with_knots from Prostep
  
uses BSplineSurface from Geom,
     BSplineSurfaceWithKnots from StepGeom
     
raises NotDone from StdFail
     
is 

Create ( Bsplin : BSplineSurface from Geom ) returns
    MakeBSplineSurfaceWithKnots;

Value (me) returns
    BSplineSurfaceWithKnots from StepGeom
    raises NotDone
    is static;
    ---C++: return const&

fields

    theBSplineSurfaceWithKnots :
    	BSplineSurfaceWithKnots from StepGeom;
    	-- The solution from StepGeom
    	
end MakeBSplineSurfaceWithKnots;


