-- Created on: 1993-07-02
-- Created by: Laurent BUCHARD
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

generic class SurfaceTool from IntCurveSurface 
    ( TheSurface       as any)
                                 
				 
uses 
   
   Shape        from GeomAbs,
   SurfaceType  from GeomAbs,
   Pln          from gp,
   Cone         from gp,
   Cylinder     from gp,
   Sphere       from gp,
   Torus        from gp, 
   Pnt          from gp,
   Vec          from gp,
   Array1OfReal from TColStd,
   BezierSurface   from Geom,
   BSplineSurface  from Geom,
   HSurface     from Adaptor3d,
   HCurve       from Adaptor3d,
   Ax1          from gp,
   Dir          from gp

raises 
   NoSuchObject from Standard,
   OutOfRange   from Standard


is 
  
    FirstUParameter(myclass; S: TheSurface)
        ---C++: inline
        returns Real from Standard;
	
    FirstVParameter(myclass; S: TheSurface)
        ---C++: inline
        returns Real from Standard;

    LastUParameter(myclass; S: TheSurface)
        ---C++: inline
        returns Real from Standard;

    LastVParameter(myclass; S: TheSurface)
        ---C++: inline
        returns Real from Standard;



    NbUIntervals(myclass; S: TheSurface;
    	    	          Sh : Shape from GeomAbs)
    	---C++: inline
    	returns Integer from Standard;

    NbVIntervals(myclass; S: TheSurface;
    	    	    	  Sh : Shape from GeomAbs) 
    	---C++: inline 
        returns Integer from Standard;



    UIntervals(myclass; S  : TheSurface;
    	    	    	T  : in out Array1OfReal from TColStd; 
    	    	    	Sh : Shape from GeomAbs);
    	---C++: inline

    VIntervals(myclass; S  : TheSurface;
    	    	    	T  : in out Array1OfReal from TColStd; 
    	    	    	Sh : Shape from GeomAbs) ;
    	---C++: inline 


   UTrim(myclass; S : TheSurface;
                  First, Last, Tol : Real) 
	---C++: inline
    returns HSurface from Adaptor3d
    raises
    	OutOfRange from Standard;
	---Purpose: If <First> >= <Last> 
    
   VTrim(myclass; S : TheSurface;
                  First, Last, Tol : Real) 
	---C++: inline
    returns HSurface from Adaptor3d
    raises
    	OutOfRange from Standard;
	---Purpose: If <First> >= <Last> 
    

    IsUClosed(myclass; S: TheSurface) 
    	---C++: inline
    	returns Boolean from Standard;

    IsVClosed(myclass; S: TheSurface) 
    	---C++: inline
    	returns Boolean from Standard;
    

    IsUPeriodic(myclass; S: TheSurface) 
    	---C++: inline
    	returns Boolean from Standard;

    UPeriod(myclass; S: TheSurface) 
    	---C++: inline
    	returns Real from Standard;
	
    IsVPeriodic(myclass; S: TheSurface) 
    	---C++: inline
    	returns Boolean from Standard;
    
    VPeriod(myclass; S: TheSurface) 
    	---C++: inline
    	returns Real from Standard;
	


    Value(myclass; S   : TheSurface;
    	           u,v : Real from Standard)
	---C++: inline
	returns Pnt from gp;

    D0(myclass; S   : TheSurface; 
                u,v : Real from Standard;
		P   : out Pnt from gp);
    	---C++: inline 

    D1(myclass; S      : TheSurface; 
                u,v    : Real from Standard; 
                P      : out Pnt from gp;
                D1u,D1v: out Vec from gp); 
    	---C++: inline 
    	
    D2(myclass; S      : TheSurface; 
                u,v    : Real from Standard; 
                P      : out Pnt from gp;
                D1U,D1V,D2U,D2V,D2UV: out Vec from gp); 
    	---C++: inline 
    	
    D3(myclass; S      : TheSurface; 
                u,v    : Real from Standard; 
                P      : out Pnt from gp;
                D1U, D1V, D2U, D2V, D2UV, D3U, D3V, D3UUV, D3UVV: out Vec from gp); 
    	---C++: inline 
    	
    DN(myclass; S      : TheSurface; 
                u,v    : Real from Standard; 
                Nu,Nv  : Integer from Standard)
    	---C++: inline 
    returns Vec from gp;
	


    UResolution(myclass; S:TheSurface; R3d: Real from Standard) 
        ---C++: inline
        returns Real from Standard;

    VResolution(myclass; S:TheSurface; R3d: Real from Standard)
        ---C++: inline
        returns Real from Standard;

    GetType(myclass; S: TheSurface)
    	---C++: inline
    	returns SurfaceType from GeomAbs;


    Plane(myclass; S: TheSurface) 
    	---C++: inline
    	returns Pln from gp;
        
    Cylinder(myclass; S : TheSurface) returns Cylinder from gp
      raises NoSuchObject from Standard;
    	---C++: inline

    
    Cone(myclass; S : TheSurface) returns Cone from gp
      raises NoSuchObject from Standard;
    	---C++: inline

    Torus(myclass; S : TheSurface) returns Torus from gp    
      raises NoSuchObject from Standard;
    	---C++: inline


    Sphere(myclass; S : TheSurface) returns Sphere from gp
      raises NoSuchObject from Standard;
    	---C++: inline

    Bezier(myclass; S : TheSurface) returns BezierSurface from  Geom
      raises NoSuchObject from Standard;
    	---C++: inline

    BSpline(myclass; S : TheSurface) returns BSplineSurface  from  Geom
      raises NoSuchObject from Standard;
    	---C++: inline
    
    AxeOfRevolution(myclass; S: TheSurface) returns Ax1 from  gp 
      raises NoSuchObject from Standard;
        ---C++: inline

    Direction(myclass; S: TheSurface) returns Dir from gp
      raises NoSuchObject from Standard;
        ---C++: inline

    BasisCurve(myclass; S:TheSurface) returns HCurve from Adaptor3d 
      raises NoSuchObject from Standard;
        ---C++: inline
  

--------------------------------------------------------------------------------


    NbSamplesU(myclass; S : TheSurface) returns Integer from Standard; 

       
    NbSamplesV(myclass; S : TheSurface) returns Integer from Standard;    


    NbSamplesU(myclass; S : TheSurface; u1,u2: Real from Standard) returns Integer from Standard; 

       
    NbSamplesV(myclass; S : TheSurface; v1,v2: Real from Standard) returns Integer from Standard;    



end SurfaceTool;
