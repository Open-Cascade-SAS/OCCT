-- Created by: Peter KURNEV
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package BOPCol 

 ---Purpose:  
     -- The package contains collection classes 
     -- that are used by  
     -- partition and  boolean operation algorithms     
uses 
    TCollection
 
is 
    imported BaseAllocator from BOPCol; 
    imported DataMapOfShapeInteger from BOPCol; 
    imported DataMapOfShapeReal from BOPCol; 
    imported MapOfInteger from BOPCol; 
    imported ListOfInteger from BOPCol; 
    imported PInteger from BOPCol; 
    imported DataMapOfIntegerInteger from BOPCol; 
    imported DataMapOfIntegerReal from BOPCol; 
    imported DataMapOfIntegerListOfInteger from BOPCol; 
    imported IndexedDataMapOfShapeBox from BOPCol; 
    imported IndexedMapOfInteger from BOPCol; 
    imported ListOfShape from BOPCol;   
    imported DataMapOfShapeAddress from BOPCol;   
    imported DataMapOfTransientAddress from BOPCol;   
    imported PListOfInteger from BOPCol;  
    imported MapOfShape from BOPCol;  
    imported DataMapOfShapeShape from BOPCol;  
    imported DataMapOfShapeListOfShape from BOPCol;  
    imported MapOfOrientedShape from BOPCol;  
    imported IndexedDataMapOfShapeListOfShape from BOPCol;  
    imported IndexedMapOfShape from BOPCol;  
    imported ListOfListOfShape from BOPCol;  
    imported SequenceOfShape from BOPCol;  
    imported SequenceOfPnt2d from BOPCol;  
    imported DataMapOfIntegerListOfShape from BOPCol;
    imported IndexedDataMapOfIntegerListOfInteger from BOPCol;
    imported IndexedDataMapOfShapeInteger from BOPCol;  
   
    
end BOPCol;
