-- Created on: 1992-05-13
-- Created by: NW,JPB,CAL
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class GenId from Aspect

  ---Purpose: This class permits the creation and control of integer identifiers.

uses

  ListOfInteger from TColStd

raises

  IdentDefinitionError from Aspect

is

  Create
  returns GenId from Aspect;
  ---Purpose: Creates an available set of identifiers with the lower bound 0 and the upper bound INT_MAX / 2.

  Create (theLow, theUpper : Integer from Standard)
  returns GenId from Aspect
  ---Purpose: Creates an available set of identifiers with specified range.
  -- Raises IdentDefinitionError if theUpper is less than theLow.
  raises IdentDefinitionError from Aspect;

  Free (me : in out);
  ---Level: Internal
  ---Purpose: Free all identifiers - make the whole range available again.

  Free (me    : in out;
        theId : Integer from Standard);
  ---Purpose: Free specified identifier. Warning - method has no protection against double-freeing!

  HasFree (me)
  returns Boolean from Standard;
  ---Purpose: Returns true if there are available identifiers in range.

  Available (me)
  returns Integer from Standard;
  ---Purpose: Returns the number of available identifiers.

  Lower (me)
  returns Integer from Standard;
  ---Purpose: Returns the lower identifier in range.

  Next (me : in out)
  returns Integer from Standard
  ---Purpose: Returns the next available identifier.
  -- Warning: Raises IdentDefinitionError if all identifiers are busy.
  raises IdentDefinitionError from Aspect;

  Upper (me)
  returns Integer from Standard;
  ---Purpose: Returns the upper identifier in range.

fields

  myFreeCount  : Integer from Standard;      -- the current number of available identifiers in range, excluding freed numbers
  myLength     : Integer from Standard;      -- the number of identifiers
  myLowerBound : Integer from Standard;      -- the lower limit for identifiers
  myUpperBound : Integer from Standard;      -- the upper limit for identifiers
  myFreeIds    : ListOfInteger from TColStd; -- to save free identifiers

end GenId;
