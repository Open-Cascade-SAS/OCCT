-- Created on: 1992-05-22
-- Created by: Jean Claude VAUTHIER
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class BezierCurve2d


from DrawTrSurf


inherits Curve2d from DrawTrSurf


uses BezierCurve from Geom2d,
     Color from Draw,
     Display from Draw,
     Drawable3D from Draw


is


  Create (C : BezierCurve from Geom2d)
        --- Purpose :
        --  creates a drawable Bezier curve from a Bezier curve of 
        --  package Geom2d.
     returns mutable BezierCurve2d from DrawTrSurf;


  Create (C : BezierCurve from Geom2d;
          CurvColor, PolesColor : Color from Draw;
          ShowPoles : Boolean; Discret : Integer)
     returns mutable BezierCurve2d from DrawTrSurf;


  DrawOn (me; dis : in out Display from Draw)
     is redefined static;


  ShowPoles (me : mutable)
     is static;


  ClearPoles (me : mutable)
     is static;
     
  
  FindPole(me; X,Y : Real; D : Display from Draw; Prec : Real; 
           Index : in out Integer)
        --- Purpose :
        --  Returns in <Index> the index of the first pole  of the
        --  curve projected by the Display <D> at a distance lower
        --  than <Prec> from <X,Y>. If no pole  is found  index is
        --  set to 0, else index is always  greater than the input
        --  value of index.
  is static;
  
  
  SetPolesColor (me : mutable; aColor : Color from Draw)
        ---C++: inline
     is static;

  PolesColor (me)  returns Color from Draw
        ---C++: inline
     is static;
    
  Copy(me) returns mutable Drawable3D from Draw
	---Purpose: For variable copy.
  is redefined;
  
      
fields

  drawPoles  : Boolean;
  polesLook  : Color from Draw;

end BezierCurve2d;
