-- Created on: 1996-01-10
-- Created by: Denis PASCAL
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class PlanarDistance from DrawDim inherits PlanarDimension from DrawDim

	---Purpose: PlanarDistance point/point
	--          PlanarDistance point/line
	--          PlanarDistance line/line

uses Face    from TopoDS,
     Pnt     from gp,
     Shape   from TopoDS,
     Edge    from TopoDS,
     Color   from Draw,
     Display from Draw

is

    Create (plane  : Face from TopoDS;
            point1 : Shape from TopoDS;
            point2 : Shape from TopoDS)
    returns mutable PlanarDistance from DrawDim;
    
    Create (geom1 : Shape from TopoDS;
            geom2 : Shape from TopoDS)
    returns mutable PlanarDistance from DrawDim; 
    
    DrawOn(me; dis : in out Display);

    ---Purpose: private
    Draw (me; p : Pnt from gp;
              e : Edge from TopoDS;
              d : in out Display) is private;
    
fields

    myGeom1 : Shape from TopoDS;
    myGeom2 : Shape from TopoDS;
    
end PlanarDistance;
