-- Created on: 1998-01-07
-- Created by: Philippe MANGIN
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred  class SectionLaw from BRepFill  inherits TShared from MMgt

	---Purpose: Build Section Law, with an Vertex, or an Wire
        ---Level: Advanced
       
uses 
 SectionLaw          from GeomFill,  
 HArray1OfSectionLaw from  GeomFill, 
 Shape               from  GeomAbs, 
 Shape               from  TopoDS,
 Wire                from  TopoDS,  
 Edge                from  TopoDS, 
 Vertex              from  TopoDS,  
 WireExplorer        from  BRepTools 
  
 
is  
  NbLaw(me)  returns  Integer;  
   
  Law(me; Index  :  Integer)  
   ---C++: return const &
    returns SectionLaw from GeomFill; 
     
  IsConstant(me)  returns  Boolean 
  is  deferred; 
  
  IsUClosed(me)  returns  Boolean; 
   
  IsVClosed(me)  returns  Boolean; 
   
  IsVertex(me) 
    ---Purpose: Say if the input sahpe is a  vertex. 
  returns  Boolean   
  is  deferred;   
   
  ConcatenedLaw(me)  
  returns SectionLaw from GeomFill 
  is  deferred;        

  Continuity(me; Index  :  Integer; 
    	         TolAngular  :  Real)
  returns  Shape  from  GeomAbs 
  is  deferred;  
   
  VertexTol(me; Index  :  Integer;   
                Param  :  Real) 
  returns  Real 
  is  deferred; 	   
  
  Vertex(me;  Index  :  Integer; 
              Param  :  Real) 
  returns Vertex  from  TopoDS 
  is deferred;	 
   
  D0(me:mutable;  U  :  Real;   
     S  :  out  Shape  from  TopoDS) 
  is  deferred;  
   
  Init(me:  mutable;  W  :  Wire  from  TopoDS);  
       
  
  CurrentEdge(me  :  mutable)   
  returns  Edge  from  TopoDS;   
  
fields  
  myLaws      :  HArray1OfSectionLaw from  GeomFill is  protected; 
  uclosed     :  Boolean       from  Standard is  protected;  
  vclosed     :  Boolean       from  Standard is  protected;   
  myIterator  :  WireExplorer  from  BRepTools;  
end SectionLaw;
