-- Created on: 1993-03-10
-- Created by: JCV
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



deferred class Curve from Geom inherits Geometry from Geom

    	---Purpose : The abstract class Curve describes the common
    	-- behavior of curves in 3D space. The Geom package
    	-- provides numerous concrete classes of derived
    	-- curves, including lines, circles, conics, Bezier or
    	-- BSpline curves, etc.
    	-- The main characteristic of these curves is that they
    	-- are parameterized. The Geom_Curve class shows:
    	-- - how to work with the parametric equation of a curve
    	--   in order to calculate the point of parameter u,
    	--   together with the vector tangent and the derivative
    	--   vectors of order 2, 3,..., N at this point;
    	-- - how to obtain general information about the curve
    	--   (for example, level of continuity, closed
    	--   characteristics, periodicity, bounds of the parameter field);
    	-- - how the parameter changes when a geometric
    	--   transformation is applied to the curve or when the
    	--   orientation of the curve is inverted.
    	--   All curves must have a geometric continuity: a curve is
    	--   at least "C0". Generally, this property is checked at
    	-- the time of construction or when the curve is edited.
    	-- Where this is not the case, the documentation states so explicitly.
    	-- Warning
    	-- The Geom package does not prevent the
    	-- construction of curves with null length or curves which
    	-- self-intersect.
       

uses Pnt   from gp,
     Vec   from gp,
     Trsf  from gp,
     Shape from GeomAbs

raises RangeError          from Standard,
       NoSuchObject        from Standard,
       UndefinedDerivative from Geom,
       UndefinedValue      from Geom


is


  Reverse (me : mutable) 
        ---Purpose :
        --  Changes the direction of parametrization of <me>. 
        --  The "FirstParameter" and the "LastParameter" are not changed
        --  but the orientation  of the curve is modified. If the curve
        --  is bounded the StartPoint of the initial curve becomes the
        --  EndPoint of the reversed curve  and the EndPoint of the initial
        --  curve becomes the StartPoint of the reversed curve.
     is deferred;  
     
  ReversedParameter(me; U : Real) returns Real
	---Purpose: Returns the  parameter on the  reversed  curve for
	--          the point of parameter U on <me>.
	--          
	--          me->Reversed()->Value(me->ReversedParameter(U))
	--          
	--          is the same point as
	--          
	--          me->Value(U)
     is deferred;  

  TransformedParameter(me; U : Real; T : Trsf from gp) returns Real
	---Purpose: Returns the  parameter on the  transformed  curve for
	--          the transform of the point of parameter U on <me>.
	--          
	--          me->Transformed(T)->Value(me->TransformedParameter(U,T))
	--          
	--          is the same point as
	--          
	--          me->Value(U).Transformed(T)
	--          
	--          This methods returns <U>
	--          
	--          It can be redefined. For example on the Line.
     is virtual;  


  ParametricTransformation(me; T : Trsf from gp) returns Real
	---Purpose: Returns a  coefficient to compute the parameter on
	--          the transformed  curve  for  the transform  of the
	--          point on <me>.
	--          
	--          Transformed(T)->Value(U * ParametricTransformation(T))
	--          
	--          is the same point as
	--          
	--          Value(U).Transformed(T)
	--          
	--          This methods returns 1.
	--          
	--          It can be redefined. For example on the Line.
     is virtual;  


  Reversed (me)  returns mutable like me 
        ---Purpose : Returns a copy of <me> reversed.
     is static;


  FirstParameter (me)   returns Real
        ---Purpose : Returns the value of the first parameter.
        --  Warnings :
        --  It can be RealFirst from package Standard 
        --  if the curve is infinite
     is deferred;


  LastParameter (me)   returns Real
        ---Purpose :  Returns the value of the last parameter.
        --  Warnings :
        --  It can be RealLast from package Standard 
        --  if the curve is infinite
     is deferred;


  IsClosed (me)   returns Boolean
        ---Purpose : Returns true if the curve is closed.
        --  Some curves such as circle are always closed, others such as line
        --  are never closed (by definition).
        --  Some Curves such as OffsetCurve can be closed or not. These curves
        --  are considered as closed if the distance between the first point
        --  and the last point of the curve is lower or equal to the Resolution
        --  from package gp wich is a fixed criterion independant of the
        --  application.
     is deferred;


  IsPeriodic (me)  returns Boolean
        ---Purpose : Is the parametrization of the curve periodic ?
        --  It is possible only if the curve is closed and if the
        --  following relation is satisfied :
        --  for each parametric value U the distance between the point
        --  P(u) and the point P (u + T) is lower or equal to Resolution
        --  from package gp, T is the period and must be a constant.
        --  There are three possibilities :
        --   . the curve is never periodic by definition (SegmentLine)
        --   . the curve is always periodic by definition (Circle)
        --   . the curve can be defined as periodic (BSpline). In this case
        --     a function SetPeriodic allows you to give the shape of the
        --     curve.  The general rule for this case is : if a curve can be 
        --     periodic or not the default periodicity set is non periodic
        --     and you have to turn (explicitly) the curve into a periodic 
        --     curve  if you want the curve to be periodic.
     is deferred;


  Period (me)   returns Real from Standard
	---Purpose: Returns the period of this curve.
    	-- Exceptions Standard_NoSuchObject if this curve is not periodic.
  raises
    	NoSuchObject from Standard
  is virtual;


  Continuity (me)   returns Shape from GeomAbs
        ---Purpose : It is the global continuity of the curve 
        --  C0 : only geometric continuity,
        --  C1 : continuity of the first derivative all along the Curve,
        --  C2 : continuity of the second derivative all along the Curve,
        --  C3 : continuity of the third derivative all along the Curve,
        --  G1 : tangency continuity all along the Curve,
        --  G2 : curvature continuity all along the Curve,
        --  CN : the order of continuity is infinite.
     is deferred;

  IsCN (me; N : Integer)  returns Boolean
        ---Purpose : Returns true if the degree of continuity of this curve is at least N.
    	-- Exceptions -  Standard_RangeError if N is less than 0.
     raises RangeError
     is deferred;


  D0(me; U : Real; P : out Pnt)
	---Purpose: Returns in P the point of parameter U.
        --  If the curve is periodic  then the returned point is P(U) with 
        --  U = Ustart + (U - Uend)  where Ustart and Uend are the 
        --  parametric bounds of the curve.
     raises  UndefinedValue
        ---Purpose :
        --  Raised only for the "OffsetCurve" if it is not possible to 
        --  compute the current point. For example when the first 
        --  derivative on the basis curve and the offset direction
        --  are parallel.
     is deferred;


  D1 (me; U : Real; P : out Pnt; V1 : out Vec)
        ---Purpose :
        --  Returns the point P of parameter U and the first derivative V1.
     raises UndefinedDerivative
        ---Purpose : Raised if the continuity of the curve is not C1.
     is deferred;


  D2 (me; U : Real; P : out Pnt; V1, V2 : out Vec)
        ---Purpose :
        --  Returns the point P of parameter U, the first and second
        --  derivatives V1 and V2.
     raises UndefinedDerivative
        ---Purpose : Raised if the continuity of the curve is not C2.
     is deferred;


  D3 (me; U : Real; P : out Pnt; V1, V2, V3 : out Vec)
        ---Purpose :
        --  Returns the point P of parameter U, the first, the second 
        --  and the third derivative.
     raises UndefinedDerivative
        ---Purpose : Raised if the continuity of the curve is not C3.
     is deferred;
        

  DN (me; U : Real; N : Integer)   returns Vec
        ---Purpose :
    	-- The returned vector gives the value of the derivative for the 
        --  order of derivation N.
     raises  UndefinedDerivative,
    	---Purpose : Raised if the continuity of the curve is not CN.
        --         
    	---Purpose :  Raised if the   derivative  cannot  be  computed
        --         easily. e.g. rational bspline and n > 3.
             RangeError
        ---Purpose : Raised if N < 1.            
     is deferred;


  Value (me; U : Real)    returns Pnt 
        ---Purpose : Computes the point of parameter U on <me>.
    	--  If the curve is periodic  then the returned point is P(U) with 
    	--  U = Ustart + (U - Uend)  where Ustart and Uend are the 
        --  parametric bounds of the curve.
        --  it is implemented with D0.
     raises  UndefinedValue
        ---Purpose :
    	--  Raised only for the "OffsetCurve" if it is not possible to 
        --  compute the current point. For example when the first
     	--  derivative on the basis curve and the offset direction are parallel.
     is static;


end;







