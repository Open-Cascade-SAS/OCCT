-- Created on: 1999-07-12
-- Created by: Denis PASCAL
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

private class Modified from TDocStd inherits Attribute from TDF

    ---Purpose:   Transient     attribute   wich     register modified
    --          labels. This attribute is attached to root label.


uses Label           from TDF,
     Attribute       from TDF,
     LabelMap        from TDF,
     RelocationTable from TDF


is

    ---Purpose: API class methods
    --          =================

    IsEmpty (myclass; access : Label from TDF)
    returns Boolean;   

    Add (myclass; alabel : Label from TDF)
    returns Boolean;    

    Remove (myclass; alabel : Label from TDF)
    returns Boolean;    

    Contains (myclass; alabel : Label from TDF)
    returns Boolean;

    Get (myclass; access : Label from TDF)
    ---Purpose: if <IsEmpty> raise an exception.
    ---C++: return const &
    returns LabelMap from TDF;

    Clear (myclass; access : Label from TDF);
    ---Purpose: remove all modified labels. becomes empty

    GetID (myclass)   
    ---C++: return const &  
    returns GUID from Standard;

    ---Purpose: Modified methods
    --          ================
    
    Create
    returns Modified from TDocStd;  
    
    IsEmpty (me)
    returns Boolean from Standard;    

    Clear (me : mutable);

    AddLabel (me : mutable; L : Label from TDF)
    ---Purpose: add <L> as modified 
    returns Boolean from Standard;

    RemoveLabel (me : mutable; L : Label from TDF)    
    ---Purpose: remove  <L> as modified 
    returns Boolean from Standard;
    
    Get (me)  
    ---Purpose: returns modified label map
    ---C++: return const & 
    returns LabelMap from TDF; 
        
    ---Category: methodes de TDF_Attribute
    --           =========================
    
    ID (me)
    ---C++: return const & 
    returns GUID from Standard;

    Restore (me: mutable; With : Attribute from TDF);

    NewEmpty (me)
    returns Attribute from TDF;

    Paste (me; Into : Attribute from TDF;
	       RT   : RelocationTable from TDF);    

    Dump (me; anOS : in out OStream from Standard)
    returns OStream from Standard
    is redefined;
    ---C++: return &

fields

    myModified : LabelMap from TDF;

end Modified;
