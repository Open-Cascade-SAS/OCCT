-- Created on: 1992-06-30
-- Created by: Laurent BUCHARD
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package IntAna

    ---Purpose: This package provides the intersections between :
    --          
    --          - Natural Quadrics when the result is a conic (QuadQuadGeo)
    --          
    --          - A natural Quadric and a Quadric defined by its Coefficients
    --            (IntQuadQuad)
    --            
    --          - 3 Pln   (Int3Pln)
    --          
    --          - a Line and a Torus   (IntLinTorus)
    --          
    --          - a Conic from gp and  a Quadric  defined by its Coefficients
    --            (IntConicQuad)
    --            

    ---Level: Public
    --
    -- All the methods of the classes of this package are public.
    --

  
uses TCollection, math, gp, StdFail, IntAna2d, GeomAbs

is

    enumeration ResultType  is Point,
                               Line,
                               Circle,
                               PointAndCircle,
                               Ellipse,
                               Parabola,
                               Hyperbola,
                               Empty,
			       Same,
                               NoGeometricSolution;
    

    
    class QuadQuadGeo;
    
    class IntQuadQuad;

    class Int3Pln;

    class IntLinTorus;
    
    class IntConicQuad;

    class Curve;
    
    class Quadric;
    --
    class ListOfCurve  instantiates  
    	List from TCollection(Curve from IntAna);    
    --
end IntAna;


 
