-- Created on: 1993-03-23
-- Created by: BBL
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class EuclidAlienData from AlienImage inherits AlienImageData from AlienImage

	---Version: 0.0

	---Level: Public
	---Purpose: This class defines an Euclid .PIX Alien image.
	---Keywords:
	---Warning:
	---References:

uses
	File 			from OSD,
	AsciiString 		from TCollection,
	ColorImage 		from Image,
	PseudoColorImage 	from Image,
	Image			from Image,
	HArray2OfInteger	from TColStd

raises
	OutOfRange 	from Standard,
	TypeMismatch 	from Standard

is
	Create returns mutable EuclidAlienData from AlienImage ;

	Clear( me : in out mutable ) ;
	---Level: Public
	---Purpose: Frees memory allocated by EuclidAlienData
	---C++: alias ~

	Read ( me : in out mutable ; afile : in out File from OSD )
	  returns Boolean from Standard ;
	---Level: Public
	  ---Purpose: Read content of a  EuclidAlienData object from a file .
	  --          Returns True if file is a XWD file .

	Write( me : in immutable; afile : in out File from OSD )
	  returns Boolean from Standard ;
	---Level: Public
	  ---Purpose: Write content of a  EuclidAlienData object to a file .

	ToImage( me : in  immutable) 
	  returns mutable Image from Image 
          raises TypeMismatch from Standard ;
	---Level: Public
	  ---Purpose : convert a EuclidAlienData object to a Image object.

	FromImage( me : in out mutable ; anImage : in Image from Image )
          raises TypeMismatch from Standard ;
	---Level: Public
	  ---Purpose : convert a Image object to a EuclidAlienData object.

	--
	--			Private Method
	--


	FromPseudoColorImage( me : in out mutable ; 
			      anImage : in PseudoColorImage from Image );
	---Level: Internal
	  ---Purpose : convert a Image object to a EuclidAlienData object.

	FromColorImage( me : in out mutable ; 
				anImage : in ColorImage from Image );
	---Level: Internal
	  ---Purpose : convert a Image object to a EuclidAlienData object.

fields

	myX1, myY1, myX2, myY2 	: Integer from Standard ;
	myNumberOfColor 	: Integer from Standard ;
	myColors 		: Address from Standard ;
	myPixels 		: HArray2OfInteger from TColStd ;
	myPixelsIsDef		: Boolean from Standard ;
end ;
 
