-- Created on: 1993-03-23
-- Created by: BBL,JLF
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class XWD from ImageUtility

	---Version: 0.0

	---Purpose: Performs a "xwd" and creates a XAlienImage and an Image

	---Keywords:
	---Warning:
	---References:

uses
	XAlienImage	from AlienImage,
	File		from OSD,
	Image 		from Image

raises
	TypeMismatch 	from Standard

is
	Create returns XWD from ImageUtility ;
	---Level: Internal
	---Purpose: Create a XWD object .

	XWD( me : in out ; xwdOptions : CString from Standard = "" )
		returns Boolean from Standard
		is static;
	---Level: Internal
	---Purpose: execute a Spawn "xwd xwudOptions -out aTmpFile" .

	XAlienImage( me )
		returns XAlienImage from AlienImage
		is static;
	---Level: Internal
	---Purpose: returns the XAlienImage created from "xwd".

	Image( me )
		returns Image from Image
		is static;
	---Level: Internal
	---Purpose: returns the Image created from "xwd".

fields
	myXAlienImage : XAlienImage from AlienImage;
	myImage : Image		from Image;
end ;
