-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ProductDefinition from StepBasic 

inherits TShared from MMgt

uses

	HAsciiString from TCollection, 
	ProductDefinitionFormation from StepBasic, 
	ProductDefinitionContext from StepBasic
is

	Create returns ProductDefinition;
	---Purpose: Returns a ProductDefinition

	Init (me : mutable;
	      aId : HAsciiString from TCollection;
	      aDescription : HAsciiString from TCollection;
	      aFormation : ProductDefinitionFormation from StepBasic;
	      aFrameOfReference : ProductDefinitionContext from StepBasic) is virtual;

	-- Specific Methods for Field Data Access --

	SetId(me : mutable; aId : HAsciiString);
	Id (me) returns HAsciiString;
	SetDescription(me : mutable; aDescription : HAsciiString);
	Description (me) returns HAsciiString;
	SetFormation(me : mutable; aFormation : ProductDefinitionFormation);
	Formation (me) returns ProductDefinitionFormation;
	SetFrameOfReference(me : mutable; aFrameOfReference : ProductDefinitionContext);
	FrameOfReference (me) returns ProductDefinitionContext;

fields

	id : HAsciiString from TCollection;
	description : HAsciiString from TCollection;
	formation : ProductDefinitionFormation from StepBasic;
	frameOfReference : ProductDefinitionContext from StepBasic;

end ProductDefinition;
