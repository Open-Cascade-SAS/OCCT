-- Created on: 1991-10-02
-- Created by: NW,JPB,CAL
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Background from Aspect


	---Purpose: This class allows the definition of
	--	    a window background.

uses

	Color	from Quantity

is

	Create
		returns Background from Aspect;
	---Level: Public
	---Purpose: Creates a window background.
	--	    Default color : NOC_MATRAGRAY.

	Create ( AColor : Color from Quantity )
		returns Background from Aspect;
	---Level: Public
	---Purpose: Creates a window background with the colour <AColor>.

	---------------------------------------------------
	-- Category: Methods to modify the class definition
	---------------------------------------------------

	SetColor ( me		: in out;
		   AColor	: Color from Quantity );
	---Level: Public
	---Purpose: Modifies the colour of the window background <me>.
	---Category: Methods to modify the class definition

	----------------------------
	-- Category: Inquire methods
	----------------------------

	Color ( me )
		returns Color from Quantity;
	---Level: Public
	---Purpose: Returns the colour of the window background <me>.
	---Category: Inquire methods

--

fields

--
-- Class	:	Aspect_Background
--
-- Purpose	:	Declaration of variables specific to the window
--			background.
--
-- Reminder	:	A background is defined by one colour
--

	-- the colour associated with the window background
	MyColor	:	Color from Quantity;

end Background;
