-- Created on: 1995-03-28
-- Created by: Yves FRICAUD
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Substitution from BRepTools 

	---Purpose: A tool to substitute subshapes by other shapes.
	--          
    	--          
    	--          The user use the method Substitute to define the
    	--          modifications. 
    	--          A set of shapes is designated to replace a initial
    	--          shape. 
    	--
    	--          The method Build reconstructs a new Shape with the
    	--          modifications.The Shape and the new shape are 
    	--          registered.
    	--          

uses
    Shape                     from TopoDS,
    ListOfShape               from TopTools,	
    DataMapOfShapeListOfShape from TopTools
    
raises
    
    NoSuchObject from Standard
is
    
    Create returns Substitution from BRepTools;
    
    Clear ( me : in out)
    	---Purpose: Reset all the fields.
    is static;

    Substitute (me : in out; 
    	    	OldShape  : Shape from TopoDS;
    	    	NewShapes : ListOfShape from TopTools)
    	---Purpose: <Oldshape> will be replaced by <NewShapes>.
    	--          
    	--          <NewShapes> can be empty , in this case <OldShape>
    	--          will disparate from its ancestors.
    	--          
    	--          if an item of <NewShapes> is oriented FORWARD.
    	--          it will be oriented as <OldShape> in its ancestors.
    	--          else it will be reversed.
    is static;
    
    
    Build (me : in out; S : Shape from TopoDS)
	---Purpose: Build NewShape from <S> if its subshapes has modified.
	--          
	--          The methods <IsCopied> and <Copy> allows you to keep
	--          the resul of <Build>
    is static;	    
    
    IsCopied(me; S : Shape from TopoDS) returns Boolean
	---Purpose: Returns   True if <S> has   been  replaced .
    is static;
    
    Copy(me; S : Shape from TopoDS) returns ListOfShape from TopTools
	---Purpose: Returns the set of shapes  substitued to <S> .
	---C++: return const &
    raises
    	NoSuchObject from Standard -- if ! IsCopied(S)
    is static;
    
fields

    myMap    : DataMapOfShapeListOfShape from TopTools;
    
end Substitution;
