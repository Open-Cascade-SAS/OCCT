-- Created on: 1993-04-26
-- Created by: Jean-Louis Frenkel
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

--   GG  : GER61351 17/11/1999 Change SetColor() with a compatible Quantity_Color instead
--				       the restricted NameOfColor.
--			  Parameters the color model rule (not especially the front & back side)
--			  Add the SetTransparency() method.
--			  Add the Color(),Material() and Transparency() methods


class ShadingAspect from Prs3d inherits BasicAspect from Prs3d
    	---Purpose: A framework to define the display of shading.
    	-- The attributes which make up this definition include:
    	-- -   fill aspect
    	-- -   color, and
    	-- -   material
uses 

    TypeOfFacingModel	   from Aspect,
    AspectFillArea3d       from Graphic3d,
    NameOfColor            from Quantity,
    Color			   from Quantity,
    NameOfMaterial   from Graphic3d,
    --NameOfMaterialPhysic   from Graphic3d,
    MaterialAspect         from Graphic3d,
    TypeOfLine             from Aspect

is
    Create
    	---Purpose: Constructs an empty framework to display shading.
    returns ShadingAspect from Prs3d;
    
    SetColor (me: mutable; aColor: Color from Quantity;
				   aModel: TypeOfFacingModel from Aspect = Aspect_TOFM_BOTH_SIDE)
    is static;
    	--- Purpose: Change the polygons interior color and material ambient color.

    SetColor (me: mutable; aColor: NameOfColor from Quantity;
		  		   aModel: TypeOfFacingModel from Aspect = Aspect_TOFM_BOTH_SIDE)
    is static;
    	--- Purpose: Change the polygons interior color and material ambient color.
    	
    SetMaterial(me: mutable; aMaterial: MaterialAspect from Graphic3d;
				     aModel: TypeOfFacingModel from Aspect = Aspect_TOFM_BOTH_SIDE)
    is static;
    	--- Purpose: Change the polygons material aspect.

    SetMaterial(me: mutable; aMaterial: NameOfMaterial from Graphic3d;
				     aModel: TypeOfFacingModel from Aspect = Aspect_TOFM_BOTH_SIDE)
    is static;

    SetTransparency(me: mutable; aValue: Real from Standard;
				         aModel: TypeOfFacingModel from Aspect = Aspect_TOFM_BOTH_SIDE)
    is static;
    	--- Purpose: Change the polygons transparency value.
    	--  Warning : aValue must be in the range 0,1. 0 is the default (NO transparent)

    SetAspect(me:mutable; Asp : AspectFillArea3d from Graphic3d);
    	--- Purpose: Change the polygons aspect properties.

    Color (me; aModel: TypeOfFacingModel from Aspect = Aspect_TOFM_FRONT_SIDE) 
    returns Color from Quantity is static;
    	--- Purpose: Returns the polygons color.

    Material (me; aModel: TypeOfFacingModel from Aspect = Aspect_TOFM_FRONT_SIDE) 
    returns MaterialAspect from Graphic3d is static;
    	--- Purpose: Returns the polygons material aspect.

    Transparency (me; aModel: TypeOfFacingModel from Aspect = Aspect_TOFM_FRONT_SIDE) 
    returns Real from Standard is static;
    	--- Purpose: Returns the polygons transparency value.

    Aspect (me) returns AspectFillArea3d from Graphic3d;
    	--- Purpose: Returns the polygons aspect properties.
    
fields

    myAspect: AspectFillArea3d from Graphic3d;

end ShadingAspect from Prs3d;
