-- File:        SphericalSurface.cdl
-- Created:     Mon Dec  4 12:02:31 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWSphericalSurface from RWStepGeom

	---Purpose : Read & Write Module for SphericalSurface

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     SphericalSurface from StepGeom,
     EntityIterator from Interface

is

	Create returns RWSphericalSurface;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable SphericalSurface from StepGeom);

	WriteStep (me; SW : in out StepWriter; ent : SphericalSurface from StepGeom);

	Share(me; ent : SphericalSurface from StepGeom; iter : in out EntityIterator);

end RWSphericalSurface;
