-- Created on: 1999-12-20
-- Created by: data exchange team
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MakeTriangulation from ShapeConstruct  inherits MakeShape from BRepBuilderAPI

	---Purpose: 

uses

    Array1OfPnt from TColgp,
    Wire from TopoDS

is

    Create (pnts : Array1OfPnt from TColgp; prec : Real = 0.0)
    returns MakeTriangulation from ShapeConstruct;

    Create (wire : Wire from TopoDS; prec : Real = 0.0)
    returns MakeTriangulation from ShapeConstruct;

    Build (me : in out) is redefined;

    IsDone (me) returns Boolean is redefined;

    Triangulate (me : in out; wire : Wire from TopoDS) is private;

    AddFacet (me : in out; wire : Wire from TopoDS) is private;

fields

    myPrecision : Real from Standard;
    myWire      : Wire from TopoDS;

end MakeTriangulation;
