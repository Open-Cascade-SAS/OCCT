-- Created on: 1998-06-03
-- Created by: data exchange team
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class ReShape from ShapeBuild inherits ReShape from BRepTools

    ---Purpose: Rebuilds a Shape by making pre-defined substitutions on some
    --          of its components
    --
    --          In a first phase, it records requests to replace or remove
    --          some individual shapes
    --          For each shape, the last given request is recorded
    --          Requests may be applied "Oriented" (i.e. only to an item with
    --          the SAME orientation) or not (the orientation of replacing
    --          shape is respectful of that of the original one)
    --           
    --          Then, these requests may be applied to any shape which may
    --          contain one or more of these individual shapes

uses 
    ShapeEnum from TopAbs, 
    Shape     from TopoDS,
    Status from ShapeExtend

is

    Create returns mutable ReShape from ShapeBuild;
    	---Purpose: Returns an empty Reshape

    Apply (me: mutable; shape: Shape from TopoDS; until: ShapeEnum from TopAbs; buildmode: Integer)
    returns Shape from TopoDS is redefined;
    	---Purpose: Applies the substitutions requests to a shape
    	--         
    	--          <until> gives the level of type until which requests are taken
    	--          into account. For subshapes of the type <until> no rebuild 
        --          and futher exploring are done.
    	--          ACTUALLY, NOT IMPLEMENTED BELOW  TopAbs_FACE
    	--           
    	--          <buildmode> says how to do on a SOLID,SHELL ... if one of its
    	--          sub-shapes has been changed:
    	--          0: at least one Replace or Remove -> COMPOUND, else as such
    	--          1: at least one Remove (Replace are ignored) -> COMPOUND
    	--          2: Replace and Remove are both ignored
    	--          If Replace/Remove are ignored or absent, the result as same
    	--          type as the starting shape

    Apply (me: mutable; shape: Shape from TopoDS; until: ShapeEnum from TopAbs = TopAbs_SHAPE)
    returns Shape from TopoDS is redefined;
    	---Purpose: Applies the substitutions requests to a shape.
    	--         
    	--          <until> gives the level of type until which requests are taken
    	--          into account. For subshapes of the type <until> no rebuild 
        --          and futher exploring are done.
	--
	--          NOTE: each subshape can be replaced by shape of the same type
	--          or by shape containing only shapes of that type (for 
	--          example, TopoDS_Edge can be replaced by TopoDS_Edge,
	--          TopoDS_Wire or TopoDS_Compound containing TopoDS_Edges).
	--          If incompatible shape type is encountered, it is ignored
	--          and flag FAIL1 is set in Status.
    
    Status (me: mutable; shape: Shape from TopoDS; newsh: out Shape from TopoDS; last : Boolean = Standard_False)
    returns Integer is redefined;
    	---Purpose: Returns a complete substitution status for a shape
    	--          0  : not recorded,   <newsh> = original <shape>
    	--          < 0: to be removed,  <newsh> is NULL
    	--          > 0: to be replaced, <newsh> is a new item
	--          If <last> is False, returns status and new shape recorded in
	--          the map directly for the shape, if True and status > 0 then
	--          recursively searches for the last status and new shape.

    Status (me; status: Status from ShapeExtend) returns Boolean;
    	---Purpose: Queries the status of last call to Apply(shape,enum)
    	--          OK   : no (sub)shapes replaced or removed
    	--          DONE1: source (starting) shape replaced
    	--          DONE2: source (starting) shape removed
    	--          DONE3: some subshapes replaced
    	--          DONE4: some subshapes removed
    	--          FAIL1: some replacements not done because of bad type of subshape

end ReShape;
