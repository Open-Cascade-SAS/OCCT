-- Created on: 1995-04-25
-- Created by: Marie Jose MARTZ
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



package BRepToIGESBRep

    ---Purpose : Provides tools in order to transfer CAS.CADE entities
    --         to IGESBRep.

uses 
    Interface,
    IGESData,
    IGESBasic,
    IGESGeom,
    IGESSolid,
    Geom,
    Geom2d,
    GeomAbs,
    GeomToIGES,
    Geom2dToIGES,
    TColStd,
    TopoDS,
    TopTools,
    TopLoc,
    TopAbs,
    Transfer,
    TransferBRep,
    BRep,
    BRepTools, 
    gp,
    TCollection,
    BRepToIGES

is

--  ------------------------------------------------------
--  Package Classes
--  ------------------------------------------------------

    class Entity;


end BRepToIGESBRep;
