-- Created on: 1996-09-23
-- Created by: Philippe MANGIN
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Modified:	Fri Jul 10 11:23:35 1998
--              JCT : Add WithRatio,MinM


class CompCurveToBSplineCurve from GeomConvert 

	---Purpose: Concat several curve in an BSplineCurve

uses
 ParameterisationType from Convert,
 BoundedCurve from Geom,
 BSplineCurve from Geom

--raises

is

    Create(Parameterisation : ParameterisationType from Convert =  Convert_TgtThetaOver2);
    ---Purpose: Initialize the algorithme
    --        - Parameterisation is used to convert


    Create (BasisCurve : BoundedCurve from Geom; 
     	    Parameterisation : ParameterisationType from Convert 
    	    	       =  Convert_TgtThetaOver2)
	 ---Purpose: Initialize the algorithme with one curve
	 --        - Parameterisation is used to convert 
    returns CompCurveToBSplineCurve;
    

    Add (me : in out; 
         NewCurve   :  BoundedCurve from Geom;
         Tolerance  :  Real from Standard;
         After      :  Boolean from Standard = Standard_False; 
         WithRatio  :  Boolean from Standard = Standard_True; 
         MinM       :  Integer  from  Standard  =  0)
	---Purpose: Append a curve in  the BSpline Return False if the
	--          curve is not G0  with the BSplineCurve.  Tolerance
	--             is   used to   check   continuity  and decrease
	--          Multiplicity at the common Knot until MinM
	--          if MinM = 0, the common Knot can be removed
    returns Boolean;
       
    
    Add (me : in out; 
         FirstCurve : in out BSplineCurve from Geom;
    	 SecondCurve: in out BSplineCurve from Geom;
         After      : Boolean from Standard; 
         WithRatio  : Boolean from Standard; 
         MinM       : Integer from Standard)
	---Purpose: Concat two BSplineCurves.
    	is private;    
    
    BSplineCurve(me) returns BSplineCurve from Geom;

    Clear(me : in out);
    ---Purpose: Clear a result curve

fields
 myCurve :  BSplineCurve from Geom;
 myTol   :  Real;
 myType  :  ParameterisationType from Convert;

end CompCurveToBSplineCurve;
