-- Created on: 1994-12-09
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class NurbsConvert from BRepBuilderAPI inherits ModifyShape from BRepBuilderAPI

	---Purpose: Conversion of the complete geometry of a shape into
    	-- NURBS geometry. For example, all curves supporting
    	-- edges of the basis shape are converted into BSpline
    	-- curves, and all surfaces supporting its faces are
    	-- converted into BSpline surfaces.

uses 

    Shape             from TopoDS,
    Face              from TopoDS,
    ShapeModification from BRepBuilderAPI,
    ListOfShape       from TopTools
     
is

    Create returns NurbsConvert from BRepBuilderAPI;
    	---Purpose: Constructs a framework for converting the geometry of a
    	-- shape into NURBS geometry. Use the function Perform
    	-- to define the shape to convert.
    Create(S: Shape from TopoDS; 
           Copy: Boolean from Standard  =  Standard_False)

    	returns NurbsConvert from BRepBuilderAPI;
	---Purpose:  Builds a new shape by converting the geometry of the
    	-- shape S into NURBS geometry. Specifically, all curves
    	-- supporting edges of S are converted into BSpline
    	-- curves, and all surfaces supporting its faces are
    	-- converted into BSpline surfaces.
    	-- Use the function Shape to access the new shape.
    	-- Note: the constructed framework can be reused to
    	-- convert other shapes. You specify these with the
    	-- function Perform.

    Perform(me: in out; S   : Shape   from TopoDS; 
                        Copy: Boolean from Standard  =  Standard_False)

	---Purpose: Builds a new shape by converting the geometry of the
    	-- shape S into NURBS geometry.
    	-- Specifically, all curves supporting edges of S are
    	-- converted into BSpline curves, and all surfaces
    	-- supporting its faces are converted into BSpline surfaces.
    	-- Use the function Shape to access the new shape.
    	-- Note: this framework can be reused to convert other
    	-- shapes: you specify them by calling the function Perform again.
    	is static;

end NurbsConvert;
