-- File:	RWStepFEA_RWNodeSet.cdl
-- Created:	Thu Dec 12 17:51:06 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWNodeSet from RWStepFEA

    ---Purpose: Read & Write tool for NodeSet

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    NodeSet from StepFEA

is
    Create returns RWNodeSet from RWStepFEA;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : NodeSet from StepFEA);
	---Purpose: Reads NodeSet

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: NodeSet from StepFEA);
	---Purpose: Writes NodeSet

    Share (me; ent : NodeSet from StepFEA;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWNodeSet;
