-- Created on: 1995-02-01
-- Created by: Marie Jose MARTZ
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Geom2dCurve from Geom2dToIGES inherits Geom2dEntity from Geom2dToIGES

    ---Purpose: This class implements the transfer of the Curve Entity from Geom2d
    --          To IGES. These can be :
    --          Curve
    --            . BoundedCurve
    --               * BSplineCurve
    --               * BezierCurve
    --               * TrimmedCurve
    --            . Conic     
    --               * Circle
    --               * Ellipse
    --               * Hyperbloa
    --               * Line
    --               * Parabola
    --            . OffsetCurve     
  

uses

    Curve                from Geom2d,
    BoundedCurve         from Geom2d,
    BSplineCurve         from Geom2d,
    BezierCurve          from Geom2d,
    TrimmedCurve         from Geom2d,
    Conic                from Geom2d,
    Circle               from Geom2d,
    Ellipse              from Geom2d,
    Hyperbola            from Geom2d,
    Line                 from Geom2d,
    Parabola             from Geom2d,
    OffsetCurve          from Geom2d,
    IGESEntity           from IGESData,
    Geom2dEntity         from Geom2dToIGES
    
    
is 
    
    Create returns Geom2dCurve from Geom2dToIGES;


    Create(G2dE : Geom2dEntity from Geom2dToIGES)  
    	 returns Geom2dCurve from Geom2dToIGES;
    ---Purpose : Creates a tool Geom2dCurve ready to run and sets its
    --         fields as G2dE's.

    Transfer2dCurve (me    : in out;
                     start : Curve from Geom2d;
		     Udeb  : Real  from Standard;
		     Ufin  : Real  from Standard)
    	 returns mutable IGESEntity from IGESData;
    ---Purpose :  Transfert  an Entity from Geom2d to IGES. If this
    --            Entity could not be converted, this member returns a NullEntity.

end Geom2dCurve;


