-- Created on: 1998-10-19
-- Created by: Christian CAILLET
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class SelectSuite  from IFSelect    inherits SelectDeduct  from IFSelect

    ---Purpose : A SelectSuite can describe a suite of SelectDeduct as a unique
    --           one : in other words, it can be seen as a "macro selection"
    --           
    --           It works by applying each of its items (which is a
    --           SelectDeduct) on the result computed by the previous one
    --           (by using Alternate Input)
    --           
    --           But each of these Selections used as items may be used
    --           independently, it will then give its own result
    --           
    --           Hence, SelectSuite gives a way of defining a new Selection
    --           from existing ones, without having to do copies or saves

uses CString, AsciiString from TCollection,
     SequenceOfTransient from TColStd,
     Graph from Interface, EntityIterator from Interface,
     Selection from IFSelect

raises InterfaceError

is

    Create returns SelectSuite;
    ---Purpose : Creates an empty SelectSuite

    AddInput (me : mutable; item : Selection) returns Boolean;
    ---Purpose : Adds an input selection. I.E. :
    --           If <item> is a SelectDeduct, adds it as Previous, not as Input
    --           Else, sets it as Input
    --           Returns True when done
    --           Returns False and refuses to work if Input is already defined

    AddPrevious (me : mutable; item : SelectDeduct);
    ---Purpose : Adds a new first item (prepends to the list). The Input is not
    --           touched
    --           If <item> is null, does nothing

    AddNext     (me : mutable; item : SelectDeduct);
    ---Purpose : Adds a new last item (prepends to the list)
    --           If <item> is null, does nothing

    NbItems (me) returns Integer;
    ---Purpose : Returns the count of Items

    Item    (me; num : Integer) returns SelectDeduct;
    ---Purpose : Returns an item from its rank in the list
    --           (the Input is always apart)

    SetLabel (me : mutable; lab : CString);
    ---Purpose : Sets a value for the Label

    	--  Definitions for Selecting

    RootResult (me; G : Graph) returns EntityIterator
        raises InterfaceError;
    ---Purpose : Returns the list of selected entities
    --           To do this, once InputResult has been taken (if Input or
    --           Alternate has been defined, else the first Item gives it) :
    --           this result is set as alternate input for the first item,
    --           which computes its result : this result is set as alternate
    --           input for the second item, etc...

    Label (me) returns AsciiString from TCollection;
    ---Purpose : Returns the Label
    --           Either it has been defined by SetLabel, or it will give
    --           "Suite of nn Selections"

fields

    thelab : AsciiString;
    thesel : SequenceOfTransient;

end SelectSuite;
