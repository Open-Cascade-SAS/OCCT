-- Created on: 1998-04-07
-- Created by: Jean-Pierre COMBE
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- modified     Sergey Zaritchny

class Position from PDataXtd inherits Attribute from PDF

	---Purpose: Position of a Label

uses Pnt from gp

is

    Create returns Position from PDataXtd;
    
    GetPosition (me)
    ---C++: inline
    returns Pnt from gp;
    
    SetPosition (me: mutable ; aPosition : Pnt from gp);
    ---C++: inline

fields

    myPosition : Pnt  from gp;	
    
end Position;

