-- File:	StepAP214_ExternalIdentificationItem.cdl
-- Created:	Wed May 10 15:09:05 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class ExternalIdentificationItem from StepAP214
inherits SelectType from StepData

    ---Purpose: Representation of STEP SELECT type ExternalIdentificationItem

uses
    DocumentFile from StepBasic,
    ExternallyDefinedClass from StepAP214,
    ExternallyDefinedGeneralProperty from StepAP214,
    ProductDefinition from StepBasic

is
    Create returns ExternalIdentificationItem from StepAP214;
	---Purpose: Empty constructor

    CaseNum (me; ent: Transient) returns Integer;
	---Purpose: Recognizes a kind of ExternalIdentificationItem select type
	--          1 -> DocumentFile from StepBasic
	--          2 -> ExternallyDefinedClass from StepAP214
	--          3 -> ExternallyDefinedGeneralProperty from StepAP214
	--          4 -> ProductDefinition from StepBasic
	--          0 else

    DocumentFile (me) returns DocumentFile from StepBasic;
	---Purpose: Returns Value as DocumentFile (or Null if another type)

    ExternallyDefinedClass (me) returns ExternallyDefinedClass from StepAP214;
	---Purpose: Returns Value as ExternallyDefinedClass (or Null if another type)

    ExternallyDefinedGeneralProperty (me) returns ExternallyDefinedGeneralProperty from StepAP214;
	---Purpose: Returns Value as ExternallyDefinedGeneralProperty (or Null if another type)

    ProductDefinition (me) returns ProductDefinition from StepBasic;
	---Purpose: Returns Value as ProductDefinition (or Null if another type)

end ExternalIdentificationItem;
