-- Created on: 1996-01-29
-- Created by: Kernel
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class BaseArray from DBC
inherits Storable from Standard

uses DBVArray from DBC

raises NullObject,
    NegativeValue,
    DimensionMismatch

is
    Create returns BaseArray;
    ---Purpose: Creates an BaseArray of NULL size
    
    Create (Size : Integer) returns BaseArray;
    ---Purpose: Creates  an BaseArray of lower bound 0 and
    --          upper bound <Size>-1.

    Create (BaseArray: BaseArray) returns BaseArray;
    ---Purpose: Creates an array which  is the copy of the given
    --          argument.

    Delete ( me : out ) is redefined;
    ---C++: alias "Standard_EXPORT virtual ~DBC_BaseArray(){Delete();}"

    Length (me) returns Integer is static ;
    ---C++: inline

    Upper (me) returns Integer is static;
    ---Purpose: Returns the upper bound
    ---C++: inline
              
    Lock (me) returns Address is static ;
    ---Purpose: Locks the array <me> in memory and 
    --          returns its virtual address
		

    Unlock (me) is static;
    ---Purpose: unlocks the array <me> from memory
		
    ShallowDump (me; S: in out OStream)
    --Purpose: Prints the contents at the first level of <me> on
    --         the stream <s>. The Root version of ShallowDump prints
    --         the name of the class <me> is an instance of, 
    --         followed by its memory address.
    ---C++:  function call
      is redefined;


fields
    mySize : Integer is protected;
    myData : DBVArray from DBC is protected;
end BaseArray;
