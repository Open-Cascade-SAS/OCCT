-- File:	IntParam.cdl
-- Created:	Mon Nov 30 16:57:11 1992
-- Author:	Christian CAILLET
--		<cky@sdsun1>
---Copyright:	 Matra Datavision 1992


class IntParam  from IFSelect  inherits TShared

    ---Purpose : This class simply allows to access an Integer value through a
    --           Handle, as a String can be (by using HString).
    --           Hence, this value can be accessed : read and modified, without
    --           passing through the specific object which detains it. Thus,
    --           parameters of a Selection or a Dispatch (according its type)
    --           can be controlled directly from the ShareOut which contains them
    --           
    --           Additionnaly, an IntParam can be bound to a Static.
    --           Remember that for a String, binding is immediate, because the
    --           string value of a Static is a HAsciiString, it then suffices
    --           to get its Handle.
    --           For an Integer, an IntParam can designate (by its name) a
    --           Static : each time its value is required or set, the Static
    --           is aknowledged

uses Integer, CString, AsciiString

is
 
    Create returns mutable IntParam;
    ---Purpose : Creates an IntParam. Initial value is set to zer

    SetStaticName (me : mutable; statname : CString);
    ---Purpose : Commands this IntParam to be bound to a Static
    --           Hence, Value will return the value if this Static if it is set
    --           Else, Value works on the locally stored value
    --           SetValue also will set the value of the Static
    --           This works only for a present static of type integer or enum
    --           Else, it is ignored
    --           
    --           If <statname> is empty, disconnects the IntParam from Static

    StaticName (me) returns CString;
    ---Purpose : Returns the name of static parameter to which this IntParam
    --           is bound, empty if none

    Value (me) returns Integer is static;
    ---Purpose : Reads Integer Value of the IntParam. If a StaticName is
    --           defined and the Static is set, looks in priority the value
    --           of the static

    SetValue (me : mutable; val : Integer) is static;
    ---Purpose : Sets a new Integer Value for the IntParam. If a StaticName is
    --           defined and the Static is set, also sets the value of the static

fields

    theval : Integer;
    thestn : AsciiString;

end IntParam;
