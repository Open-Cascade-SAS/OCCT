-- Created on: 2002-12-12
-- Created by: data exchange team
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class SurfaceSection from StepElement
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity SurfaceSection

uses
    MeasureOrUnspecifiedValue from StepElement

is
    Create returns SurfaceSection from StepElement;
	---Purpose: Empty constructor

    Init (me: mutable; aOffset: MeasureOrUnspecifiedValue from StepElement;
                       aNonStructuralMass: MeasureOrUnspecifiedValue from StepElement;
                       aNonStructuralMassOffset: MeasureOrUnspecifiedValue from StepElement);
	---Purpose: Initialize all fields (own and inherited)

    Offset (me) returns MeasureOrUnspecifiedValue from StepElement;
	---Purpose: Returns field Offset
    SetOffset (me: mutable; Offset: MeasureOrUnspecifiedValue from StepElement);
	---Purpose: Set field Offset

    NonStructuralMass (me) returns MeasureOrUnspecifiedValue from StepElement;
	---Purpose: Returns field NonStructuralMass
    SetNonStructuralMass (me: mutable; NonStructuralMass: MeasureOrUnspecifiedValue from StepElement);
	---Purpose: Set field NonStructuralMass

    NonStructuralMassOffset (me) returns MeasureOrUnspecifiedValue from StepElement;
	---Purpose: Returns field NonStructuralMassOffset
    SetNonStructuralMassOffset (me: mutable; NonStructuralMassOffset: MeasureOrUnspecifiedValue from StepElement);
	---Purpose: Set field NonStructuralMassOffset

fields
    theOffset: MeasureOrUnspecifiedValue from StepElement;
    theNonStructuralMass: MeasureOrUnspecifiedValue from StepElement;
    theNonStructuralMassOffset: MeasureOrUnspecifiedValue from StepElement;

end SurfaceSection;
