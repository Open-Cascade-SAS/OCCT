-- Created on: 1994-06-01
-- Created by: Christian CAILLET
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ComputeStatus  from IGESSelect  inherits ModelModifier from IGESSelect

    ---Purpose : Computes Status of IGES Entities for a whole IGESModel.
    --           This concerns SubordinateStatus and UseFlag, which must have
    --           some definite values according the way they are referenced.
    --           (see definitions of Logical use, Physical use, etc...)
    --           
    --           Works by calling a BasicEditor from IGESData. Works on the
    --           whole produced (target) model, because computation is global.

uses AsciiString from TCollection,
     IGESModel, CopyTool, ContextModif

is

    Create returns mutable ComputeStatus;
    ---Purpose : Creates an ComputeStatus, which uses the system Date


    Performing (me; ctx : in out ContextModif;
    	        target  : mutable IGESModel;
                TC      : in out CopyTool);
    ---Purpose : Specific action : it first evaluates the required values for
    --           Subordinate Status and Use Flag (in Directory Part of each
    --           IGES Entity). Then it corrects them, for the whole target.
    --           Works with a Protocol. Implementation uses BasicEditor

    Label (me) returns AsciiString from TCollection;
    ---Purpose : Returns a text which is
    --           "Compute Subordinate Status and Use Flag"

end ComputeStatus;
