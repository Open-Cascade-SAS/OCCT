-- File:        OrdinalDate.cdl
-- Created:     Mon Dec  4 12:02:28 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWOrdinalDate from RWStepBasic

	---Purpose : Read & Write Module for OrdinalDate

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     OrdinalDate from StepBasic

is

	Create returns RWOrdinalDate;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable OrdinalDate from StepBasic);

	WriteStep (me; SW : in out StepWriter; ent : OrdinalDate from StepBasic);

end RWOrdinalDate;
