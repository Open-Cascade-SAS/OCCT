-- Created on: 2008-09-01
-- Created by: Vladislav ROMASHKO
-- Copyright (c) 2008-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


private class SplitData from Voxel

    ---Purpose: A container of split information.
    --          An instance of this class is used as a slice 
    --          in inner representation of recursive octtree voxels.

is

    Create
    ---Purpose: An empty constructor.
    returns SplitData from Voxel;

    GetValues(me : in out)
    ---Purpose: Gives access to the values.
    ---C++: return &
    returns Address from Standard;

    GetSplitData(me : in out)
    ---Purpose: Gives access to the next split data.
    ---C++: return &
    returns Address from Standard;

fields

    myValues    : Address from Standard;
    mySplitData : Address from Standard;
    
end SplitData;

