-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MarkerSelect from StepVisual inherits SelectType from StepData

	-- <MarkerSelect> is an EXPRESS Select Type construct translation.
	-- it gathers : enum MarkerType

uses Transient, SelectMember from StepData, MarkerMember from StepVisual

is

	Create returns MarkerSelect;
	---Purpose : Returns a MarkerSelect SelectType

	CaseNum (me; ent : Transient) returns Integer;
	---Purpose: Recognizes a MarkerSelect Kind Entity that is :
	--        0 else

    NewMember (me) returns SelectMember from StepData  is redefined;
    ---Purpose : Returns a new MarkerMember

    CaseMem (me; sm : SelectMember from StepData) returns Integer is redefined;
    ---Purpose : Returns 1 for a SelectMember enum, named MARKER_TYPE

    MarkerMember (me) returns MarkerMember  from StepVisual;
    ---Purpose : Gives access to the MarkerMember in order to get/set its value

end MarkerSelect;
