-- Created on: 1998-08-17
-- Created by: Philippe MANGIN
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class ShapeLaw from BRepFill inherits  SectionLaw  from  BRepFill

	---Purpose: Build Section Law, with an Vertex, or an Wire
        ---Level: Advanced
       
uses 
 SectionLaw          from GeomFill,  
 HArray1OfSectionLaw from  GeomFill, 
 HArray1OfShape      from  TopTools,  
 Shape               from  GeomAbs,
 Vertex              from  TopoDS, 
 Wire                from  TopoDS,  
 Edge                from  TopoDS,  
 Shape               from  TopoDS, 
 Function            from  Law

is  
  Create (V:  Vertex  from  TopoDS;   
          Build  :  Boolean = Standard_True )  
    ---Purpose: Construct an constant Law  
  returns  ShapeLaw  from BRepFill;   

  Create (W:Wire  from  TopoDS;   
          Build :  Boolean = Standard_True)   
     ---Purpose: Construct an constant Law   
  returns ShapeLaw from BRepFill;  
   
  Create  (W:  Wire  from  TopoDS;  
           L:  Function  from  Law; 
           Build :  Boolean = Standard_True)   
    ---Purpose: Construct an evolutive Law         
  returns ShapeLaw from BRepFill;      

  IsVertex(me) 
    ---Purpose: Say if the input shape is a  vertex. 
  returns  Boolean   
  is  redefined; 
   
  IsConstant(me) 
    ---Purpose: Say if the Law is  Constant.        
  returns  Boolean   
  is  redefined;        

  ConcatenedLaw(me)  
   ---Purpose: Give the law build on a concaneted section         
  returns SectionLaw from GeomFill 
  is  redefined;    
  
  Continuity(me; Index  :  Integer; 
    	         TolAngular  :  Real)
  returns  Shape  from  GeomAbs  
  is  redefined;  
   
  VertexTol(me; Index  :  Integer;   
                Param  :  Real) 
  returns  Real   
  is  redefined;  
  
  Vertex(me;  Index  :  Integer; 
              Param  :  Real) 
  returns Vertex  from  TopoDS 
  is  redefined;	    
   
  D0(me:mutable;  Param  :  Real;   
     S  :  out  Shape  from  TopoDS)   
    is  redefined;  
   
  Edge(me; Index  :  Integer)  
   ---C++: return const &
   ---C++: inline
  returns  Edge  from  TopoDS;  
   
  Init(me  :  mutable;  B  :  Boolean)  is  private;
   
fields
  myShape:  Shape          from  TopoDS;
  myEdges:  HArray1OfShape from  TopTools;   
  TheLaw :  Function       from  Law;   
  vertex :  Boolean        from  Standard is  protected; 
end ShapeLaw;
