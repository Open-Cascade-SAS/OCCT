-- Created on: 1996-01-29
-- Created by: Robert COUBLANC
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class CompositionFilter from SelectMgr inherits Filter from SelectMgr
    	---Purpose: A framework to define a compound filter composed of
    	-- two or more simple filters.

uses
    Boolean      from Standard,
    ListOfFilter from SelectMgr,
    ShapeEnum from TopAbs
is

    Add(me : mutable; afilter : Filter from SelectMgr);
    	--- Purpose: Adds the filter afilter to a filter object created by a
    	-- filter class inheriting this framework.   
    Remove(me:mutable;aFilter : Filter from SelectMgr);

    	--- Purpose: Removes the filter aFilter from this framework.
    IsEmpty(me) returns Boolean;
    	---Purpose: Returns true if this framework is empty.
    IsIn(me;aFilter : Filter from SelectMgr)
    returns Boolean;

    	--- Purpose: Returns true if the filter aFilter is in this framework.
    
    StoredFilters(me) returns ListOfFilter from SelectMgr;
    	---C++: return const &
    	---C++: inline
    	---Purpose: Returns the list of stored filters from this framework.

    Clear(me:mutable);
    	---Purpose: Clears the filters used in this framework.
    ActsOn(me; aStandardMode : ShapeEnum from TopAbs)
    returns Boolean from Standard is redefined virtual;


fields

    myFilters : ListOfFilter from SelectMgr is protected;

end CompositionFilter;
