-- Created on: 1994-11-08
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class EdgeInterferenceTool from TopOpeBRepDS 

	---Purpose: a tool computing complex transition on Edge.

uses

    Orientation from TopAbs,
    CurveTransition from TopTrans,
    Interference from TopOpeBRepDS,
    Point from TopOpeBRepDS,
    Shape from TopoDS

is

    Create returns EdgeInterferenceTool from TopOpeBRepDS;
    
    Init(me : in out; 
         E : Shape from TopoDS; 
         I : Interference from TopOpeBRepDS)
    is static;
    
    Add(me : in out; 
        E : Shape from TopoDS;
        V : Shape from TopoDS;
        I : Interference from TopOpeBRepDS)
    is static;
    
    Add(me : in out; 
        E : Shape from TopoDS;
	P : Point from TopOpeBRepDS;
        I : Interference from TopOpeBRepDS)
    is static;
    
    Transition(me; I : Interference from TopOpeBRepDS)
    is static;
    
fields
    
    myEdgeOrientation : Orientation from TopAbs;
    myEdgeOriented    : Integer from Standard;
    myTool            : CurveTransition from TopTrans;

end EdgeInterferenceTool from TopOpeBRepDS;
