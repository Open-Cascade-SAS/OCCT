-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class AutoDesignPresentedItem from StepAP214 

    -- updated for CC1 Rev4 (usage of Select)

inherits PresentedItem from StepVisual

uses

	HArray1OfAutoDesignPresentedItemSelect from StepAP214, 
	AutoDesignPresentedItemSelect from StepAP214
is

	Create returns mutable AutoDesignPresentedItem;
	---Purpose: Returns a AutoDesignPresentedItem

	Init (me : mutable;
	      aItems : mutable HArray1OfAutoDesignPresentedItemSelect from StepAP214) is virtual;

	-- Specific Methods for Field Data Access --

	SetItems(me : mutable; aItems : mutable HArray1OfAutoDesignPresentedItemSelect);
	Items (me) returns mutable HArray1OfAutoDesignPresentedItemSelect;
	ItemsValue (me; num : Integer) returns AutoDesignPresentedItemSelect;
	NbItems (me) returns Integer;

fields

	items : HArray1OfAutoDesignPresentedItemSelect from StepAP214;

end AutoDesignPresentedItem;
