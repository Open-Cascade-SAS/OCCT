-- Created on: 1993-01-09
-- Created by: CKY / Contract Toubro-Larsen ( Anand NATRAJAN )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ExternalRefName from IGESBasic  inherits IGESEntity

        ---Purpose: defines ExternalRefName, Type <416> Form <3>
        --          in package IGESBasic
        --          Used when it is assumed that a copy of the subfigure
        --          exists in native form on the receiving system

uses

        HAsciiString from TCollection

is

        Create returns mutable ExternalRefName;

        -- Specific Methods pertaining to the class

        Init (me : mutable; anExtName : HAsciiString);
        ---Purpose : This method is used to set the fields of the class
        --           ExternalRefName
        --       - anExtName : External Reference Entity Symbolic Name

        ReferenceName (me) returns HAsciiString from TCollection;
        ---Purpose : returns External Reference Entity Symbolic Name

fields

--
-- Class    : IGESBasic_ExternalRefName
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class ExternalRefName.
--
-- Reminder : A ExternalRefName instance is defined by :
--            - External Reference Entity Symbolic Name

        theExtRefEntitySymbName : HAsciiString from TCollection;

end ExternalRefName;
