-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class OrganizationalAddress from StepBasic 

inherits Address from StepBasic 

uses

	HArray1OfOrganization from StepBasic, 
	HAsciiString from TCollection, 
	Organization from StepBasic
is

	Create returns mutable OrganizationalAddress;
	---Purpose: Returns a OrganizationalAddress


	Init (me : mutable;
	      hasAinternalLocation : Boolean from Standard;
	      aInternalLocation : mutable HAsciiString from TCollection;
	      hasAstreetNumber : Boolean from Standard;
	      aStreetNumber : mutable HAsciiString from TCollection;
	      hasAstreet : Boolean from Standard;
	      aStreet : mutable HAsciiString from TCollection;
	      hasApostalBox : Boolean from Standard;
	      aPostalBox : mutable HAsciiString from TCollection;
	      hasAtown : Boolean from Standard;
	      aTown : mutable HAsciiString from TCollection;
	      hasAregion : Boolean from Standard;
	      aRegion : mutable HAsciiString from TCollection;
	      hasApostalCode : Boolean from Standard;
	      aPostalCode : mutable HAsciiString from TCollection;
	      hasAcountry : Boolean from Standard;
	      aCountry : mutable HAsciiString from TCollection;
	      hasAfacsimileNumber : Boolean from Standard;
	      aFacsimileNumber : mutable HAsciiString from TCollection;
	      hasAtelephoneNumber : Boolean from Standard;
	      aTelephoneNumber : mutable HAsciiString from TCollection;
	      hasAelectronicMailAddress : Boolean from Standard;
	      aElectronicMailAddress : mutable HAsciiString from TCollection;
	      hasAtelexNumber : Boolean from Standard;
	      aTelexNumber : mutable HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      hasAinternalLocation : Boolean from Standard;
	      aInternalLocation : mutable HAsciiString from TCollection;
	      hasAstreetNumber : Boolean from Standard;
	      aStreetNumber : mutable HAsciiString from TCollection;
	      hasAstreet : Boolean from Standard;
	      aStreet : mutable HAsciiString from TCollection;
	      hasApostalBox : Boolean from Standard;
	      aPostalBox : mutable HAsciiString from TCollection;
	      hasAtown : Boolean from Standard;
	      aTown : mutable HAsciiString from TCollection;
	      hasAregion : Boolean from Standard;
	      aRegion : mutable HAsciiString from TCollection;
	      hasApostalCode : Boolean from Standard;
	      aPostalCode : mutable HAsciiString from TCollection;
	      hasAcountry : Boolean from Standard;
	      aCountry : mutable HAsciiString from TCollection;
	      hasAfacsimileNumber : Boolean from Standard;
	      aFacsimileNumber : mutable HAsciiString from TCollection;
	      hasAtelephoneNumber : Boolean from Standard;
	      aTelephoneNumber : mutable HAsciiString from TCollection;
	      hasAelectronicMailAddress : Boolean from Standard;
	      aElectronicMailAddress : mutable HAsciiString from TCollection;
	      hasAtelexNumber : Boolean from Standard;
	      aTelexNumber : mutable HAsciiString from TCollection;
	      aOrganizations : mutable HArray1OfOrganization from StepBasic;
	      aDescription : mutable HAsciiString from TCollection) is virtual;

	-- Specific Methods for Field Data Access --

	SetOrganizations(me : mutable; aOrganizations : mutable HArray1OfOrganization);
	Organizations (me) returns mutable HArray1OfOrganization;
	OrganizationsValue (me; num : Integer) returns mutable Organization;
	NbOrganizations (me) returns Integer;
	SetDescription(me : mutable; aDescription : mutable HAsciiString);
	Description (me) returns mutable HAsciiString;

fields

	organizations : HArray1OfOrganization from StepBasic;
	description : HAsciiString from TCollection;

end OrganizationalAddress;
