-- Created on: 1997-02-12
-- Created by: Alexander BRIVIN
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Rotation from Vrml 

	---Purpose:  defines a Rotation node of VRML specifying matrix and transform properties.
    	--  This  node  defines  a  3D  rotation  about  an  arbitrary  axis  through  the  origin. 
    	--  By  default  :  myRotation  =  (0 0 1 0)

uses
 
    SFRotation  from  Vrml

is
 
    Create returns   Rotation from Vrml;

    Create  (  aRotation  :  SFRotation  from  Vrml ) 
    	returns   Rotation from Vrml;
      
    SetRotation ( me : in out; aRotation : SFRotation  from  Vrml );
    Rotation ( me )  returns  SFRotation  from  Vrml;

    Print  ( me;  anOStream: in out OStream from Standard) returns OStream from Standard;
    ---C++:  return  & 

fields
 
    myRotation  :  SFRotation  from  Vrml; -- Rotation

end Rotation;
