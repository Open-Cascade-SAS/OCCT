-- File:	StepFEA_CurveElementEndOffset.cdl
-- Created:	Thu Dec 12 17:51:03 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class CurveElementEndOffset from StepFEA
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity CurveElementEndOffset

uses
    CurveElementEndCoordinateSystem from StepFEA,
    HArray1OfReal from TColStd

is
    Create returns CurveElementEndOffset from StepFEA;
	---Purpose: Empty constructor

    Init (me: mutable; aCoordinateSystem: CurveElementEndCoordinateSystem from StepFEA;
                       aOffsetVector: HArray1OfReal from TColStd);
	---Purpose: Initialize all fields (own and inherited)

    CoordinateSystem (me) returns CurveElementEndCoordinateSystem from StepFEA;
	---Purpose: Returns field CoordinateSystem
    SetCoordinateSystem (me: mutable; CoordinateSystem: CurveElementEndCoordinateSystem from StepFEA);
	---Purpose: Set field CoordinateSystem

    OffsetVector (me) returns HArray1OfReal from TColStd;
	---Purpose: Returns field OffsetVector
    SetOffsetVector (me: mutable; OffsetVector: HArray1OfReal from TColStd);
	---Purpose: Set field OffsetVector

fields
    theCoordinateSystem: CurveElementEndCoordinateSystem from StepFEA;
    theOffsetVector: HArray1OfReal from TColStd;

end CurveElementEndOffset;
