-- File:	IGESGeom_ToolBoundedSurface.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolBoundedSurface  from IGESGeom

    ---Purpose : Tool to work on a BoundedSurface. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses BoundedSurface from IGESGeom,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolBoundedSurface;
    ---Purpose : Returns a ToolBoundedSurface, ready to work


    ReadOwnParams (me; ent : mutable BoundedSurface;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : BoundedSurface;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : BoundedSurface;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a BoundedSurface <ent>, from
    --           its specific (own) parameters

    DirChecker (me; ent : BoundedSurface) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : BoundedSurface;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : BoundedSurface; entto : mutable BoundedSurface;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : BoundedSurface;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolBoundedSurface;
