-- File:	StepToTopoDS_TranslateCompositeCurve.cdl
-- Created:	Fri Feb 12 13:17:04 1999
-- Author:	Andrey BETENEV
--		<abv@doomox.nnov.matra-dtv.fr>
---Copyright:	 Matra Datavision 1999


class TranslateCompositeCurve from StepToTopoDS 
    inherits Root from StepToTopoDS
	---Purpose: Translate STEP entity composite_curve to TopoDS_Wire
	--          If surface is given, the curve is assumed to lie on that
        --          surface and in case if any segment of it is a
	--          curve_on_surface, the pcurve for that segment will be taken.
	--          Note: a segment of composite_curve may be itself 
        --                composite_curve. Only one-level protection against 
        --                cyclic references is implemented.

uses
    TransientProcess from Transfer,
    CompositeCurve   from StepGeom,
    Surface          from StepGeom,
    Surface          from Geom,
    Wire             from TopoDS
    
is

    Create returns TranslateCompositeCurve;
        ---Purpose: Empty constructor
	
    Create (CC: CompositeCurve from StepGeom;
    	    TP: TransientProcess from Transfer)
    	returns TranslateCompositeCurve;
        ---Purpose: Translates standalone composite_curve

    Create (CC: CompositeCurve from StepGeom;
    	    TP: TransientProcess from Transfer;
    	    S : Surface from StepGeom;
    	    Surf: Surface from Geom)
    	returns TranslateCompositeCurve;
        ---Purpose: Translates composite_curve lying on surface 
	
    Init (me: in out;
          CC: CompositeCurve from StepGeom;
    	  TP: TransientProcess from Transfer)
    	returns Boolean;
        ---Purpose: Translates standalone composite_curve

    Init (me: in out;
          CC: CompositeCurve from StepGeom;
    	  TP: TransientProcess from Transfer;
    	  S : Surface from StepGeom;
    	  Surf: Surface from Geom)
    	returns Boolean;
        ---Purpose: Translates composite_curve lying on surface 

    Value (me) returns Wire from TopoDS;
        ---Purpose: Returns result of last translation or null wire if failed.
	---C++: return const &

    IsInfiniteSegment (me) returns Boolean;
        ---Purpose: Returns True if composite_curve contains a segment with infinite parameters.
        ---C++: inline 

fields

    myWire: Wire from TopoDS;
    myInfiniteSegment: Boolean;

end TranslateCompositeCurve;
