-- Created on: 1993-06-23
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Curve from TopOpeBRepDS

    ---Purpose: A Geom curve and a tolerance.

uses

    Shape from TopoDS,
    Curve from Geom,
    Curve from Geom2d,
    Interference from TopOpeBRepDS

is

    Create returns Curve from TopOpeBRepDS; 

    Create(P : Curve from Geom; 
     	   T : Real from Standard; 
    	   IsWalk : Boolean from Standard = Standard_False)  
    returns Curve from TopOpeBRepDS; 
 
    DefineCurve(me : in out; 
           P : Curve from Geom; 
     	   T : Real from Standard; 
    	   IsWalk : Boolean from Standard);

    Tolerance(me : in out; tol : Real)
    ---Purpose: Update the tolerance
    is static;
	
    SetSCI(me : in out; I1,I2 : Interference from TopOpeBRepDS)
    ---Purpose: define the interferences face/curve.
    is static;

    GetSCI1(me) returns any Interference from TopOpeBRepDS
    ---C++: return const &
    is static;

    GetSCI2(me) returns any Interference from TopOpeBRepDS
    ---C++: return const &
    is static;

    GetSCI(me; I1,I2 : in out Interference from TopOpeBRepDS)
    is static;

    SetShapes(me : in out; S1,S2 : Shape from TopoDS)
    is static; 
    
    GetShapes(me; S1,S2 : in out Shape from TopoDS)
    is static;

    Shape1(me) returns Shape from TopoDS
    ---C++: return const &
    is static;
 
    ChangeShape1(me : in out) returns Shape from TopoDS
    ---C++: return &
    is static;
    Shape2(me) returns Shape from TopoDS
    ---C++: return const &
    is static;

    ChangeShape2(me : in out) returns Shape from TopoDS
    ---C++: return &
    is static;

    Curve(me) returns any Curve from Geom
    ---C++: return const &
    is static;

    SetRange(me : in out ; First, Last : Real from Standard)
    is static;
    
    Range(me; First, Last : out Real from Standard) 
    returns Boolean from Standard
    is static;

    Tolerance(me) returns Real from Standard
    is static;

    ChangeCurve(me : in out) returns any Curve from Geom
    ---C++: return &
    is static;
	
    Curve(me : in out; C3D : Curve from Geom; Tol : Real from Standard)
    is static;
    
    Curve1(me) returns any Curve from Geom2d
    ---C++: return const &
    is static;

    Curve1(me : in out; PC1 : Curve from Geom2d)
    is static;
    
    Curve2(me) returns any Curve from Geom2d
    ---C++: return const &
    is static;

    Curve2(me : in out; PC2 : Curve from Geom2d)
    is static;
    
    IsWalk(me) returns Boolean from Standard;
    ChangeIsWalk(me: in out; B : Boolean from Standard);

    Keep(me) returns Boolean from Standard
    is static;
    ChangeKeep(me : in out; B : Boolean from Standard)
    is static;

    Mother(me) returns Integer from Standard
    is static;
    ChangeMother(me : in out; I : Integer from Standard)
    is static;

    DSIndex(me) returns Integer from Standard
    is static;
    ChangeDSIndex(me : in out; I : Integer from Standard)
    is static;

    Dump(me; OS : in out OStream from Standard; 
    	     index : Integer from Standard;
             compact : Boolean = Standard_True)
    ---C++: return &
    returns OStream from Standard
    is static;
	  

fields

    myCurve         : Curve from Geom;
    myFirst,myLast  : Real from Standard;
    myRangeDefined  : Boolean from Standard;
    myTolerance     : Real from Standard;
    myIsWalk        : Boolean from Standard;
    
    myS1    : Shape from TopoDS;
    myS2    : Shape from TopoDS;
    mySCI1  : Interference from TopOpeBRepDS;
    mySCI2  : Interference from TopOpeBRepDS;

    myKeep          : Boolean from Standard;
    myMother        : Integer;
    myDSIndex       : Integer;
    
end Curve;
