-- Created on: 1992-12-15
-- Created by: Jean Louis FRENKEL
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



deferred class Root from Prs3d

    	---Purpose: A root class for the standard presentation algorithms
    	-- of the StdPrs package.
    	--          
uses
    Presentation from Prs3d,
    Structure from Graphic3d,
    Group from Graphic3d

is
    CurrentGroup(myclass; Prs3d: Presentation from Prs3d) returns Group from Graphic3d;
    	---Purpose: Returns the current group of primititves inside graphic
    	-- objects in the display.
    	-- A group also contains the attributes whose ranges are
    	-- limited to the primitives in it. 
    
    NewGroup (myclass; Prs3d: Presentation from Prs3d ) returns Group from Graphic3d ;
    	---Purpose: Returns the new group of primitives inside graphic
    	-- objects in the display.
    	-- A group also contains the attributes whose ranges are limited to the primitives in it.
    
end Root from Prs3d;
