-- Created on: 1993-01-09
-- Created by: CKY / Contract Toubro-Larsen ( SIVA )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SolidInstance from IGESSolid  inherits IGESEntity

        ---Purpose: defines SolidInstance, Type <430> Form Number <0>
        --          in package IGESSolid
        --          This provides a mechanism for replicating a solid
        --          representation.
        --          
        --          From IGES-5.3, Form may be <1> for a BREP
        --          Else it is for a Boolean Tree, Primitive, other Solid Inst.

uses  Integer  -- no one specific type


is

        Create returns mutable SolidInstance;

        -- Specific Methods pertaining to the class

        Init (me       : mutable; 
              anEntity : IGESEntity);
        ---Purpose : This method is used to set the fields of the class
        --           SolidInstance
        --       - anEntity : the entity corresponding to the solid

    	IsBrep (me) returns Boolean;
	---Purpose : Tells if a SolidInstance is for a BREP
	--           Default is False

    	SetBrep (me : mutable; brep : Boolean);
	---Purpose : Sets or unsets the Brep status (FormNumber = 1 else 0)

        Entity(me) returns IGESEntity;
        ---Purpose : returns the solid entity

fields

--
-- Class    : IGESSolid_SolidInstance
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class SolidInstance.
--
-- Reminder : A SolidInstance instance is defined by :
--            a pointer to a solid entity
--

        theEntity : IGESEntity;
            -- the solid entity

end SolidInstance;
