-- Created on: 1994-06-16
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class FileDescription from HeaderSection 

inherits TShared from MMgt

uses

	HArray1OfHAsciiString from Interface,
	HAsciiString from TCollection
is

	Create returns mutable FileDescription;
	---Purpose: Returns a FileDescription

	Init (me : mutable;
	      aDescription : mutable HArray1OfHAsciiString from Interface;
	      aImplementationLevel : mutable HAsciiString from TCollection);

	-- Specific Methods for Field Data Access --

	SetDescription(me : mutable; aDescription : mutable HArray1OfHAsciiString);
	Description (me) returns mutable HArray1OfHAsciiString;
	DescriptionValue (me; num : Integer) returns mutable HAsciiString;
	NbDescription (me) returns Integer;
	SetImplementationLevel(me : mutable; aImplementationLevel : mutable HAsciiString);
	ImplementationLevel (me) returns mutable HAsciiString;

fields

	description : HArray1OfHAsciiString from Interface;
	implementationLevel : HAsciiString from TCollection;

end FileDescription;
