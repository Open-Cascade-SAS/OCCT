-- Created on: 1999-07-08
-- Created by: Sergey RUIN
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class AISPresentation_1 from PPrsStd 
    inherits Attribute from PDF

	---Purpose: 
    
uses    HExtendedString from PCollection
is

    Create returns mutable AISPresentation_1 from PPrsStd;
	
    IsDisplayed(me) returns Boolean from Standard;
    SetDisplayed(me : mutable; B : Boolean from Standard);

    SetDriverGUID(me: mutable; guid: HExtendedString from PCollection );     
    GetDriverGUID(me) returns HExtendedString from PCollection; 
    
    Color(me) returns Integer from Standard;
    SetColor(me : mutable; C : Integer from Standard);
    
    Transparency(me) returns Real from Standard;
    SetTransparency(me : mutable; T : Real from Standard);    
    
    Material(me) returns Integer from Standard;
    SetMaterial(me : mutable; M : Integer from Standard);    
   
    Width(me) returns Real from Standard;
    SetWidth(me : mutable; W : Real from Standard);
 
    Mode(me)    returns Integer from Standard; 
    SetMode(me : mutable; M : Integer from Standard);    
fields

    myIsDisplayed         : Boolean              from Standard;
    myDriverGUID          : HExtendedString      from PCollection; 
    myTransparency        : Real                 from Standard;
    myColor               : Integer              from Standard;
    myMaterial            : Integer              from Standard;
    myWidth               : Real                 from Standard; 
    myMode                : Integer              from Standard;
end AISPresentation_1;
