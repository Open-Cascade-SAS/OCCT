-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ConversionBasedUnitAndPlaneAngleUnit from StepBasic inherits ConversionBasedUnit from StepBasic 

	--- This classe is an implementation of EXPRESS
	--  ANDOR Subtype Declaration.
uses

    PlaneAngleUnit from StepBasic, 
    DimensionalExponents from StepBasic, 
    HAsciiString from TCollection, 
    MeasureWithUnit from StepBasic
    
is

    Create returns mutable ConversionBasedUnitAndPlaneAngleUnit;
	---Purpose: Returns a ConversionBasedUnitAndPlaneAngleUnit

    Init (me: mutable; aDimensions: mutable DimensionalExponents from StepBasic)
    is redefined;

    Init (me: mutable; aDimensions: mutable DimensionalExponents from StepBasic;
		       aName      : mutable HAsciiString from TCollection;
		       aConversionFactor: mutable MeasureWithUnit from StepBasic) is redefined;

    -- Specific Methods for Field Data Access --

    SetPlaneAngleUnit(me: mutable; aPlaneAngleUnit: mutable PlaneAngleUnit);
    
    PlaneAngleUnit (me) returns mutable PlaneAngleUnit;

fields

    planeAngleUnit: PlaneAngleUnit from StepBasic;

end ConversionBasedUnitAndPlaneAngleUnit;
