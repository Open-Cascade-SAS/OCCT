-- File:        FacetedBrep.cdl
-- Created:     Mon Dec  4 12:02:26 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWFacetedBrep from RWStepShape

	---Purpose : Read & Write Module for FacetedBrep

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     FacetedBrep from StepShape,
     EntityIterator from Interface

is

	Create returns RWFacetedBrep;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable FacetedBrep from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : FacetedBrep from StepShape);

	Share(me; ent : FacetedBrep from StepShape; iter : in out EntityIterator);

end RWFacetedBrep;
