-- File:	IGESDimen_ToolDimensionUnits.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolDimensionUnits  from IGESDimen

    ---Purpose : Tool to work on a DimensionUnits. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses DimensionUnits from IGESDimen,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolDimensionUnits;
    ---Purpose : Returns a ToolDimensionUnits, ready to work


    ReadOwnParams (me; ent : mutable DimensionUnits;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : DimensionUnits;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : DimensionUnits;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a DimensionUnits <ent>, from
    --           its specific (own) parameters

    OwnCorrect (me; ent : mutable DimensionUnits) returns Boolean  is static;
    ---Purpose : Sets automatic unambiguous Correction on a DimensionUnits
    --           (NbPropertyValues forced to 6)

    DirChecker (me; ent : DimensionUnits) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : DimensionUnits;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : DimensionUnits; entto : mutable DimensionUnits;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : DimensionUnits;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolDimensionUnits;
