-- Created on: 2000-02-07
-- Created by: data exchange team
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class AlgoContainer from IGESToBRep inherits TShared from MMgt

    ---Purpose: 

uses

    ToolContainer from IGESToBRep
    
is

    Create returns mutable AlgoContainer from IGESToBRep;
    	---Purpose: Empty constructor
	
    SetToolContainer (me: mutable; TC: ToolContainer from IGESToBRep);
    	---C++    : inline
    	---Purpose: Sets ToolContainer
	
    ToolContainer (me) returns ToolContainer from IGESToBRep;
    	---C++    : inline
    	---Purpose: Returns ToolContainer
	
	
fields

    myTC     : ToolContainer from IGESToBRep;
    
end AlgoContainer;
