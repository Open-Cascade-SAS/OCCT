-- File:        CylindricalSurface.cdl
-- Created:     Mon Dec  4 12:02:25 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWCylindricalSurface from RWStepGeom

	---Purpose : Read & Write Module for CylindricalSurface

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     CylindricalSurface from StepGeom,
     EntityIterator from Interface

is

	Create returns RWCylindricalSurface;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable CylindricalSurface from StepGeom);

	WriteStep (me; SW : in out StepWriter; ent : CylindricalSurface from StepGeom);

	Share(me; ent : CylindricalSurface from StepGeom; iter : in out EntityIterator);

end RWCylindricalSurface;
