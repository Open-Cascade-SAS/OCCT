--
-- File      :  OrdinateDimension.cdl
-- Created   :  Mon 11 Jan 1993
-- Author    : CKY / Contract Toubro-Larsen ( SIVA )
--
---Copyright : MATRA-DATAVISION  1993
--

class OrdinateDimension from IGESDimen  inherits IGESEntity

        ---Purpose: defines IGES Ordinate Dimension, Type <218> Form <0, 1>,
        --          in package IGESDimen
        -- Note   : The ordinate dimension entity is used to
        --          indicate dimensions from a common base line.
        --          Dimensioning is only permitted along the XT
        --          or YT axis.

uses

        LeaderArrow from IGESDimen,
        WitnessLine from IGESDimen,
        GeneralNote from IGESDimen

is

        Create returns mutable OrdinateDimension;

            -- --specific-- --

        Init(me       : mutable;
             aNote    : GeneralNote;
             aType    : Boolean;
             aLine    : WitnessLine;
             anArrow  : LeaderArrow);
        -- This method is used to set fields of the
        -- class OrdinateDimension
        --       - aNote    : Note for the dimension
        --       - aType    : Type (Witness line or leader arrow)
        --                    (Ignored if form no. = 1)
        --       - aLine    : Witness line used for the dimension
        --       - anArrow  : Leader arrow used for the dimension

        IsLine(me) returns Boolean;
        ---Purpose : returns True if Witness Line and False if Leader (only for Form 0)

        IsLeader(me) returns Boolean;
        ---Purpose : returns True if Leader and False if Witness Line (only for Form 0)

        Note(me) returns GeneralNote;
        ---Purpose : returns the General Note entity associated.

        WitnessLine(me) returns WitnessLine;
        ---Purpose : returns the Witness Line associated or Null handle

        Leader(me) returns LeaderArrow;
        ---Purpose : returns the Leader associated or Null handle

fields

--
-- Class    : IGESDimen_OrdinateDimension
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class OrdinateDimension.
--
-- Reminder : A OrdinateDimension instance is defined by :
--            - A General Note
--            - A Boolean field determining whether a Witness Line
--                                or Leader is present
--            - A Witness Line
--            - A Leader Arrow
--

        theNote        : GeneralNote;
        isItLine       : Boolean;     --True if Witness Line, False if Leader
        theWitnessLine : WitnessLine;
        theLeader      : LeaderArrow;

end OrdinateDimension;
