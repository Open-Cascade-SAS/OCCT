-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PresentationLayerAssignment from StepVisual 

inherits TShared from MMgt

uses

	HAsciiString from TCollection, 
	HArray1OfLayeredItem from StepVisual, 
	LayeredItem from StepVisual
is

	Create returns PresentationLayerAssignment;
	---Purpose: Returns a PresentationLayerAssignment

	Init (me : mutable;
	      aName : HAsciiString from TCollection;
	      aDescription : HAsciiString from TCollection;
	      aAssignedItems : HArray1OfLayeredItem from StepVisual) is virtual;

	-- Specific Methods for Field Data Access --

	SetName(me : mutable; aName : HAsciiString);
	Name (me) returns HAsciiString;
	SetDescription(me : mutable; aDescription : HAsciiString);
	Description (me) returns HAsciiString;
	SetAssignedItems(me : mutable; aAssignedItems : HArray1OfLayeredItem);
	AssignedItems (me) returns HArray1OfLayeredItem;
	AssignedItemsValue (me; num : Integer) returns LayeredItem;
	NbAssignedItems (me) returns Integer;

fields

	name : HAsciiString from TCollection;
	description : HAsciiString from TCollection;
	assignedItems : HArray1OfLayeredItem from StepVisual; -- a SelectType

end PresentationLayerAssignment;
