-- File:	Blend_CSWalking.cdl
-- Created:	Thu Dec  2 11:33:03 1993
-- Author:	Jacques GOUSSARD
--		<jag@topsn2>
---Copyright:	 Matra Datavision 1993



generic class CSWalking from Blend 
    (TheVertex        as any;
     TheArc           as any;
     TheSurface       as any;
     TheCurve         as any;
     TheVertexTool    as any;
     TheArcTool       as any;
     TheSurfaceTool   as any;
     TheCurveTool     as any;
     TheTopolTool     as Transient;
     TheBlendTool     as any;
     ThePointOnRst    as any; -- as PointOnRst from Blend(TheArc)
     TheSeqPointOnRst as any; -- as Iterator from Blend(ThePointOnRst)
     TheExtremity     as any; -- as Extremity from Blend(TheVertex,TheArc,
                              --    ThePointOnRst,TheSeqPointOnRst)
     TheLine          as Transient) -- as Line from Blend(TheVertex,TheArc,
                                    --   ThePointOnRst,TheSeqPointOnRst,
                                    --   TheExtremity)
 


	---Purpose: 

uses Point            from Blend,
     Status           from Blend,
     Vector           from math,
     Matrix           from math,
     Pnt              from gp,
     Pnt2d            from gp,
     Vec              from gp,
     Vec2d            from gp,
     HArray1OfReal    from TColStd,
     Transition       from IntSurf,
     CSFunction       from Blend
--     CSFuncInv          from Blend
     

raises NotDone from StdFail


is

    Create(Curv : TheCurve; Surf: TheSurface; Domain: TheTopolTool)
    
    	returns CSWalking from Blend;


    Perform(me: in out; F       : in out CSFunction from Blend;
--                        FInv    : in out CSFuncInv  from Blend;
                        Pdep    : Real from Standard;
                        Pmax    : Real from Standard;
			MaxStep : Real from Standard;
			TolGuide: Real from Standard;
                        Soldep  : Vector from math;
                        Tolesp  : Real from Standard;
                        Fleche  : Real from Standard;
                        Appro   : Boolean from Standard = Standard_False)

    
    	is static;


    Complete(me: in out;F       : in out CSFunction from Blend;
--                        FInv    : in out FuncInv  from Blend;
                        Pmin    : Real from Standard)
			
	returns Boolean from Standard
	raises NotDone from StdFail
	is static;


    InternalPerform (me: in out;F       : in out CSFunction from Blend;
--                                FInv    : in out CSFuncInv  from Blend;
                                Sol     : in out Vector from math;
                                Bound   : Real from Standard)
			
	is static private;


    IsDone(me)
    
    	returns Boolean from Standard
	---C++: inline

	is static;




    Line(me)
    
    	returns TheLine
	---C++: inline
	---C++: return const&
	
    	raises NotDone from StdFail

	is static;





--    Recadre(me: in out; FInv : in out CSFuncInv from Blend;
--                        Sol: Vector from math;
--			Solrst : out Vector from math;
--			Indexsol: out Integer from Standard;
--   	    	    	IsVtx: out Boolean from Standard;
--                        Vtx: out TheVertex)
			
--        returns Boolean from Standard
--	is static private;


    Transition(me:in out; A: TheArc; Param: Real from Standard;
			  TLine,TArc: out Transition from IntSurf)

    	is static private;


    MakeExtremity(me:in out; Extrem : in out TheExtremity;
                             Index  : Integer from Standard;
    	                     Param  : Real from Standard;
			     IsVtx  : Boolean from Standard;
			     Vtx    : TheVertex)

    	is static private;


    CheckDeflectionOnSurf(me: in out; Psurf   : Pnt from gp;
                                      Ponsurf : Pnt2d from gp;
    	                              Tgsurf  : Vec from gp;
			              Tgonsurf: Vec2d from gp)
					
					
	returns Status from Blend
	is static private;


    CheckDeflectionOnCurv(me: in out; Pcurv   : Pnt from gp;
                                      Poncurv : Real from Standard;
    	                              Tgcurv  : Vec from gp)
					
					
	returns Status from Blend
	is static private;


    TestArret(me: in out; F    : in out CSFunction from Blend;
    	                  Sol  : Vector from math;
                          TestDeflection : Boolean from Standard;
                          State: Status from Blend)
    
    	returns Status from Blend
	is static private;



fields

    done         : Boolean          from Standard;
    line         : TheLine;
    surf         : TheSurface;
    curv         : TheCurve;
    domain       : TheTopolTool;

    tolesp       : Real             from Standard;
    tolgui       : Real             from Standard;
    pasmax       : Real             from Standard;
    fleche       : Real             from Standard;
    param        : Real             from Standard;
    firstparam   : Real             from Standard;
    firstsol     : HArray1OfReal    from TColStd;
    previousP    : Point            from Blend;
    rebrou       : Boolean          from Standard;
    iscomplete   : Boolean          from Standard;
    comptra      : Boolean          from Standard;
    sens         : Real             from Standard;

end CSWalking;
