-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class GP from XmlObjMgt

        ---Purpose: Translation of gp (simple geometry) objects
uses
    Trsf        from gp,
    Mat         from gp,
    XYZ         from gp,
    DOMString   from XmlObjMgt
is

    -- ---------------
    -- Package Methods
    -- ---------------

    -- from gp to string

    Translate (myclass; aTrsf : Trsf from gp)
    returns DOMString from XmlObjMgt;
        ---Level: Advanced 
    
    Translate (myclass; aMat : Mat from gp)
    returns DOMString from XmlObjMgt;
        ---Level: Advanced 
    
    Translate (myclass; anXYZ : XYZ from gp)
    returns DOMString from XmlObjMgt;
        ---Level: Advanced 
    
    -- from string to gp

    Translate (myclass; aStr : DOMString from XmlObjMgt; T : out Trsf from gp)
        returns Boolean from Standard;
        ---Level: Advanced 
    
    Translate (myclass; aStr : DOMString from XmlObjMgt; T : out Mat from gp)
        returns Boolean from Standard;
        ---Level: Advanced 
    
    Translate (myclass; aStr : DOMString from XmlObjMgt; T : out XYZ from gp)
        returns Boolean from Standard;
        ---Level: Advanced 
    
end;
