-- File:        GeometricRepresentationContextAndGlobalUnitAssignedContext.cdl
-- Created:     Thu Dec  7 14:30:30 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWGeometricRepresentationContextAndGlobalUnitAssignedContext from RWStepGeom

	---Purpose : Read & Write Module for GeometricRepresentationContextAndGlobalUnitAssignedContext

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     GeometricRepresentationContextAndGlobalUnitAssignedContext from StepGeom,
     EntityIterator from Interface

is

	Create returns RWGeometricRepresentationContextAndGlobalUnitAssignedContext;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable GeometricRepresentationContextAndGlobalUnitAssignedContext from StepGeom);

	WriteStep (me; SW : in out StepWriter; ent : GeometricRepresentationContextAndGlobalUnitAssignedContext from StepGeom);

	Share(me; ent : GeometricRepresentationContextAndGlobalUnitAssignedContext from StepGeom; iter : in out EntityIterator);

end RWGeometricRepresentationContextAndGlobalUnitAssignedContext;
