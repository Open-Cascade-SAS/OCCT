-- Created on: 1991-02-20
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class IntPoint from IntAna2d inherits Storable from Standard

    ---Purpose: Geometrical intersection between two 2d elements.


uses Pnt2d from gp

raises DomainError from Standard

is

    Create(X,Y: Real; U1,U2: Real)
    
    	---Purpose: Create an intersection point between 2 parametric 2d lines.
    	--          X,Y are the coordinate of the point. U1 is the parameter
    	--          on the first element, U2 the parameter on the second one.
    
    	returns IntPoint;


    Create(X,Y: Real; U1: Real)
    
    	---Purpose: Create an intersection point between a parametric 2d line,
    	--          and a line given by an implicit equation (ImplicitCurve).
    	--          X,Y are the coordinate of the point. U1 is the parameter
    	--          on the parametric element.
    
    	returns IntPoint;


    Create

	---Purpose: Empty constructor. It's necessary to use one of
	--          the SetValue method after this one.

    	returns IntPoint;


    SetValue(me : in out; X,Y: Real; U1,U2: Real)
    
	---Purpose: Set the values for a "non-implicit" point.
    is virtual;


    SetValue(me : in out; X,Y:Real; U1: Real)
    
	---Purpose: Set the values for an "implicit" point.
    is virtual;

    Value(me)
    
	---Purpose: Returns the geometric point.
    	---C++: inline
    	---C++: return const&
    	returns Pnt2d from gp

    is static;
    
    
    SecondIsImplicit(me)
    
    	---Purpose: Returns True if the second curve is implicit.
    	---C++: inline
    	returns Boolean from Standard
	
   is static;
	
    
    ParamOnFirst(me)
    
    	---Purpose: Returns the parameter on the first element.
    	---C++: inline
    	returns Real
	
    is static;

 
    ParamOnSecond(me)
    
    	---Purpose: Returns the parameter on the second element.
    	--          If the second element is an implicit curve, an exception
    	--          is raised.
    	---C++: inline
    	returns Real
	
	raises DomainError from Standard
    
    is static;



fields

    myu1        : Real  from Standard;
    myu2        : Real  from Standard;
    myp         : Pnt2d from gp;
    myimplicit  : Boolean from Standard;

end IntPoint;
