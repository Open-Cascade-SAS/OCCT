-- Created by: Peter KURNEV
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Objects from BOPTest 

 ---Purpose: 

uses  
    ListOfShape from BOPCol, 
    PDS from BOPDS,
    PaveFiller from BOPAlgo,
    Builder from BOPAlgo, 
    PBuilder from BOPAlgo, 
    BOP from BOPAlgo, 
    Section from BOPAlgo  
 
--raises

is 
    PaveFiller(myclass) 
     returns PaveFiller from BOPAlgo;  
    ---C++: return &   

    Init(myclass); 

    Clear(myclass); 

    PDS(myclass) 
     returns PDS from BOPDS; 
  
    Builder(myclass) 
     returns Builder from BOPAlgo; 
    ---C++: return & 
    
    BOP(myclass) 
     returns BOP from BOPAlgo; 
    ---C++: return & 
 
    Section(myclass) 
     returns Section from BOPAlgo;  
    ---C++: return &  
 
    Shapes(myclass)   
     returns ListOfShape from BOPCol; 
    ---C++: return &  
     
    Tools(myclass)   
     returns ListOfShape from BOPCol; 
    ---C++: return &  
    -- 
    SetBuilder(myclass; 
         theBuilder:PBuilder from BOPAlgo); 
  
    SetBuilderDefault(myclass); 
 
    SetRunParallel(myclass; 
            theFlag: Boolean from Standard); 
       
    RunParallel(myclass) 
        returns  Boolean from Standard; 
      
    SetFuzzyValue(myclass; 
            theValue: Real from Standard); 
       
    FuzzyValue(myclass) 
        returns  Real from Standard;     
 
--fields

end Objects;
