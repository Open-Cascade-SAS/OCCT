-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Hypr2d   from gp   inherits Storable

        ---Purpose:
        -- Describes a branch of a hyperbola in the plane (2D space).
        -- A hyperbola is defined by its major and minor radii, and
        -- positioned in the plane with a coordinate system (a
        -- gp_Ax22d object) of which:
        -- -   the origin is the center of the hyperbola,
        -- -   the "X Direction" defines the major axis of the hyperbola, and
        -- -   the "Y Direction" defines the minor axis of the hyperbola.
        --   This coordinate system is the "local coordinate system"
        -- of the hyperbola. The orientation of this coordinate
        -- system (direct or indirect) gives an implicit orientation to
        -- the hyperbola. In this coordinate system, the equation of
        -- the hyperbola is:
        -- X*X/(MajorRadius**2)-Y*Y/(MinorRadius**2) = 1.0
        -- The branch of the hyperbola described is the one located
        -- on the positive side of the major axis.
        -- The following schema shows the plane of the hyperbola,
        -- and in it, the respective positions of the three branches of
        -- hyperbolas constructed with the functions OtherBranch,
        -- ConjugateBranch1, and ConjugateBranch2:     
        --                         ^YAxis                
        --                         |                   
        --                  FirstConjugateBranch     
        --                         |        
        --        Other            |                Main
        --   --------------------- C ------------------------------>XAxis
        --        Branch           |                Branch
        --                         |
        --                         |         
        --                   SecondConjugateBranch
        --                         |         
        --
        -- Warning
        -- The major radius can be less than the minor radius.
        -- See Also
        -- gce_MakeHypr2d which provides functions for more
        -- complex hyperbola constructions
        -- Geom2d_Hyperbola which provides additional functions
        -- for constructing hyperbolas and works, in particular, with
        -- the parametric equations of hyperbolas

uses Ax2d   from gp,
     Ax22d  from gp, 
     Pnt2d  from gp,
     Trsf2d from gp,
     Vec2d  from gp

raises ConstructionError from Standard,
       DomainError       from Standard

is

  Create   returns Hypr2d;
        ---C++: inline
        --- Purpose : Creates of an indefinite hyperbola.


  Create (MajorAxis : Ax2d; 
    	  MajorRadius, MinorRadius : Real;
    	  Sense : Boolean from Standard = Standard_True)
     returns Hypr2d
        --- Purpose :
	--  Creates a hyperbola with radii MajorRadius and
        --   MinorRadius, centered on the origin of MajorAxis
        --   and where the unit vector of MajorAxis is the "X
        --   Direction" of the local coordinate system of the
        --   hyperbola. This coordinate system is direct if Sense
        --   is true (the default value), and indirect if Sense is false.
        --  Warnings :
        --  It is yet  possible to create an Hyperbola with 
        --  MajorRadius <= MinorRadius. 
        -- Raises ConstructionError if MajorRadius < 0.0 or MinorRadius < 0.0
     raises ConstructionError;

  Create (A : Ax22d; MajorRadius, MinorRadius : Real)
     returns Hypr2d
        ---C++: inline
        --- Purpose :
	--  a hyperbola with radii MajorRadius and
        --   MinorRadius, positioned in the plane by coordinate system A where:
        --   -   the origin of A is the center of the hyperbola,
        --   -   the "X Direction" of A defines the major axis of
        --    the hyperbola, that is, the major radius
        --    MajorRadius is measured along this axis, and
        --   -   the "Y Direction" of A defines the minor axis of
        --    the hyperbola, that is, the minor radius
        --    MinorRadius is measured along this axis, and
        --   -   the orientation (direct or indirect sense) of A
        --    gives the implicit orientation of the hyperbola.
        --  Warnings :
        --  It is yet  possible to create an Hyperbola with 
        --  MajorRadius <= MinorRadius.  
        -- Raises ConstructionError if MajorRadius < 0.0 or MinorRadius < 0.0
     raises ConstructionError;
	

  SetLocation (me : in out; P : Pnt2d)   is static;
        ---C++: inline
        --- Purpose : Modifies this hyperbola, by redefining its local
        -- coordinate system so that its origin becomes P.


  SetMajorRadius (me : in out; MajorRadius : Real)
     raises ConstructionError
        ---C++: inline
        ---Purpose: Modifies the major or minor radius of this hyperbola.
        -- Exceptions
        -- Standard_ConstructionError if MajorRadius or
        -- MinorRadius is negative.
     is static;


  SetMinorRadius (me : in out; MinorRadius : Real)
     raises ConstructionError
        ---C++: inline
        ---Purpose: Modifies the major or minor radius of this hyperbola.
        -- Exceptions
        -- Standard_ConstructionError if MajorRadius or
        -- MinorRadius is negative.
     is static;


  SetAxis (me : in out; A : Ax22d)   is static;
        ---C++: inline
        --- Purpose : Modifies this hyperbola, by redefining its local
        -- coordinate system so that it becomes A.


  SetXAxis (me : in out; A : Ax2d)   is static;
        ---C++: inline
        --- Purpose :
        --  Changes the major axis of the hyperbola. The minor axis is
        --  recomputed and the location of the hyperbola too.


  SetYAxis (me : in out; A : Ax2d) is static;
        ---C++: inline
        --- Purpose :
        --  Changes the minor axis of the hyperbola.The minor axis is
        --  recomputed and the location of the hyperbola too.


  Asymptote1 (me)   returns Ax2d
        ---C++: inline
	--- Purpose :
	--  In the local coordinate system of the hyperbola the equation of
	--  the hyperbola is (X*X)/(A*A) - (Y*Y)/(B*B) = 1.0 and the
        --  equation of the first asymptote is Y = (B/A)*X
        --  where A is the major radius of the hyperbola and B the minor
        --  radius of the hyperbola. 
        -- Raises ConstructionError if MajorRadius = 0.0
     raises ConstructionError
     is static;


  Asymptote2 (me)  returns Ax2d
        ---C++: inline
	--- Purpose :
	--  In the local coordinate system of the hyperbola the equation of
	--  the hyperbola is (X*X)/(A*A) - (Y*Y)/(B*B) = 1.0 and the
        --  equation of the first asymptote is Y = -(B/A)*X
        --  where A is the major radius of the hyperbola and B the minor
        --  radius of the hyperbola. 
        -- Raises ConstructionError if MajorRadius = 0.0
     raises ConstructionError
     is static;


  Coefficients (me; A, B, C, D, E, F : out Real)   is static;
        --- Purpose :
        --  Computes the coefficients of the implicit equation of 
        --  the hyperbola :
        --  A * (X**2) + B * (Y**2) + 2*C*(X*Y) + 2*D*X + 2*E*Y + F = 0.


  ConjugateBranch1 (me)  returns Hypr2d   is static;
        ---C++: inline
	--- Purpose :
	--  Computes the branch of hyperbola which is on the positive side of the 
	--  "YAxis" of <me>.


  ConjugateBranch2 (me)   returns Hypr2d  is static;
        ---C++: inline
	--- Purpose :
	-- Computes the branch of hyperbola which is on the negative side of the 
	--  "YAxis" of <me>.


  Directrix1 (me)   returns Ax2d   is static;
        ---C++: inline
        --- Purpose :
        --  Computes the directrix which is the line normal to the XAxis of the hyperbola
        --  in the local plane (Z = 0) at a distance d = MajorRadius / e 
        --  from the center of the hyperbola, where e is the eccentricity of
        --  the hyperbola.
        --  This line is parallel to the "YAxis". The intersection point
        --  between the "Directrix1" and the "XAxis" is the "Location" point
        --  of the "Directrix1".
        --  This point is on the positive side of the "XAxis".


  Directrix2 (me)  returns Ax2d is static;
        ---C++: inline
        --- Purpose :
        --  This line is obtained by the symmetrical transformation 
        --  of "Directrix1" with respect to the "YAxis" of the hyperbola.


  Eccentricity (me)  returns Real
        ---C++: inline
	--- Purpose :
	--  Returns the excentricity of the hyperbola (e > 1).
	--  If f is the distance between the location of the hyperbola
	--  and the Focus1 then the eccentricity e = f / MajorRadius. Raises DomainError if MajorRadius = 0.0.
     raises DomainError
     is static;


  Focal (me)   returns Real  is static;
        ---C++: inline
	--- Purpose :
	--  Computes the focal distance. It is the distance between the
        --  "Location" of the hyperbola and "Focus1" or "Focus2".


  Focus1 (me)    returns Pnt2d  is static;
        ---C++: inline
	--- Purpose :
	--  Returns the first focus of the hyperbola. This focus is on the
        --  positive side of the "XAxis" of the hyperbola.


  Focus2 (me)  returns Pnt2d  is static;
        ---C++: inline
        --- Purpose :
	--  Returns the second focus of the hyperbola. This focus is on the
        --  negative side of the "XAxis" of the hyperbola.


  Location (me)   returns Pnt2d  is static;
        ---C++: inline
        --- Purpose : 
        --  Returns  the location point of the hyperbola.
        --  It is the intersection point between the "XAxis" and 
        --  the "YAxis".
        ---C++: return const&


  MajorRadius (me)   returns Real  is static;
        ---C++: inline
	--- Purpose :
	--  Returns the major radius of the hyperbola (it is the radius
	--  corresponding to the "XAxis" of the hyperbola).


  MinorRadius (me)   returns Real  is static;
        ---C++: inline
	--- Purpose :
	--  Returns the minor radius of the hyperbola (it is the radius
	--  corresponding to the "YAxis" of the hyperbola).


  OtherBranch (me)   returns Hypr2d   is static;
        ---C++: inline
        --- Purpose :
	--  Returns the branch of hyperbola obtained by doing the 
	--  symmetrical transformation of <me> with respect to the 
	--  "YAxis" of <me>.


  Parameter (me)   returns Real
        ---C++: inline
        --- Purpose :
        --  Returns p = (e * e - 1) * MajorRadius where e is the 
        --  eccentricity of the hyperbola.
        -- Raises DomainError if MajorRadius = 0.0
     raises DomainError
     is static;


  Axis (me)   returns Ax22d   is static;
	--- Purpose : Returns the axisplacement of the hyperbola.
        ---C++: inline
        ---C++: return const&
  


  XAxis (me)   returns Ax2d   is static;
	--- Purpose : Computes an axis whose
        -- -   the origin is the center of this hyperbola, and
        -- -   the unit vector is the "X Direction" or "Y Direction"
        -- respectively of the local coordinate system of this hyperbola
        --        Returns the major axis of the hyperbola.


  YAxis (me)   returns Ax2d   is static;
        ---C++: inline
	--- Purpose : Computes an axis whose
        -- -   the origin is the center of this hyperbola, and
        -- -   the unit vector is the "X Direction" or "Y Direction"
        --  respectively of the local coordinate system of this hyperbola
        --  Returns the minor axis of the hyperbola.



  Reverse (me : in out)         is static;
        ---C++: inline

  Reversed (me)  returns Hypr2d  is static;
        ---C++: inline
        ---Purpose: Reverses the orientation of the local coordinate system
        -- of this hyperbola (the "Y Axis" is reversed). Therefore,
        -- the implicit orientation of this hyperbola is reversed.
        -- Note:
        -- -   Reverse assigns the result to this hyperbola, while
        -- -   Reversed creates a new one.
    
  IsDirect (me)  returns Boolean  is static;
        ---C++: inline
        --- Purpose : Returns true if the local coordinate system is direct
        --            and false in the other case.




  Mirror (me : in out; P : Pnt2d)            is static;

  Mirrored (me; P : Pnt2d)   returns Hypr2d  is static;

        --- Purpose :
        --  Performs the symmetrical transformation of an hyperbola with 
        --  respect  to the point P which is the center of the symmetry.



  Mirror (me : in out; A : Ax2d)             is static;

  Mirrored (me; A : Ax2d)   returns Hypr2d   is static;

        --- Purpose :
        --  Performs the symmetrical transformation of an hyperbola with 
        --  respect to an axis placement which is the axis of the symmetry.
      
  Rotate (me : in out; P : Pnt2d; Ang : Real)           is static;
        ---C++: inline
  
  Rotated (me; P : Pnt2d; Ang : Real)  returns Hypr2d   is static;
        ---C++: inline
        --- Purpose :
        --  Rotates an hyperbola. P is the center of the rotation.
        --  Ang is the angular value of the rotation in radians.
     
   

  Scale (me : in out; P : Pnt2d; S : Real)           is static;
        ---C++: inline

  Scaled (me; P : Pnt2d; S : Real)  returns Hypr2d   is static;
        ---C++: inline  
        --- Purpose : 
        --  Scales an hyperbola. <S> is the scaling value.
        --  If <S> is positive only the location point is 
        --  modified. But if <S> is negative the "XAxis" is 
        --  reversed and the "YAxis" too.   



  Transform (me : in out; T : Trsf2d)            is static;
        ---C++: inline

  Transformed (me; T : Trsf2d)  returns Hypr2d   is static;
        ---C++: inline
        --- Purpose :
        --  Transforms an hyperbola with the transformation T from 
        --  class Trsf2d.


  

  Translate (me : in out; V : Vec2d)            is static;
        ---C++: inline

  Translated (me; V : Vec2d)   returns Hypr2d   is static;
        ---C++: inline
        --- Purpose :
        --  Translates an hyperbola in the direction of the vector V.
        --  The magnitude of the translation is the vector's magnitude.


   
  Translate (me : in out; P1, P2 : Pnt2d)           is static;
        ---C++: inline

  Translated (me; P1, P2 : Pnt2d)   returns Hypr2d  is static;
        ---C++: inline
        --- Purpose :
        --  Translates an hyperbola from the point P1 to the point P2.


fields

  pos         : Ax22d;
  majorRadius : Real;
  minorRadius : Real;


end;

