-- Created on: 1991-02-21
-- Created by: Isabelle GRIGNON
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ExtSS from Extrema 
    	---Purpose: It calculates all the extremum distances
    	--          between two surfaces.
    	--          These distances can be minimum or maximum.

uses  	POnSurf           from Extrema,
    	ExtElSS           from Extrema,
    	Pnt               from gp,
	SurfaceType       from GeomAbs,
	SequenceOfPOnSurf from Extrema,
	SequenceOfReal    from TColStd,
	Surface           from Adaptor3d,
	SurfacePtr        from Adaptor3d
	

raises  NotDone      from StdFail,
    	OutOfRange   from Standard,
	TypeMismatch from Standard
	
	
is
    Create returns ExtSS;


    Create (S1, S2: Surface from Adaptor3d; TolS1, TolS2: Real)
    	returns ExtSS;
      	---Purpose: It calculates all the distances between S1 and S2.
    

    Create (S1, S2: Surface from Adaptor3d;
    	    Uinf1, Usup1, Vinf1, Vsup1: Real;
    	    Uinf2, Usup2, Vinf2, Vsup2: Real;
    	    TolS1, TolS2: Real)
    	returns ExtSS;
      	---Purpose: It calculates all the distances between S1 and S2.
    

    Initialize(me: in out; S2: Surface from Adaptor3d;
    	       Uinf2, Usup2, Vinf2, Vsup2: Real; TolS1: Real)
	---Purpose: Initializes the fields of the algorithm.
    
    is static;
    
    Perform(me: in out; S1: Surface from Adaptor3d; 
    	    Uinf1, Usup1, Vinf1, Vsup1: Real; TolS1: Real)
    	---Purpose: Computes the distances.
    	--          An exception is raised if the fieds have not been 
    	--          initialized.
    
    raises TypeMismatch from Standard
    is static;
    
    
    IsDone (me) returns Boolean
    	---Purpose: Returns True if the distances are found.
    	is static;
    
    IsParallel (me) returns Boolean
    	---Purpose: Returns True if the curve is on a parallel surface.
    	raises  NotDone from StdFail
    	    	-- if IsDone(me)=False.
    	is static;


    NbExt (me) returns Integer
    	---Purpose: Returns the number of extremum distances.
    	raises  NotDone from StdFail
	    	-- if IsDone(me)=False.
    	is static;

    SquareDistance (me; N: Integer) returns Real
    	---Purpose: Returns the value of the Nth resulting square distance.
    	raises  NotDone from StdFail,
    	    	-- if IsDone(me)=False.
    	        OutOfRange
		-- if N < 1 or N > NbPoints(me).
    	is static;

    Points (me; N: Integer; P1: out POnSurf; P2: out POnSurf) 
    	---Purpose: Returns the point of the Nth resulting distance.
    	raises  NotDone from StdFail,
    	    	-- if IsDone(me)=False.
    	        OutOfRange from Standard
		-- if N < 1 or N > NbPoints(me).
    	is static;

    Bidon(me) returns SurfacePtr from Adaptor3d
    is static private;


fields
    myS2     : SurfacePtr        from Adaptor3d;
    myDone   : Boolean           from Standard;
    myIsPar  : Boolean           from Standard;
    myExtElSS: ExtElSS           from Extrema;
    myPOnS1  : SequenceOfPOnSurf from Extrema;
    myPOnS2  : SequenceOfPOnSurf from Extrema;
    myuinf1  : Real              from Standard;
    myusup1  : Real              from Standard;
    myvinf1  : Real              from Standard;
    myvsup1  : Real              from Standard;
    myuinf2  : Real              from Standard;
    myusup2  : Real              from Standard;
    myvinf2  : Real              from Standard;
    myvsup2  : Real              from Standard;
    mytolS1  : Real              from Standard;
    mytolS2  : Real              from Standard;
    mySqDist : SequenceOfReal    from TColStd;
    myStype  : SurfaceType       from GeomAbs;

end ExtSS;
