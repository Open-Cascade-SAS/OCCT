-- Created on: 1991-01-14
-- Created by: Arnaud BOUZY
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class RelationIterator from Expr

	---Purpose: Iterates on every basic relation contained in
	--          a GeneralRelation.
        ---Level : Internal

uses GeneralRelation from Expr,
    SingleRelation from Expr,
    Array1OfSingleRelation from Expr

raises NoMoreObject from Standard,
    NoSuchObject from Standard

is

    Create(rel : GeneralRelation)
    returns RelationIterator;
    
    More(me)
    ---Purpose: Returns False if no other relation remains.
    returns Boolean
    is static;
    
    Next(me : in out)
    raises NoMoreObject
    is static;
    
    Value(me)
    ---Purpose: Returns current basic relation.
    --          Exception is raised if no more relation remains.
    returns  SingleRelation
    raises NoSuchObject
    is static;

fields

    myRelation : Array1OfSingleRelation;
    current : Integer;

end RelationIterator;
