-- Created on: 1993-12-08
-- Created by: Isabelle GRIGNON
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package ChFiKPart  

	---Purpose: Fonctions de remplissage pour une SurfData, dans
	--          les cas particulers de conges/chanfreins suivants :
	--          - cylindre/plan entre 2 surfaces planes,
	--          - tore/sphere/cone entre un plan et un cylindre othogonal,
	--          - tore/sphere/cone entre un plan et un cone othogonal,
	--          - tore/sphere/cone entre un plan et un tore othogonal,
	--          - tore/cone entre un plan et une sphere.

uses 
    ChFiDS, 
    TopOpeBRepDS,
    Adaptor2d,
    Adaptor3d,
    TopoDS,
    TopAbs,
    gp,
    TCollection,
    TColStd,
    Standard

is

    class RstMap instantiates DataMap from TCollection 
    	(Integer from Standard, 
    	 HCurve2d from Adaptor2d, 
    	 MapIntegerHasher  from  TColStd);

    class ComputeData;
    ---Purpose: Contient toutes  les   methodes de classe  destinees a
    --          remplir  une SurfData   dans  les  cas  particuliers
    --          enumeres ci-dessus.

end ChFiKPart;


