-- File:	StepFEA_FeaAreaDensity.cdl
-- Created:	Thu Dec 12 17:51:05 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class FeaAreaDensity from StepFEA
inherits FeaMaterialPropertyRepresentationItem from StepFEA

    ---Purpose: Representation of STEP entity FeaAreaDensity

uses
    HAsciiString from TCollection

is
    Create returns FeaAreaDensity from StepFEA;
	---Purpose: Empty constructor

    Init (me: mutable; aRepresentationItem_Name: HAsciiString from TCollection;
                       aFeaConstant: Real);
	---Purpose: Initialize all fields (own and inherited)

    FeaConstant (me) returns Real;
	---Purpose: Returns field FeaConstant
    SetFeaConstant (me: mutable; FeaConstant: Real);
	---Purpose: Set field FeaConstant

fields
    theFeaConstant: Real;

end FeaAreaDensity;
