-- Created on: 2000-11-21
-- Created by: Peter KURNEV
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class InterferenceLine from BOPTools 

	---Purpose: class for storing information about all  
    	---         interferences for given shape. 
	---         So,  for each shape in the DS, we will have 
        ---         the  following interference list 
	---         (i1, t1, r1), (i2, t2, r2),...(iN, tN, rN), 
	---         where    
	---         (iN, tN, rN) - object of type  BOPTools_Interference 
        ---         The  class 	BOPTools_InterferenceLine is  dedicated 
	---         to provide convinient tools to  manage this info. 
        --- 
	 
uses
    KindOfInterference from BooleanOperations, 
    ListOfInterference from BOPTools,
    Interference from BOPTools


is
    Create  
    	returns InterferenceLine from BOPTools; 
    	---Purpose:  
    	--- Empty constructor 
    	---
    GetOnType(me;  
    	    	    aType :KindOfInterference from BooleanOperations) 
    	returns ListOfInterference from BOPTools; 
    	---C++: return  const & 
    	---Purpose:  
    	--- Returns info. list for interferences of given type 
    	---
    IsComputed(me;  
    	    	    aWith :Integer from Standard; 
    	            aType :KindOfInterference from BooleanOperations) 
	returns Boolean from Standard; 
    	---Purpose:  
    	--- Returns  TRUE if the interference of type <aType> 
    	--- with the shape <aWith> has already been computed.           
    	---
    AddInterference  (me:out;  
    	    	    anInterference  :Interference from BOPTools);	    	  
    	---Purpose:  
    	--- Adds  info. about the Interference to the list
    	---
    AddInterference  (me:out;  
    	    	    aWith :Integer from Standard; 
    	            aType :KindOfInterference from BooleanOperations;  
    	    	    anIndex:Integer from Standard);
    	---Purpose:  
    	--- Adds  info. about the Interference to the list
    	---
    List(me) 
    	returns ListOfInterference from BOPTools;  
    	---C++: return const & 
    	---Purpose:  
    	--- Selector  
    	---
     RealList(me) 
    	returns ListOfInterference from BOPTools;  
    	---C++: return const & 
    	---Purpose:  
    	--- Selector     
    	---
    HasInterference(me)    	    
    	returns Boolean from Standard;       	
    	---Purpose:  
    	--- Returns  TRUE if the list contains at least one  interference   
    	--- with non-empty result            
    	---
fields
     
    myList            : ListOfInterference from BOPTools; 
    mySSList          : ListOfInterference from BOPTools; 
    myESList          : ListOfInterference from BOPTools; 
    myVSList          : ListOfInterference from BOPTools; 
    myEEList          : ListOfInterference from BOPTools; 
    myVEList          : ListOfInterference from BOPTools; 
    myVVList          : ListOfInterference from BOPTools; 
    myEmptyList       : ListOfInterference from BOPTools;  
    
end InterferenceLine;
