-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class SensitivePoly from Select3D 
inherits SensitiveEntity from Select3D

    ---Purpose: Sensitive Entity to make a face selectable.
    -- In some cases this class can raise Standard_ConstructionError and 
    -- Standard_OutOfRange exceptions from its member Select3D_PointData 
    -- mypolyg.

uses
    EntityOwner       from SelectBasics,
    Projector         from Select3D,
    ListOfBox2d       from SelectBasics,
    Array1OfPnt       from TColgp,
    HArray1OfPnt      from TColgp,
    Array1OfPnt2d     from TColgp,
    Box2d             from Select3D,
    PointData         from Select3D

raises    
    ConstructionError from Standard,
    OutOfRange        from Standard

is

    Initialize (OwnerId      : EntityOwner from SelectBasics;
            ThePoints    : Array1OfPnt from TColgp)
     returns mutable SensitivePoly;
        ---Level: Public 
        ---Purpose: Constructs a sensitive face object defined by the
        -- owner OwnerId, the array of points ThePoints, and
        -- the sensitivity type Sensitivity.
        -- The array of points is the outer polygon of the geometric face.

    Initialize (OwnerId      : EntityOwner from SelectBasics;
            ThePoints    : HArray1OfPnt from TColgp)
     returns mutable SensitivePoly;
        ---Level: Public 
        ---Purpose: Constructs a sensitive face object defined by the
        -- owner OwnerId, the array of points ThePoints, and
        -- the sensitivity type Sensitivity.
        -- The array of points is the outer polygon of the geometric face.

    Initialize(OwnerId      : EntityOwner from SelectBasics;
            NbOfPoints   : Integer = 6)
     returns mutable SensitivePoly;
        ---Level: Public 
        ---Purpose: Constructs the sensitive circle object defined by the
        -- owner OwnerId, the circle Circle, the Boolean
        -- FilledCircle and the number of points NbOfPoints. 

    Project (me:mutable;aProjector : Projector from Select3D) is redefined virtual;
    ---Level: Public 
    ---Purpose: projection of the sensitive primitive in order to
    --          get 2D boxes for the Sort Algorithm
    
    Areas   (me:mutable ; boxes : in out ListOfBox2d from SelectBasics) is redefined static;
    ---Level: Public 
    ---Purpose: stores in <boxes> the 2D Boxes which represent the sensitive face
    --          in the selection algorithm.

    Points3D(me:mutable; theHArrayOfPnt : in out HArray1OfPnt from TColgp);
    ---Purpose: Returns the 3D points of the array used at construction time.
    ---C++: inline

    Points2D(me:mutable; theArrayOfPnt2d : in out Array1OfPnt2d from TColgp);
    ---Purpose: Returns the 2D points of the array used at construction time.
    ---C++: inline

fields
 
    mybox2d         : Box2d     from Select3D is protected;
    mypolyg         : PointData from Select3D is protected;
end SensitivePoly;
