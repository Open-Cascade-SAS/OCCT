-- File:	BRepExtrema_DistanceSS.cdl
-- Created:	Wed Apr 17 16:03:05 1996
-- Author:	Maria PUMBORIOS
-- Author:      Herve LOUESSARD
--		<mps@sgi30>
---Copyright:	 Matra Datavision 1996
--           	 

private class DistanceSS from BRepExtrema


  ---Purpose:  This class allows to compute minimum distance between two shapes 
  -- (face edge vertex) and is used in DistShapeShape class. 

uses
  Shape   from  TopoDS,
  Box     from  Bnd,
  Vertex  from  TopoDS,
  Edge    from  TopoDS,
  Face    from  TopoDS,
  Pnt     from  gp,
  SeqOfSolution from BRepExtrema,
  Real from Standard

  
is 
  Create( S1: Shape from TopoDS; S2: Shape from TopoDS;
    	    B1, B2: Box from Bnd; DstRef: Real from Standard)
	---Purpose: computes the distance between two Shapes
        -- ( face edge vertex)        
  returns DistanceSS  from   BRepExtrema;
	              
  Create( S1: Shape from TopoDS; S2: Shape from TopoDS;
    	    B1, B2: Box from Bnd; DstRef: Real from Standard;
            aDeflection: Real from Standard)
	---Purpose: computes the distance between two Shapes
        -- ( face edge vertex). Parameter theDeflection is used 
        -- to specify a maximum deviation of extreme distances 
    	-- from the minimum one. 
    	-- Default value is Precision::Confusion().
  returns DistanceSS  from   BRepExtrema;


  Perform(me:in out; S1: Shape from TopoDS; S2: Shape from TopoDS;
    	  B1, B2: Box from Bnd; DstRef: Real from Standard)
	---Purpose: computes the distance between two Shapes
        -- ( face edge vertex)        
  is private;

  Perform (me:in out; S1: Vertex from TopoDS; S2: Vertex from TopoDS; 
    	    B1, B2: Box from Bnd; DstRef: Real from Standard)
	---Purpose:   computes the distance between two vertices  
  is private;


  Perform( me:in out;S1: Vertex from TopoDS; S2: Edge from TopoDS;
    	    B1, B2: Box from Bnd; DstRef: Real from Standard)
	---Purpose: computes the minimum distance between a vertex and an edge
 
  is private;      

  
  Perform( me:in out; S1: Vertex from TopoDS; S2: Face from TopoDS;
    	    B1, B2: Box from Bnd; DstRef: Real from Standard )
	---Purpose:computes the minimum distance between a vertex and a face  
  is private;

  
  Perform(me:in out; S1: Edge from TopoDS; S2: Vertex from TopoDS; 
    	    B1, B2: Box from Bnd; DstRef: Real from Standard)
	---Purpose: computes the minimum distance between an edge and a vertex  
  is private;

  Perform( me:in out;S1:Edge from TopoDS; S2: Edge from TopoDS; 
    	    B1, B2: Box from Bnd; DstRef: Real from Standard)
	    
	---Purpose:                        
  is private;

  Perform(me:in out; S1: Edge from TopoDS; S2: Face from TopoDS; 
    	    B1, B2: Box from Bnd; DstRef: Real from Standard )
	---Purpose:computes the minimum distance an edge and a face  
  is private; 

  Perform( me:in out; S1: Face from TopoDS; S2: Vertex from TopoDS; 
    	    B1, B2: Box from Bnd; DstRef: Real from Standard)
	---Purpose:computes the minimum distance betwwen a face and a vertex  
  is private;

  Perform( me: in out ;S1: Face from TopoDS; S2: Edge from TopoDS; 
    	    B1, B2: Box from Bnd; DstRef: Real from Standard)
	---Purpose:computes the minimum distance between a face and an edge  
                     
  is private;

  Perform( me:in out; S1: Face from TopoDS; S2: Face from TopoDS; 
    	    B1, B2: Box from Bnd ; DstRef: Real from Standard)
	---Purpose:computes the minimum distance between a face and a face   
                     
  is private;

  IsDone(me) returns Boolean from Standard;
    	---Purpose: True if the distance has been computed 

  
  DistValue(me) returns Real from Standard;
    	---Purpose: returns the distance value 
 
  Seq1Value(me) returns  SeqOfSolution from BRepExtrema;
  ---C++: return const& 
        ---Purpose : returns the list of solutions on the first shape
  
  Seq2Value(me) returns  SeqOfSolution from BRepExtrema; 
  ---C++: return const& 
       ---Purpose returns the list of solutions on the second shape 
        
 
fields

    SeqSolShape1 :  SeqOfSolution from BRepExtrema;
    SeqSolShape2 :  SeqOfSolution from BRepExtrema;  
    myDstRef: Real from Standard;
    myModif : Boolean from Standard;
    myEps   : Real    from Standard;
    

  
end;
