-- Created on: 1995-09-13
-- Created by: Marie Jose MARTZ
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class GeomEntity from GeomToIGES


    ---Purpose : provides methods to transfer Geom entity from CASCADE to IGES.

uses

    Real                     from Standard,
    IGESEntity               from IGESData,
    IGESModel                from IGESData

is

    Create 
    	returns GeomEntity from GeomToIGES;
    ---Purpose : Creates a tool GeomEntity

    Create(GE : GeomEntity from GeomToIGES)
        returns GeomEntity from GeomToIGES;
    ---Purpose : Creates a tool ready to run and sets its 
    --         fields as GE's.

    SetModel(me : in out; model : IGESModel from IGESData);
    ---Purpose : Set the value of "TheModel"

    GetModel(me) 
    	returns IGESModel from IGESData;
    ---Purpose : Returns the value of "TheModel"

    SetUnit(me: in out; unit: Real);
    ---Purpose : Sets the value of the UnitFlag 
    
    GetUnit(me)
    	returns Real from Standard;
    ---Purpose : Returns the value of the UnitFlag of the header of the model
    --           in meters.
    
fields

    TheModel      : IGESModel from IGESData ;

    TheUnitFactor : Real from Standard;

end GeomEntity;

