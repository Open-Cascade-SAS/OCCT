-- Created on: 1994-05-31
-- Created by: Christian CAILLET
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SelectFromSingleView  from IGESSelect  inherits SelectDeduct

    ---Purpose : This selection gets in all the model, the entities which are
    --           attached to the views given as input. Only Single Views are
    --           considered. This information is kept from Directory Part
    --           (View Item).

uses AsciiString from TCollection, EntityIterator, Graph

raises InterfaceError

is

    Create returns mutable SelectFromSingleView;
    ---Purpose : Creates a SelectFromSingleView

    RootResult (me; G : Graph) returns EntityIterator  raises InterfaceError;
    ---Purpose : Selects the Entities which are attached to the Single View(s)
    --           present in the Input

    Label (me) returns AsciiString from TCollection;
    ---Purpose : Returns the label, with is "Entities attached to single View"

end SelectFromSingleView;
