-- File:        Torus.cdl
-- Created:     Fri Dec  1 11:11:30 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class Torus from StepShape 

inherits GeometricRepresentationItem from StepGeom

uses

	Axis1Placement from StepGeom,
	Real from Standard, 
	HAsciiString from TCollection
is

	Create returns mutable Torus;
	---Purpose: Returns a Torus


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aPosition : mutable Axis1Placement from StepGeom;
	      aMajorRadius : Real from Standard;
	      aMinorRadius : Real from Standard) is virtual;

	-- Specific Methods for Field Data Access --

	SetPosition(me : mutable; aPosition : mutable Axis1Placement);
	Position (me) returns mutable Axis1Placement;
	SetMajorRadius(me : mutable; aMajorRadius : Real);
	MajorRadius (me) returns Real;
	SetMinorRadius(me : mutable; aMinorRadius : Real);
	MinorRadius (me) returns Real;

fields

	position : Axis1Placement from StepGeom;
	majorRadius : Real from Standard;
	minorRadius : Real from Standard;

end Torus;
