-- Created on: 1999-11-26
-- Created by: Andrey BETENEV
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0

class DateTimeItem from StepAP203
inherits SelectType from StepData

    ---Purpose: Representation of STEP SELECT type DateTimeItem

uses
    ProductDefinition from StepBasic,
    ChangeRequest from StepAP203,
    StartRequest from StepAP203,
    Change from StepAP203,
    StartWork from StepAP203,
    ApprovalPersonOrganization from StepBasic,
    Contract from StepBasic,
    SecurityClassification from StepBasic,
    Certification from StepBasic

is
    Create returns DateTimeItem from StepAP203;
	---Purpose: Empty constructor

    CaseNum (me; ent: Transient) returns Integer;
	---Purpose: Recognizes a kind of DateTimeItem select type
	--          1 -> ProductDefinition from StepBasic
	--          2 -> ChangeRequest from StepAP203
	--          3 -> StartRequest from StepAP203
	--          4 -> Change from StepAP203
	--          5 -> StartWork from StepAP203
	--          6 -> ApprovalPersonOrganization from StepBasic
	--          7 -> Contract from StepBasic
	--          8 -> SecurityClassification from StepBasic
	--          9 -> Certification from StepBasic
	--          0 else

    ProductDefinition (me) returns ProductDefinition from StepBasic;
	---Purpose: Returns Value as ProductDefinition (or Null if another type)

    ChangeRequest (me) returns ChangeRequest from StepAP203;
	---Purpose: Returns Value as ChangeRequest (or Null if another type)

    StartRequest (me) returns StartRequest from StepAP203;
	---Purpose: Returns Value as StartRequest (or Null if another type)

    Change (me) returns Change from StepAP203;
	---Purpose: Returns Value as Change (or Null if another type)

    StartWork (me) returns StartWork from StepAP203;
	---Purpose: Returns Value as StartWork (or Null if another type)

    ApprovalPersonOrganization (me) returns ApprovalPersonOrganization from StepBasic;
	---Purpose: Returns Value as ApprovalPersonOrganization (or Null if another type)

    Contract (me) returns Contract from StepBasic;
	---Purpose: Returns Value as Contract (or Null if another type)

    SecurityClassification (me) returns SecurityClassification from StepBasic;
	---Purpose: Returns Value as SecurityClassification (or Null if another type)

    Certification (me) returns Certification from StepBasic;
	---Purpose: Returns Value as Certification (or Null if another type)

end DateTimeItem;
