-- File:	QANewBRepNaming_Limitation.cdl
-- Created:	Tue Oct 31 14:42:07 2000
-- Author:	Vladislav ROMASHKO
--		<vro@flox.nnov.matra-dtv.fr>
---Copyright:	 Matra Datavision 2000

-- Lastly modified by :
-- +---------------------------------------------------------------------------+
-- !       szy ! Modified input parameter type           !18-10-2002! 3.0-00-2!
-- +---------------------------------------------------------------------------+

class Limitation from QANewBRepNaming inherits BooleanOperationFeat from QANewBRepNaming

uses

    Label from TDF, 
    MakeShape from BRepBuilderAPI,
    Limitation from QANewModTopOpe

is
 
    Create returns Limitation from QANewBRepNaming;

    Create(ResultLabel : Label from TDF) 
    returns Limitation from QANewBRepNaming;

    Load (me; MakeShape : in out Limitation from QANewModTopOpe); 
     
    LoadContent(me; MakeShape : in out Limitation from QANewModTopOpe)
    ---Purpose: Loads the content of the result.
    is protected;

    LoadResult(me; MakeShape : in out Limitation from QANewModTopOpe)
    ---Purpose: Loads the result.
    is protected;

    LoadDegenerated(me; MakeShape : in out Limitation from QANewModTopOpe)
    ---Purpose: Loads the deletion of the degenerated edges.
    is protected;    


    LoadWire(me; MakeShape : in out Limitation from QANewModTopOpe)
    ---Purpose: A default implementation for naming of a wire as an object of
    --          a boolean operation.
    is protected;

    LoadShell(me; MakeShape : in out Limitation from QANewModTopOpe)
    ---Purpose: A default implementation for naming of a shell as an object of
    --          a boolean operation.
    is protected;

end Limitation;

-- @@SDM: begin

-- Lastly modified by : vro                                    Date : 31-10-2000

-- File history synopsis (creation,modification,correction)
-- +---------------------------------------------------------------------------+
-- ! Developer !              Comments                   !   Date   ! Version  !
-- +-----------!-----------------------------------------!----------!----------+
-- !       vro ! Creation                                !31-10-2000!3.0-00-1!
-- !       szy ! Modified input parameter type of  Load  !18-10-2002! 3.0-00-2!
-- !  vladimir ! adaptation to CAS 5.0                   !  07/01/03!    4.0-2!
-- +---------------------------------------------------------------------------+
--
-- @@SDM: end
