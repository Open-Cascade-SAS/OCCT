-- Created on: 1993-01-26
-- Created by: Laurent PAINNOT
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package AdvApprox
    
     ---Purpose: This package provides algorithms approximating a function
     --          that can be multidimensional creating in the end a 
     --          BSpline function with the required continuity
     --          
               
uses gp,
     math,
     GeomAbs,
     TColStd, 
     TColgp, 
     TCollection, 
     Standard,
     StdFail, 
     PLib

    
is
    

    class ApproxAFunction from AdvApprox ;
    class SimpleApprox;
--  class ApproxAFunction;  

    imported EvaluatorFunction ;

    deferred class Cutting;

    class DichoCutting;

    class PrefCutting;

    class PrefAndRec;


end AdvApprox;
