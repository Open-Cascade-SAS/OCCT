-- Created on: 1992-05-21
-- Created by: Jean Claude VAUTHIER
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Curve from DrawTrSurf

inherits Drawable 
   
        --- Purpose :
        --  This class defines a drawable curve in 3d space.

uses Curve from Geom,
     Color from Draw,
     Display from Draw,
     Drawable3D from Draw,
     Interpretor from Draw,
     OStream

is




  Create (C : Curve from Geom; DispOrigin : Boolean from Standard = Standard_True)
        --- Purpose :
        --  creates a drawable curve from a curve of package Geom.
     returns Curve from DrawTrSurf;


  Create (C : Curve from Geom; aColor : Color from Draw; Discret : Integer;
          Deflection : Real; DrawMode : Integer;
    	  DispOrigin : Boolean from Standard = Standard_True;
          DispCurvRadius : Boolean  = Standard_False;
          RadiusMax : Real = 1.0e3;
	  RatioOfRadius : Real = 0.1)
     returns Curve from DrawTrSurf;


  DrawOn (me; dis : in out Display from Draw);
     

  GetCurve (me) returns any Curve from Geom
  ---C++: inline
  is static;

  SetColor(me : mutable; aColor : Color from Draw)
  ---C++: inline
  is static;

  DisplayOrigin(me) returns Boolean
  ---C++: inline
  is static;
    
  DisplayOrigin(me : mutable; V : Boolean)
  ---C++: inline
  is static;
    
  ShowCurvature(me : mutable)
        ---C++: inline
     is static;
     
  ClearCurvature(me : mutable)
        ---C++: inline
     is static;
  
  SetRadiusMax(me : mutable; Radius : Real)
        ---C++: inline
     is static;
     
  SetRadiusRatio(me : mutable;  Ratio : Real)
        ---C++: inline
     is static;
  Color (me)  returns Color from Draw
        ---C++: inline
     is static;
     
  RadiusMax(me)  returns Real
        ---C++: inline
     is static;
     
  RadiusRatio(me)  returns Real
        ---C++: inline
     is static;   
     
  Copy(me) returns Drawable3D from Draw
	---Purpose: For variable copy.
  is redefined;
  
  Dump(me; S : in out OStream)
	---Purpose: For variable dump.
  is redefined;

    Whatis(me; I : in out Interpretor from Draw)
    is redefined;
	---Purpose: For variable whatis command. Set  as a result  the
	--          type of the variable.

fields

  curv       : Curve   from Geom     is protected ;
  look       : Color   from Draw     is protected ;
  disporigin : Boolean from Standard is protected ;
  dispcurvradius : Boolean from Standard is protected ;
  radiusmax      : Real from  Standard is protected ;
  radiusratio    : Real from  Standard is protected ;  

end Curve;
