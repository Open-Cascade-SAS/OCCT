-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class BSplineSurface from StepGeom 

inherits BoundedSurface from StepGeom 


  -- N.B : EXPRESS Complexe SUBTYPE Declaration :

  -- ANDOR ( ONEOF ( b_spline_surface_with_knots uniform_surface quasi_uniform_surface bezier_surface ) rational_b_spline_surface ) 

uses

	Integer from Standard, 
	HArray2OfCartesianPoint from StepGeom, 
	BSplineSurfaceForm from StepGeom, 
	Logical from StepData, 
	CartesianPoint from StepGeom, 
	HAsciiString from TCollection
is

	Create returns BSplineSurface;
	---Purpose: Returns a BSplineSurface


	Init (me : mutable;
	      aName : HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      aName : HAsciiString from TCollection;
	      aUDegree : Integer from Standard;
	      aVDegree : Integer from Standard;
	      aControlPointsList : HArray2OfCartesianPoint from StepGeom;
	      aSurfaceForm : BSplineSurfaceForm from StepGeom;
	      aUClosed : Logical from StepData;
	      aVClosed : Logical from StepData;
	      aSelfIntersect : Logical from StepData) is virtual;

	-- Specific Methods for Field Data Access --

	SetUDegree(me : mutable; aUDegree : Integer);
	UDegree (me) returns Integer;
	SetVDegree(me : mutable; aVDegree : Integer);
	VDegree (me) returns Integer;
	SetControlPointsList(me : mutable; aControlPointsList : HArray2OfCartesianPoint);
	ControlPointsList (me) returns HArray2OfCartesianPoint;
	ControlPointsListValue (me; num1 : Integer;  num2 : Integer) returns CartesianPoint;
	NbControlPointsListI (me) returns Integer;
	NbControlPointsListJ (me) returns Integer;
	SetSurfaceForm(me : mutable; aSurfaceForm : BSplineSurfaceForm);
	SurfaceForm (me) returns BSplineSurfaceForm;
	SetUClosed(me : mutable; aUClosed : Logical);
	UClosed (me) returns Logical;
	SetVClosed(me : mutable; aVClosed : Logical);
	VClosed (me) returns Logical;
	SetSelfIntersect(me : mutable; aSelfIntersect : Logical);
	SelfIntersect (me) returns Logical;

fields

	uDegree : Integer from Standard;
	vDegree : Integer from Standard;
	controlPointsList : HArray2OfCartesianPoint from StepGeom;
	surfaceForm : BSplineSurfaceForm from StepGeom; -- an Enumeration
	uClosed : Logical from StepData;
	vClosed : Logical from StepData;
	selfIntersect : Logical from StepData;

end BSplineSurface;
