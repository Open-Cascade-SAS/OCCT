-- Created on: 1993-04-06
-- Created by: Philippe DAUTRY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Line from PGeom2d inherits Curve from PGeom2d

        ---Purpose :   Defines   an   infinite   line.  	   The
        --         parametrization range is ]-infinite, +infinite[.
        --         
	---See Also : Line from Geom2d.

uses Ax2d from gp

is


  Create returns Line;
        ---Purpose : Creates a line with default values.
	---Level: Internal 


  Create (aPosition : Ax2d from gp)   returns Line;
        ---Purpose : Creates   a  line  located    in  3D space   with
        --         <aPosition>.  The Location   of <aPosition> is  the
        --         origin of the line.
	---Level: Internal 


  Position (me : mutable; aPosition : Ax2d from gp);
        --- Purpose : Set the value of the field position with <aPosition>.
	---Level: Internal 


  Position (me) returns Ax2d from gp;
        --- Purpose : Returns the value of the field position.
	---Level: Internal 


fields

  position : Ax2d from gp;

end;
