-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class CsgPrimitive from StepShape inherits SelectType from StepData

	-- <CsgPrimitive> is an EXPRESS Select Type construct translation.
	-- it gathers : Sphere, Block, RightAngularWedge, Torus, RightCircularCone, RightCircularCylinder

uses

	Sphere,
	Block,
	RightAngularWedge,
	Torus,
	RightCircularCone,
	RightCircularCylinder
is

	Create returns CsgPrimitive;
	---Purpose : Returns a CsgPrimitive SelectType

	CaseNum (me; ent : Transient) returns Integer;
	---Purpose: Recognizes a CsgPrimitive Kind Entity that is :
	--        1 -> Sphere
	--        2 -> Block
	--        3 -> RightAngularWedge
	--        4 -> Torus
	--        5 -> RightCircularCone
	--        6 -> RightCircularCylinder
	--        0 else

	Sphere (me) returns any Sphere;
	---Purpose : returns Value as a Sphere (Null if another type)

	Block (me) returns any Block;
	---Purpose : returns Value as a Block (Null if another type)

	RightAngularWedge (me) returns any RightAngularWedge;
	---Purpose : returns Value as a RightAngularWedge (Null if another type)

	Torus (me) returns any Torus;
	---Purpose : returns Value as a Torus (Null if another type)

	RightCircularCone (me) returns any RightCircularCone;
	---Purpose : returns Value as a RightCircularCone (Null if another type)

	RightCircularCylinder (me) returns any RightCircularCylinder;
	---Purpose : returns Value as a RightCircularCylinder (Null if another type)


end CsgPrimitive;

