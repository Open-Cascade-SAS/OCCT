-- Created on: 2000-05-10
-- Created by: Andrey BETENEV
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1

class ExternalIdentificationAssignment from StepBasic
inherits IdentificationAssignment from StepBasic

    ---Purpose: Representation of STEP entity ExternalIdentificationAssignment

uses
    HAsciiString from TCollection,
    IdentificationRole from StepBasic,
    ExternalSource from StepBasic

is
    Create returns ExternalIdentificationAssignment from StepBasic;
	---Purpose: Empty constructor

    Init (me: mutable; aIdentificationAssignment_AssignedId: HAsciiString from TCollection;
                       aIdentificationAssignment_Role: IdentificationRole from StepBasic;
                       aSource: ExternalSource from StepBasic);
	---Purpose: Initialize all fields (own and inherited)

    Source (me) returns ExternalSource from StepBasic;
	---Purpose: Returns field Source
    SetSource (me: mutable; Source: ExternalSource from StepBasic);
	---Purpose: Set field Source

fields
    theSource: ExternalSource from StepBasic;

end ExternalIdentificationAssignment;
