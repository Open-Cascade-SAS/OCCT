-- Created on: 1994-10-03
-- Created by: Assim
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ShapeBinder  from TransferBRep  inherits BinderOfShape

    ---Purpose : A ShapeBinder is a BinderOfShape with some additional services
    --           to cast the Result under various kinds of Shapes

uses  ShapeEnum from TopAbs,  Shape from TopoDS ,
      Vertex from TopoDS,  Edge  from TopoDS,  Wire  from TopoDS,
      Face   from TopoDS,  Shell from TopoDS,  Solid from TopoDS,
      CompSolid from TopoDS,    Compound from TopoDS

raises TypeMismatch from Standard

is

    Create returns mutable ShapeBinder;
    ---Purpose : Creates an empty ShapeBinder

    Create (res : Shape) returns mutable ShapeBinder;
    ---Purpose : Creates a ShapeBinder with a result

    ShapeType (me) returns ShapeEnum;
    ---Purpose : Returns the Type of the Shape Result (under TopAbs form)

    -- different sub-types for the Result. Result returns a Shape

    Vertex    (me) returns Vertex    raises TypeMismatch from Standard;
    Edge      (me) returns Edge      raises TypeMismatch from Standard;
    Wire      (me) returns Wire      raises TypeMismatch from Standard;
    Face      (me) returns Face      raises TypeMismatch from Standard;
    Shell     (me) returns Shell     raises TypeMismatch from Standard;
    Solid     (me) returns Solid     raises TypeMismatch from Standard;
    CompSolid (me) returns CompSolid raises TypeMismatch from Standard;
    Compound  (me) returns Compound  raises TypeMismatch from Standard;

end ShapeBinder;
