-- Created on: 1996-01-26
-- Created by: Philippe MANGIN
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



private class BattenLaw from FairCurve inherits Function from math

	---Purpose: This class compute the Heigth of an batten 

is
     Create(Heigth, Slope, Sliding : Real)
    ---Purpose: Constructor of linear batten with
    --          Heigth : the Heigth at the middle point
    --          Slope  : the geometric slope of the batten
    --          Sliding : Active Length of the batten without extension
     returns BattenLaw;
     
     SetSliding(me : in out; Sliding : Real);
     ---Purpose: Change the value of sliding
     ---C++: inline
     
     SetHeigth(me : in out; Heigth : Real);
     ---Purpose: Change the value of Heigth at the middle point.
     ---C++: inline
     
     SetSlope(me : in out; Slope : Real);
     ---Purpose: Change the value of the geometric slope.
     ---C++: inline
     
    
     Value(me: in out; T: Real; THeigth: out Real) returns Boolean
     ---Purpose: computes the value of  the heigth for the parameter T
     --          on  the neutral fibber
     ---C++: inline
     is redefined;




fields
MiddleHeigth   : Real; -- the Heigth at the middle point
GeometricSlope : Real; -- the geometric slope of the batten
LengthSliding  : Real; -- the length of sliding of the batten
end BattenLaw;
