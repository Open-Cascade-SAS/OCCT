-- File:	QANewBRepNaming_Chamfer.cdl
-- Created:	Mon Sep 22 15:59:33 1997
-- Author:	VAUTHIER Jean-Claude
---Copyright:	 Matra Datavision 1997


class Chamfer from QANewBRepNaming inherits TopNaming from QANewBRepNaming

    ---Purpose: To load the Chamfer results

uses 
 
    MakeChamfer from BRepFilletAPI,
    Shape       from TopoDS,
    Label       from TDF

is
 
    Create returns Chamfer from QANewBRepNaming; 

    Create(ResultLabel : Label from TDF) 
    returns Chamfer from QANewBRepNaming; 

    Init(me : in out; ResultLabel :  Label from TDF);


    Load (me; part      : in     Shape       from TopoDS;
    	      mkChamfer : in out MakeChamfer from BRepFilletAPI);

    FacesFromEdges (me) 
    ---Purpose: Returns the label of faces generated from edges
    returns Label from TDF;
    
    ModifiedFaces (me)
    ---Purpose: Returns the label of modified faces 
    returns Label from TDF;

    DeletedFaces (me)
    ---Purpose: Returns the label of deleted faces 
    returns Label from TDF;

end Chamfer;
