-- Created on: 1994-04-18
-- Created by: Laurent BUCHARD
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



package BRepClass3d 

uses  
    gp,
    TopAbs,
    TopoDS,
    TopTools,
    TCollection,
    TopExp,
    TopClass,
    BRepClass,
    Geom2dInt,
    IntCurveSurface,
    IntCurvesFace,
    Bnd,
    BRepAdaptor


is

    class Intersector3d;

    class MapOfInter instantiates  
       DataMap from TCollection(Shape          from TopoDS,
	    	    	    	Address        from Standard,
                                ShapeMapHasher from TopTools);
				

    class SolidExplorer;
        
    class SolidPassiveClassifier instantiates Classifier3d from TopClass
    	(Intersector3d  from BRepClass3d);

    ---class SClassifier instantiates SolidClassifier from TopClass
    ---   (SolidExplorer from BRepClass3d,
    ---	Intersector3d from BRepClass3d);
     
    
    class SClassifier;       

    class SolidClassifier;
    
       
       
end BRepClass3d;
