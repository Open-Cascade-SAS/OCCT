-- Created on: 1997-02-06
-- Created by: Denis PASCAL
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Integer from TDataStd inherits Attribute from TDF

	---Purpose:  The basis to define an integer attribute.

uses Attribute       from TDF,
     Label           from TDF,
     GUID            from Standard,
     Integer         from Standard,
     RelocationTable from TDF

is 

    ---Purpose: class methods
    --          =============

    GetID (myclass)   
        ---C++: return const & 
	---Purpose: Returns the GUID for integers.  
    returns GUID from Standard;

    Set (myclass; label : Label from TDF; value : Integer from Standard)
    ---Purpose: Finds, or creates, an Integer attribute and sets <value>
    --          the Integer  attribute is returned.
    returns Integer from TDataStd;

    ---Purpose: Integer methods
    --          ===============
    
    Set (me : mutable; V : Integer from Standard);
    
    Get (me)
    returns Integer from Standard;
    ---Purpose: Returns the integer value contained in the attribute.
    IsCaptured(me) returns Boolean;
	---Purpose: Returns True if there is a reference on the same label

    ---Category: methodes de TDF_Attribute
    --           =========================
    
    ID (me)
    	---C++: return const & 
    returns GUID from Standard;

    Restore (me: mutable; With : Attribute from TDF);

    NewEmpty (me)
    returns mutable Attribute from TDF;

    Paste (me; Into : mutable Attribute from TDF;
	       RT   : mutable RelocationTable from TDF);    

    Dump(me; anOS : in out OStream from Standard)
    	returns OStream from Standard
    	is redefined;
	---C++: return &


    Create
    returns mutable Integer from TDataStd;    


fields

    myValue : Integer from Standard;

end Integer;
