-- Created on: 1995-12-04
-- Created by: Laurent BOURESCHE
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class CoonsAlgPatch from GeomFill inherits TShared from MMgt

	---Purpose: Provides  evaluation   methods on an   algorithmic
	--          patch   defined by  its   boundaries and  blending
	--          functions.

uses
    Pnt              from gp,
    Vec              from gp,
    Boundary         from GeomFill,
    Function         from Law

is

    Create(B1, B2, B3, B4 : Boundary from GeomFill) 
    ---Purpose: Constructs the  algorithmic   patch. By   Default  the
    --          constructed blending functions are linear.
    --  Warning: No control is done on the bounds.
    --          B1/B3 and B2/B4 must be same range and well oriented.
    returns mutable CoonsAlgPatch  from  GeomFill;

    Func(me;
         f1,f2 : out Function from Law)
    ---Purpose: Give the blending functions.

    is static;

    SetFunc(me    : mutable;
            f1,f2 : Function from Law)
    ---Purpose: Set the blending functions.

    is static;

    Value(me;
          U,V : Real from Standard) returns Pnt from gp
    ---Purpose: Computes  the  value   on the  algorithmic    patch at
    --          parameters U and V.
    is static;
    
    D1U(me;
    	U,V : Real from Standard)
    returns Vec from gp
    ---Purpose: Computes   the  d/dU   partial   derivative  on    the
    --          algorithmic patch at parameters U and V.
    is static;

    D1V(me;
    	U,V : Real from Standard)
    returns Vec from gp
    ---Purpose: Computes    the  d/dV    partial    derivative on  the
    --          algorithmic patch at parameters U and V.
    is static;

    DUV(me;
    	U,V : Real from Standard)
    returns Vec from gp
    ---Purpose: Computes the   d2/dUdV  partial  derivative   on   the
    --          algorithmic  patch made with linear blending functions
    --          at parameter U and V.
    is static;

    Corner(me; I : Integer from Standard) 
    ---C++: return const&
    returns Pnt from gp
    is static;

    Bound(me; I : Integer from Standard) 
    ---C++: return const&
    returns any Boundary from GeomFill
    is static;

    Func(me; I : Integer from Standard) 
    ---C++: return const&
    returns any Function from Law
    is static;

fields

    -- the boundaries.
    bound : Boundary from GeomFill [4];
    
    -- the corners.
    c   : Pnt from gp [4];
    
    -- the   blending functions.
    a : Function from Law [2];
    
end CoonsAlgPatch;
