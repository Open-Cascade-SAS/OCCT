-- Created on: 2009-03-20
-- Created by: ABD
-- Copyright (c) 2009-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

private class ColorScaleLayerItem from V3d inherits LayerItem from Visual3d

    ---Version:

    ---Purpose: This class is drawable unit of ColorScale of 2d scene
    ---Keywords:
    ---Warning:
    ---References:

uses
    ColorScale from V3d
is
    -------------------------
    -- Category: Constructors
    -------------------------

    Create ( aColorScale: ColorScale from V3d )
            returns ColorScaleLayerItem;
    ---Level: Public
    ---Purpose: Creates a layer item
    ---Category: Constructors

    ---------------------------------------------------
    -- Category: Methods to modify the class definition
    ---------------------------------------------------
    
    ComputeLayerPrs( me : mutable )
            is redefined;   
    ---Level: Public
    ---Purpose: virtual function for recompute 2D
    --        presentation (empty by default)

    RedrawLayerPrs( me : mutable )
        is redefined;
    ---Level: Public
    ---Purpose: virtual function for recompute 2D
    --        presentation (empty by default)

fields
    MyColorScale     : ColorScale from V3d;

end ColorScaleLayerItem from V3d;
