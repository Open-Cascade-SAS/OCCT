-- File:        SurfaceStyleControlGrid.cdl
-- Created:     Mon Dec  4 12:02:31 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWSurfaceStyleControlGrid from RWStepVisual

	---Purpose : Read & Write Module for SurfaceStyleControlGrid

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     SurfaceStyleControlGrid from StepVisual,
     EntityIterator from Interface

is

	Create returns RWSurfaceStyleControlGrid;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable SurfaceStyleControlGrid from StepVisual);

	WriteStep (me; SW : in out StepWriter; ent : SurfaceStyleControlGrid from StepVisual);

	Share(me; ent : SurfaceStyleControlGrid from StepVisual; iter : in out EntityIterator);

end RWSurfaceStyleControlGrid;
