-- Created on: 1996-01-22
-- Created by: Philippe MANGIN
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class GaussSetIntegration from math
    ---Purpose: -- This class implements the integration of a set of N
    --              functions of M  variables variables between the
    --              parameter bounds Lower[a..b] and Upper[a..b].
    --  Warning: - The case M>1 is not implemented.


uses Vector from math,
     IntegerVector from math, 
     FunctionSet from math,
     OStream from Standard,
     NotDone from StdFail

raises NotDone, NotImplemented

is

     Create(F: in out FunctionSet; Lower, Upper: Vector;
     	    Order: IntegerVector)
     ---Purpose:
     -- The Gauss-Legendre integration with Order = points of 
     -- integration for each unknow, is done on the function F 
     -- between the bounds Lower and Upper.
     returns GaussSetIntegration     
     raises  NotImplemented;
     
     IsDone(me)
     	---Purpose: returns True if all has been correctly done.
    	---C++: inline

     returns Boolean
     is static;
     
     Value(me)
     	---Purpose: returns the value of the integral.
    	---C++: inline
    	---C++: return const&

     returns Vector
     raises NotDone
     is static;


    Dump(me; o: in out OStream)
    	---Purpose: Prints information on the current state of the object.
    is static;




fields

Val: Vector;
Done: Boolean;

end GaussSetIntegration;
