-- Created on: 1994-06-24
-- Created by: Yves FRICAUD
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Inter from Bisector 

	---Purpose: Intersection between two <Bisec> from Bisector.

inherits 
    Intersection from IntRes2d
    
uses   
    Domain  from IntRes2d,
    Bisec   from Bisector,
    Curve   from Bisector,
    BisecCC from Bisector,
    Curve   from Geom2d,
    Line    from Geom2d
    
raises ConstructionError from Standard

is
    Create returns Inter from Bisector;
    
    Create (C1: Bisec from Bisector; D1: Domain from IntRes2d;
            C2: Bisec from Bisector; D2: Domain from IntRes2d;
    	    TolConf,Tol  : Real    from Standard;
    	    ComunElement : Boolean from Standard) 
	---Purpose: Intersection between 2 curves.  
	--          C1 separates the element A and B. 
	--          C2 separates the elements C et D.
	--          If B an C have the same geometry. <ComunElement>
	--          Has to be True. 
	--          It Permits an optimiztion of the computation.

    returns  Inter from Bisector
    raises   ConstructionError from Standard;

    
    Perform (me: in out;
             C1: Bisec from Bisector; D1: Domain from IntRes2d;
             C2: Bisec from Bisector; D2: Domain from IntRes2d;
    	     TolConf,Tol  : Real    from Standard;
    	     ComunElement : Boolean from Standard) 
	---Purpose: Intersection between 2 curves.          
    	--          C1 separates the element A and B. 
	--          C2 separates the elements C et D.
	--          If B an C have the same geometry. <ComunElement>
	--          Has to be True. 
	--          It Permits an optimiztion of the computation.

    raises   ConstructionError from Standard
    is static;
    
    SinglePerform (me: in out;
             	   C1: Curve from Geom2d ; D1: Domain from IntRes2d;
             	   C2: Curve from Geom2d ; D2: Domain from IntRes2d;
    	           TolConf,Tol  : Real    from Standard;
    	           ComunElement : Boolean from Standard) 
	---Purpose: Intersection between 2 curves.          
    
    raises   ConstructionError from Standard
    is static private;
	
    NeighbourPerform (me : in out;
    	    	      C1 : BisecCC from Bisector; D1: Domain from IntRes2d;
                      C2 : BisecCC from Bisector; D2: Domain from IntRes2d;
    	              Tol: Real    from Standard)
    is static private;
    
    TestBound (me : in out;
    	       C1 : Line  from Geom2d  ; D1      : Domain  from IntRes2d;
    	       C2 : Curve from Geom2d  ; D2      : Domain  from IntRes2d;
	       Tol: Real  from Standard; Reverse : Boolean from Standard)
    is static private;
    
end Inter;
