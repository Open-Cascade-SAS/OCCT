-- Created on: 1992-08-26
-- Created by: Jean Louis FRENKEL
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


package Prs3d

    	---Purpose: The Prs3d package provides the following services
	-- -   a presentation object (the context for all
	--   modifications to the display, its presentation will be
	--   displayed in every view of an active viewer)
	-- -   an attribute manager governing how objects such
	--   as color, width, and type of line are displayed;
	--   these are generic objects, whereas those in
	--   StdPrs are specific geometries and topologies.
	-- -   generic   algorithms providing default settings for
	--   objects such as points, curves, surfaces and shapes
	-- -   a root object which provides the abstract
	--   framework for the DsgPrs definitions at work in
	--   display of dimensions, relations and trihedra.
    
uses
  Graphic3d,
  Aspect,
  Quantity,
  MMgt,
  Standard,
  Adaptor3d,
  BRepAdaptor,
  Geom,
  CPnts,
  GCPnts,
  TopAbs,
  TopLoc,
  TopoDS,
  TopTools,
  TopExp,
  HLRAlgo,
  TCollection,
  TColgp,
  Bnd,
  gp,
  Poly,
  TColStd
is  
  exception InvalidAngle inherits RangeError from Standard;

  enumeration TypeOfLinePicking is TOLP_Point,
                                   TOLP_Segment
  end TypeOfLinePicking;
        
  enumeration TypeOfHLR is TOH_NotSet,
                           TOH_PolyAlgo,
                           TOH_Algo;
  ---Purpose: Declares types of hidden line removal algorithm.
  --          TOH_Algo enables using of exact HLR algorithm.
  --          TOH_PolyAlgo enables using of polygonal HLR algorithm.
  --          TOH_NotSet is used by AIS_Drawer class, it means that the drawer should return the global value.
  --          For more details see AIS_Drawer class, AIS_Shape::Compute() method and
  --          HLRAlgo package from TKHLR toolkit.
  
  enumeration DimensionTextHorizontalPosition is DTHP_Left, DTHP_Right, DTHP_Center, DTHP_Fit;
  ---Purpose: Specifies options for positioning dimension value label in horizontal direction.
  -- DTHP_Left   - value label located at left side on dimension extension.
  -- DTHP_Right  - value label located at right side on dimension extension.
  -- DTHP_Center - value label located at center of dimension line.
  -- DTHP_Fit    - value label located automatically at left side if does not fits
  --               the dimension space, otherwise the value label is placed at center.

  enumeration DimensionTextVerticalPosition is DTVP_Above, DTVP_Below, DTVP_Center;
  ---Purpose: Specifies options for positioning dimension value label in vertical direction
  -- with respect to dimension (extension) line.
  -- DTVP_Above - text label is located above the dimension or extension line.
  -- DTVP_Below - text label is located below the dimension or extension line.
  -- DTVP_Center - the text label middle-point is in line with dimension or extension line.

  enumeration DimensionArrowOrientation is DAO_Internal, DAO_External, DAO_Fit;
  ---Purpose: Specifies dimension arrow location and orientation.
  -- DAO_Internal - arrows "inside", pointing outwards.
  -- DAO_External - arrows "outside", pointing inwards.
  -- DAO_Fit      - arrows oriented inside if value label with arrowtips fit the dimension line,
  --                otherwise - externally

  class Presentation;
  ---Purpose: defines the presentation object. This object can be
  --          displayed, highlighted, erased, etc... The output
  --          of the presentation algorithms are sent in a
  --          presentation object. A presentation object is attached
  --          to a given Viewer.

	---Category: Aspect classes.
	---Purpose: The aspect classes qualifies how to represent
	--          a given kind of object.
	--          

  deferred class BasicAspect;	
  class PointAspect;
  class LineAspect;
	class ShadingAspect;
	class TextAspect;
  class IsoAspect;
  class ArrowAspect;
	class PlaneAspect;
  class DimensionAspect;
	class DatumAspect;

  class Drawer;
	---Purpose: qualifies how the presentation algorithms compute
	--          the presentation of a specific kind of object. 
	--          This includes for example color, width and type
	--          of lines, maximal chordial deviation, etc...
	--          A drawer includes an instance of the Aspect classes
	--          with particular default values.
	
  class Projector;
	---Purpose: defines the projection parameters for the hidden
	--          lines removal algorithm.
	
  class PlaneSet;
	---Purpose: defines a set of planes used for a presentation
	--          by sections.
	-- 

  deferred class Root;
	---Purpose: defines the root of the presentation algorithms.

  ---Category: Basis construction elements.

	class Text;

        ---Category: Class signatures.

	class ShapeTool;
	---Purpose: describes the behaviour requested for a wireframe
	--          shape presentation.

  class Arrow;
	---Purpose: draws an arrow at a given location, with respect
	--          to a given direction. 

  imported NListOfSequenceOfPnt; 
  imported NListIteratorListOfSequenceOfPnt;
  imported Point;
  imported WFShape;
  
  MatchSegment(X,Y,Z: Length from Quantity;
	            aDistance: Length from Quantity;
		          p1,p2: Pnt from gp;
              dist: out Length from Quantity)
	returns Boolean from Standard;
end Prs3d;
