-- Created on: 1993-04-23
-- Created by: Modelistation
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SLPropsATool from HLRBRep

uses
    Address from Standard,
    Pnt     from gp,
    Vec     from gp

is

    Value(myclass; A    :     Address from Standard; 
    	    	   U, V :     Real    from Standard;
                   P    : out Pnt     from gp);
    	---Purpose: Computes the point  <P> of 	parameter <U> and <V>
    	--          on the Surface <A>.
    	--
    	---C++: inline

    D1   (myclass; A        : Address from Standard;
                   U, V     : Real    from Standard;
                   P        : out Pnt from gp;
                   D1U, D1V : out Vec from gp);
    	---Purpose: Computes the point <P>  and first derivative <D1*>
    	--          of parameter <U> and <V> on the Surface <A>.
    	--          
    	---C++: inline

    D2   (myclass; A    : Address from Standard;
                   U, V : Real    from Standard; 
              P : out Pnt; D1U, D1V, D2U, D2V, DUV : out Vec);
    	---Purpose: Computes the point <P>, the first derivative <D1*>
    	--          and second  derivative <D2*> of parameter  <U> and
    	--          <V> on the Surface <A>.
    	--          
       	---C++: inline

    DN   (myclass; A      : Address from Standard;
                   U, V   : Real    from Standard;
		   Nu, Nv : Integer from Standard)
    returns Vec from gp;

    Continuity(myclass; A : Address from Standard)
    returns Integer from Standard;
    	---Purpose: returns the order of   continuity of the   Surface
    	--          <A>.  returns  1   :  first  derivative    only is
    	--          computable returns 2 : first and second derivative
    	--          only are computable.
    	--          
       	---C++: inline

    Bounds(myclass; A              :     Address from Standard;
                    U1, V1, U2, V2 : out Real    from Standard);
    	---Purpose: returns the bounds of the Surface.
    	--          
    	---C++: inline

end SLPropsATool;
