-- Created on: 2000-05-10
-- Created by: Andrey BETENEV
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1

class EffectivityAssignment from StepBasic
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity EffectivityAssignment

uses
    Effectivity from StepBasic

is
    Create returns EffectivityAssignment from StepBasic;
	---Purpose: Empty constructor

    Init (me: mutable; aAssignedEffectivity: Effectivity from StepBasic);
	---Purpose: Initialize all fields (own and inherited)

    AssignedEffectivity (me) returns Effectivity from StepBasic;
	---Purpose: Returns field AssignedEffectivity
    SetAssignedEffectivity (me: mutable; AssignedEffectivity: Effectivity from StepBasic);
	---Purpose: Set field AssignedEffectivity

fields
    theAssignedEffectivity: Effectivity from StepBasic;

end EffectivityAssignment;
