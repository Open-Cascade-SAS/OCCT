-- Created on: 1993-01-13
-- Created by: CKY / Contract Toubro-Larsen ( Deepak PRABHU )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class MacroDef from IGESDefs  inherits IGESEntity

        ---Purpose: defines IGES Macro Definition Entity, Type <306> Form <0>
        --          in package IGESDefs
        --          This Class specifies the action of a specific MACRO.
        --          After specification MACRO can be used as necessary
        --          by means of MACRO class instance entity.

uses

        HAsciiString          from TCollection,
        HArray1OfHAsciiString from Interface

raises OutOfRange

is

        Create returns mutable MacroDef;

        -- Specific methods for the entity

        Init (me             : mutable;
              macro          : HAsciiString;
              entityTypeID   : Integer;
              langStatements : HArray1OfHAsciiString;
              endMacro       : HAsciiString);
        ---Purpose : This method is used to set the fields of the class
        --           MacroDef
        --       - macro          : MACRO
        --       - entityTypeID   : Entity Type ID
        --       - langStatements : Language Statements
        --       - endMacro       : END MACRO

        NbStatements(me) returns Integer;
        ---Purpose : returns the number of language statements

        MACRO(me) returns HAsciiString from TCollection;
        ---Purpose : returns the MACRO(Literal)

        EntityTypeID(me) returns Integer;
        ---Purpose : returns the Entity Type ID

        LanguageStatement(me ; StatNum : Integer) 
        returns HAsciiString from TCollection
        raises OutOfRange;
        -- returns the StatNum'th statement
        -- raises exception if StatNum <= 0 or StatNum > NbStatements()

        ENDMACRO(me) returns HAsciiString from TCollection;
        ---Purpose : returns the ENDM(Literal)

fields

--
--  Class    : IGESDefs_MacroDef
--
--  Purpose  : Declaration of variables specific to MacroDef
--
--  Reminder : An MacroDef Entity specifies the action of a
--             specific MACRO. It consists of only language
--             statements in the parameter data.

        theMACRO          : HAsciiString;
        theEntityTypeID   : Integer;
        theLangStatements : HArray1OfHAsciiString;
        theENDMACRO       : HAsciiString;

end MacroDef;
