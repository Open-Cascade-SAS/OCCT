-- Created on: 1994-09-02
-- Created by: Christian CAILLET
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class PacketList  from IFSelect  inherits TShared

    ---Purpose : This class gives a simple way to return then consult a
    --           list of packets, determined from the content of a Model,
    --           by various criteria.
    --           
    --           It allows to describe several lists with entities from a
    --           given model, possibly more than one list knowing every entity,
    --           and to determine the remaining list (entities in no lists) and
    --           the duplications (with their count).

uses Array1OfInteger, IntList, HSequenceOfTransient, AsciiString,
     EntityIterator, InterfaceModel

raises InterfaceError

is

    Create (model : InterfaceModel) returns mutable PacketList;
    ---Purpose : Creates a PackList, empty, ready to receive entities from a
    --           given Model

    SetName (me : mutable; name : CString)  is static;
    ---Purpose : Sets a name to a packet list : this makes easier a general
    --           routine to print it. Default is "Packets"

    Name (me) returns CString  is static;
    ---Purpose : Returns the recorded name for a packet list

    Model (me) returns InterfaceModel;
    ---Purpose : Returns the Model of reference

    AddPacket (me : mutable);
    ---Purpose : Declares a new Packet, ready to be filled
    --           The entities to be added will be added to this Packet

    Add (me : mutable; ent : Transient)
    ---Purpose : Adds an entity from the Model into the current packet for Add
    	raises InterfaceError;
    --           Error if <ent> is not from the Model, or if no AddPacket was
    --           yet called

    AddList (me : mutable; list : HSequenceOfTransient)
    ---Purpose : Adds an list of entities into the current packet for Add
    	raises InterfaceError;
    --           Error if on of the items of <list> is not from the Model, or
    --           if no AddPacket was yet called

    NbPackets (me) returns Integer;
    ---Purpose : Returns the count of non-empty packets

    NbEntities (me; numpack : Integer) returns Integer;
    ---Purpose : Returns the count of entities in a Packet given its rank, or 0

    Entities (me; numpack : Integer) returns EntityIterator;
    ---Purpose : Returns the content of a Packet given its rank
    --           Null Handle if <numpack> is out of range

    HighestDuplicationCount (me) returns Integer;
    ---Purpose : Returns the highest number of packets which know a same entity
    --           For no duplication, should be one

    NbDuplicated (me; count : Integer; andmore : Boolean) returns Integer;
    ---Purpose : Returns the count of entities duplicated :
    --           <count> times, if <andmore> is False, or
    --           <count> or more times, if <andmore> is True
    --           See Duplicated for more details

    Duplicated (me; count : Integer; andmore : Boolean) returns EntityIterator;
    ---Purpose : Returns a list of entities duplicated :
    --           <count> times, if <andmore> is False, or
    --           <count> or more times, if <andmore> is True
    --           Hence, count=2 & andmore=True gives all duplicated entities
    --           count=1 gives non-duplicated entities (in only one packet)
    --           count=0 gives remaining entities (in no packet at all)

fields

    themodel : InterfaceModel;
    thedupls : Array1OfInteger;
    thepacks : IntList;
    theflags : Array1OfInteger;   -- for only once par packet !
    thelast  : Integer;
    thebegin : Boolean;
    thename  : AsciiString;

end PacketList;
