-- Created on: 1992-11-24
-- Created by: Didier PIFFAULT
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class BoundSortBox from Bnd 

	---Purpose: A tool to compare a bounding box or a plane with a set of
    	-- bounding boxes. It sorts the set of bounding boxes to give
    	-- the list of boxes which intersect the element being compared.
    	-- The boxes being sorted generally bound a set of shapes,
    	-- while the box being compared bounds a shape to be
    	-- compared. The resulting list of intersecting boxes therefore
    	-- gives the list of items which potentially intersect the shape to be compared.


uses    Integer from Standard,
    	Real from Standard,
    	ListOfInteger from TColStd,
	Pln from gp,
    	Box from Bnd,
    	HArray1OfBox from Bnd,
	DataMapOfIntegerInteger from TColStd


raises  NullValue from Standard, MultiplyDefined from Standard


is      Create      returns BoundSortBox from Bnd;
	---Purpose: Constructs an empty comparison algorithm for bounding boxes.
    	-- The bounding boxes are then defined using the Initialize function.


    	Initialize (me : in out;
    	    	    CompleteBox : Box from Bnd; 
    	    	    SetOfBox    : HArray1OfBox from Bnd)
		    is static;
	---Purpose: Initializes this comparison algorithm with
    	-- -   the set of bounding boxes SetOfBox.

    	Initialize (me : in out;
    	    	    SetOfBox    : HArray1OfBox from Bnd)
		    is static;
	---Purpose: Initializes this comparison algorithm with
    	-- -   the set of bounding boxes SetOfBox, where
    	--   CompleteBox is given as the global bounding box of SetOfBox.


    	SortBoxes  (me : in out)
		    raises NullValue from Standard is static private;
	---Purpose: Prepares  BoundSortBox and  sorts   the  boxes of
	--          <SetOfBox> .



    	Initialize (me : in out;
    	    	    CompleteBox : Box from Bnd; 
    	    	    nbComponents : Integer from Standard)
		    raises NullValue from Standard is static;
	---Purpose: Initializes this comparison algorithm, giving it only
    	-- -   the maximum number nbComponents
    	-- of the bounding boxes to be managed. Use the Add
    	-- function to define the array of bounding boxes to be sorted by this algorithm.


    	Add        (me          : in out;
    	    	    theBox      : Box from Bnd;
    	    	    boxIndex    : Integer from Standard)
		    raises MultiplyDefined from Standard is static;
	---Purpose: Adds the bounding box theBox at position boxIndex in
    	-- the array of boxes to be sorted by this comparison algorithm.
    	-- This function is used only in conjunction with the third
    	-- syntax described in the synopsis of Initialize.
	--
    	-- Exceptions:
	--
    	-- - Standard_OutOfRange if boxIndex is not in the
    	--   range [ 1,nbComponents ] where
    	--   nbComponents is the maximum number of bounding
    	--   boxes declared for this comparison algorithm at
    	--   initialization.
	--
    	-- - Standard_MultiplyDefined if a box already exists at
    	--   position boxIndex in the array of boxes to be sorted by
    	--   this comparison algorithm.
  

    	Compare    (me : in out;
    	    	    theBox      : Box from Bnd)
	    	    returns ListOfInteger from TColStd
	---Purpose: Compares the bounding box theBox, 
    	-- with the set of bounding boxes to be sorted by this
    	-- comparison algorithm, and returns the list of intersecting
    	-- bounding boxes as a list of indexes on the array of
    	-- bounding boxes used by this algorithm.                  
    		    ---C++: return const &
   raises NullValue from Standard is static;

    	Compare    (me : in out;
    	    	    P : Pln from gp)
	    	    returns ListOfInteger from TColStd
	---Purpose: Compares the plane P
        -- with the set of bounding boxes to be sorted by this
    	-- comparison algorithm, and returns the list of intersecting
    	-- bounding boxes as a list of indexes on the array of
    	-- bounding boxes used by this algorithm.
		   ---C++: return const &
   raises NullValue from Standard is static;

    	Dump       (me) is static;

    	Destroy(me: in out)
	---C++: alias ~
	    is static;

fields  myBox           : Box from Bnd;
    	myBndComponents : HArray1OfBox from Bnd;
    	Xmin            : Real from Standard;
    	Ymin            : Real from Standard;
    	Zmin            : Real from Standard;
	deltaX          : Real from Standard;
    	deltaY          : Real from Standard;
    	deltaZ          : Real from Standard;
    	discrX          : Integer from Standard;
    	discrY          : Integer from Standard;
    	discrZ          : Integer from Standard;
    	theFound        : Integer from Standard;
	Crible          : DataMapOfIntegerInteger from TColStd;
	lastResult      : ListOfInteger from TColStd;
    	TabBits         : Address from Standard;
end BoundSortBox;
