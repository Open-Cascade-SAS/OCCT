-- Created on: 1992-06-22
-- Created by: Gilles DEBARBOUILLE
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



private class UnitSentence from Units

	---Purpose: This   class describes   all    the  facilities to
	--          manipulate and compute units contained in a string
	--          expression.

inherits

    Sentence from Units

uses

    QuantitiesSequence from Units

--raises

is

    Create(astring : CString)
    
    ---Level: Internal 
    
    ---Purpose: Creates   and   returns a   UnitSentence.   The string
    --          <astring> describes in natural  language the  unit  or
    --          the composed unit to be analysed.
    
    returns UnitSentence from Units;
    
    Create(astring : CString ; aquantitiessequence : QuantitiesSequence from Units)
    
    ---Level: Internal 
    
    ---Purpose: Creates  and returns    a  UnitSentence.  The   string
    --          <astring> describes in natural language the unit to be
    --          analysed.   The    sequence     of physical quantities
    --          <asequenceofquantities>   describes    the   available
    --          dictionary of units you want to use.
    
    returns UnitSentence from Units;
    
    Analyse(me : in out)
    
    ---Level: Internal 
    
    ---Purpose: Analyzes   the sequence  of   tokens  created  by  the
    --          constructor to  find  the true significance   of  each
    --          token.
    
    is static;
    
    SetUnits(me : in out ; aquantitiessequence : QuantitiesSequence from Units)
    
    ---Level: Internal 
    
    ---Purpose: For each token which  represents a unit, finds  in the
    --          sequence    of    physical   quantities      all   the
    --          characteristics of the unit found.
    
    is static;

--fields

end UnitSentence;
