-- Created on: 1992-04-06
-- Created by: Christian CAILLET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DefSwitch  from IGESData  inherits Storable

    ---Purpose : description of a directory componant which can be either
    --           undefined (let Void), defined as a Reference to an entity,
    --           or as a Rank, integer value adressing a builtin table
    --           The entity reference is not included here, only reference
    --           status is kept (because entity type must be adapted)

uses Integer, DefType

is

    Create returns DefSwitch;
    ---Purpose : creates a DefSwitch as Void

    SetVoid (me : in out)  is static;
    ---Purpose : sets DefSwitch to "Void" status (in file : Integer = 0)

    SetReference (me : in out)  is static;
    ---Purpose : sets DefSwitch to "Reference" Status (in file : Integer < 0)

    SetRank (me : in out; val : Integer)  is static;
    ---Purpose : sets DefSwitch to "Rank" with a Value (in file : Integer > 0)

    DefType (me) returns DefType  is static;
    ---Purpose : returns DefType status (Void,Reference,Rank)

    Value (me) returns Integer  is static;
    ---Purpose : returns Value as Integer (sensefull for a Rank)

fields

    theval : Integer;

end DefSwitch;
