-- File:        BezierCurveAndRationalBSplineCurve.cdl
-- Created:     Mon Dec  4 12:02:33 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWBezierCurveAndRationalBSplineCurve from RWStepGeom

	---Purpose : Read & Write Module for BezierCurveAndRationalBSplineCurve

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     BezierCurveAndRationalBSplineCurve from StepGeom,
     EntityIterator from Interface

is

	Create returns RWBezierCurveAndRationalBSplineCurve;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable BezierCurveAndRationalBSplineCurve from StepGeom);

	WriteStep (me; SW : in out StepWriter; ent : BezierCurveAndRationalBSplineCurve from StepGeom);

	Share(me; ent : BezierCurveAndRationalBSplineCurve from StepGeom; iter : in out EntityIterator);

end RWBezierCurveAndRationalBSplineCurve;
