-- File:        BezierCurve.cdl
-- Created:     Mon Dec  4 12:02:23 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWBezierCurve from RWStepGeom

	---Purpose : Read & Write Module for BezierCurve

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     BezierCurve from StepGeom,
     EntityIterator from Interface

is

	Create returns RWBezierCurve;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable BezierCurve from StepGeom);

	WriteStep (me; SW : in out StepWriter; ent : BezierCurve from StepGeom);

	Share(me; ent : BezierCurve from StepGeom; iter : in out EntityIterator);

end RWBezierCurve;
