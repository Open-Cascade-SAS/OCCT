-- Created on: 1995-04-25
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package LocOpe

        ---Purpose: Provides  tools to implement local     topological
        --          operations on a shape.

uses MMgt,
     StdFail,
     TCollection,
     TColStd,
     gp, 
     Geom,
     TColGeom,
     TColgp,

     TopAbs,
     TopoDS,
     TopExp,
     TopTools,
     BRepFill,
     BRepSweep, 
     TopOpeBRepDS
--     TopOpeBRepBuild

is 

    class SplitShape;

    deferred class ProjectedWires;      -- inherits TShared from MMgt
    
    class WiresOnShape;                 -- inherits ProjectedWires from LocOpe


    class Spliter;

    class Generator;

    deferred class GeneratedShape;      -- inherits TShared from MMgt
    
    class GluedShape;                   -- inherits GeneratedShape from LocOpe
    class Prism;
    class Revol;

    class Pipe;

    class DPrism;

    class LinearForm;

    class RevolutionForm;

    class Gluer;

    class FindEdges;

    class FindEdgesInFace;

    class DataMapOfShapePnt instantiates DataMap from TCollection
            (Shape          from TopoDS,
         Pnt            from gp,
         ShapeMapHasher from TopTools);

    class PntFace;
    
    class CurveShapeIntersector;
    
    class CSIntersector;
    

    class BuildShape;

    class SplitDrafts;


    class SequenceOfPntFace instantiates Sequence from TCollection
            (PntFace from LocOpe);

    class SequenceOfLin instantiates Sequence from TCollection
            (Lin from gp);

    class SequenceOfCirc instantiates Sequence from TCollection
            (Circ from gp);

    private class HBuilder;    -- inherits HBuilder from TopOpeBRepBuild

    private class BuildWires;   -- used in LocOpe_Spliter

    enumeration Operation is
            FUSE,
        CUT,
        INVALID
    end Operation;


    Closed(W: Wire from TopoDS; OnF: Face from TopoDS)
        ---Purpose: Returns Standard_True  when the wire <W> is closed
        --          on the face <OnF>.
            returns Boolean from Standard;
    

    Closed(E: Edge from TopoDS; OnF: Face from TopoDS)
        ---Purpose: Returns Standard_True  when the edge <E> is closed
        --          on the face <OnF>.
            returns Boolean from Standard;

    TgtFaces(E : Edge from TopoDS; 
                 F1: Face from TopoDS;
                 F2: Face from TopoDS)
        ---Purpose: Returns Standard_True  when the faces are tangent
            returns Boolean from Standard;


    
--    IsInside(F1: Face from TopoDS; F2: Face from TopoDS)
--         ---Purpose: Returns Standard_True when  the face F1 is in  the
--         --          F2 .
--            returns Boolean from Standard;
   

    SampleEdges(S : Shape from TopoDS;
                    Pt: in out SequenceOfPnt from TColgp);


end LocOpe;





