-- Created on: 1994-06-01
-- Created by: Christian CAILLET
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class SelectBypassGroup  from IGESSelect  inherits SelectExplore

    ---Purpose : Selects a list built as follows :
    --           Groups are entities type 402, forms 1,7,14,15 (Group,
    --           Ordered or not, "WithoutBackPointer" or not)
    --           
    --           Entities which are not GROUP are taken as such
    --           For Groups, their list of Elements is explore
    --           Hence, level 0 (D) recursively explores a Group if some of
    --           its Elements are Groups. level 1 explores just at first level

uses AsciiString from TCollection, Transient, EntityIterator, Graph

raises InterfaceError

is

    Create (level : Integer = 0) returns mutable SelectBypassGroup;
    ---Purpose : Creates a SelectBypassGroup, by default all level
    --           (level = 1 explores at first level)

    Explore (me; level : Integer; ent : Transient; G : Graph;
    	     explored : in out EntityIterator)
    	returns Boolean;
    ---Purpose : Explores an entity : for a Group, gives its elements
    --           Else, takes the entity itself


    ExploreLabel (me) returns AsciiString from TCollection;
    ---Purpose : Returns a text defining the criterium : "Content of Group"

end SelectBypassGroup;
