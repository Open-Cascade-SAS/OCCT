-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SolidReplica from StepShape 

inherits SolidModel from StepShape 

uses

	CartesianTransformationOperator3d from StepGeom,
	HAsciiString from TCollection
is

	Create returns mutable SolidReplica;
	---Purpose: Returns a SolidReplica


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aParentSolid : mutable SolidModel from StepShape;
	      aTransformation : mutable CartesianTransformationOperator3d from StepGeom) is virtual;

	-- Specific Methods for Field Data Access --

	SetParentSolid(me : mutable; aParentSolid : mutable SolidModel);
	ParentSolid (me) returns mutable SolidModel;
	SetTransformation(me : mutable; aTransformation : mutable CartesianTransformationOperator3d);
	Transformation (me) returns mutable CartesianTransformationOperator3d;

fields

	parentSolid : SolidModel from StepShape;
	transformation : CartesianTransformationOperator3d from StepGeom;

end SolidReplica;
