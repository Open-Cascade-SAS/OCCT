-- File:	MDataXtd_GeometryStorageDriver.cdl
-- Created:	Wed Nov 19 15:57:14 1997
-- Author:	Denis PASCAL
--		<dp@dingox.paris1.matra-dtv.fr>
-- modified     Sergey Zaritchny
---Copyright:	 Matra Datavision 1997


class GeometryStorageDriver from MDataXtd inherits ASDriver from MDF

	---Purpose: 

uses SRelocationTable from MDF,
     Attribute        from TDF,
     Attribute        from PDF, 
     MessageDriver    from CDM


is

    Create(theMessageDriver : MessageDriver from CDM) 
    returns mutable GeometryStorageDriver from MDataXtd;


    VersionNumber(me) returns Integer from Standard;
	---Purpose: Returns the version number from which the driver
	--          is available: 0.

    SourceType(me) returns Type from Standard;
	---Purpose: Returns the type: Integer from TDataStd.

    NewEmpty (me) returns mutable Attribute from PDF;


    Paste(me;
    	  Source     :         Attribute from TDF;
    	  Target     : mutable Attribute from PDF;
    	  RelocTable : SRelocationTable from MDF);


end GeometryStorageDriver;

