
-- File:	BinMXCAFDoc_LocationDriver.cdl
-- Created:	Tue May 17 14:42:38 2005
-- Author:	Eugeny NAPALKOV <eugeny.napalkov@opencascade.com>
-- Copyright:	Open CasCade S.A. 2005

class LocationDriver from BinMXCAFDoc inherits ADriver from BinMDF

uses
    MessageDriver    from CDM,
    SRelocationTable from BinObjMgt,
    RRelocationTable from BinObjMgt,
    Persistent       from BinObjMgt,
    Location         from TopLoc,
    Attribute        from TDF,
    LocationSetPtr   from BinTools
is
    Create (theMsgDriver:MessageDriver from CDM)
    returns mutable LocationDriver from BinMXCAFDoc;

    NewEmpty (me)  returns mutable Attribute from TDF
    is redefined;

    Paste(me; theSource     : Persistent from BinObjMgt;
              theTarget     : mutable Attribute from TDF;
              theRelocTable : out RRelocationTable from BinObjMgt)
    returns Boolean from Standard is redefined;

    Paste(me; theSource     : Attribute from TDF;
              theTarget     : in out Persistent from BinObjMgt;
              theRelocTable : out SRelocationTable from BinObjMgt)
    is redefined;
    
    Translate(me; theSource     : Persistent from BinObjMgt;
	               theLoc        : in out Location from TopLoc;
         	       theMap        : out RRelocationTable from BinObjMgt)
    returns Boolean from Standard;
    
    Translate(me; theLoc        : Location from TopLoc;
    	    	       theTarget     : in out Persistent from BinObjMgt;
		       theMap        : out SRelocationTable from BinObjMgt);
    ---Purpose: Translate transient location to storable
    
    SetSharedLocations(me: mutable;
                       theLocations:  in LocationSetPtr  from BinTools);
    ---C++: inline
    
fields
    myLocations : LocationSetPtr   from BinTools;
end;
