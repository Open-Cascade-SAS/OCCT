-- Created on: 1993-06-07
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class ArcFunction from IntPatch

inherits FunctionWithDerivative from math

uses
     HCurve2d      from Adaptor2d,
     HSurface      from Adaptor3d,
     Pnt           from gp,
     SequenceOfPnt from TColgp,
     Quadric       from IntSurf

is

    Create
    
    	returns ArcFunction from IntPatch;


    SetQuadric(me: in out; Q: Quadric from IntSurf)
    
	---C++: inline
    	is static;


    Set(me: in out; A: HCurve2d from Adaptor2d)
    
	---C++: inline
    	is static;


    Set(me: in out; S: HSurface from Adaptor3d)
    
	---C++: inline
    	is static;


    Value(me: in out; X: Real from Standard; F: out Real from Standard)
    
    	returns Boolean from Standard;
    

    Derivative(me: in out; X: Real from Standard; D: out Real from Standard)
    
    	returns Boolean from Standard;
    

    Values(me: in out; X: Real from Standard; F,D: out Real from Standard)
    
    	returns Boolean from Standard;
    

    NbSamples(me)
    
    	returns Integer from Standard
	is static;


    GetStateNumber(me: in out)

    	returns Integer from Standard
    	is redefined;
	
	
    Valpoint(me; Index: Integer from Standard)
    
    	returns Pnt from gp
	---C++: return const&
	---C++: inline
	is static;
    
    Quadric(me) 
    	returns Quadric from IntSurf
	---C++: return const&
	---C++: inline
	is static;
       
    Arc(me)
   	returns HCurve2d from Adaptor2d
	---C++: return const&
	---C++: inline
	is static;
       
    Surface(me)
   	returns HSurface from Adaptor3d
	---C++: return const&
	---C++: inline
	is static;
	    
fields

    myArc  : HCurve2d      from Adaptor2d;
    mySurf : HSurface      from Adaptor3d;
    myQuad : Quadric       from IntSurf;
    ptsol  : Pnt           from gp;
    seqpt  : SequenceOfPnt from TColgp;

end ArcFunction;
