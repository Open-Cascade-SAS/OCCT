-- Created on: 2009-06-17
-- Created by: Sergey ZARITCHNY <sergey.zaritchny@opencascade.com>
-- Copyright (c) 2009-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class RevolutionDriver from DNaming inherits Driver from TFunction

	---Purpose: 
uses
     Label       from TDF, 
     Logbook     from TFunction,
     Function    from TFunction,
     ExtendedString from TCollection,
     MakeRevol   from BRepPrimAPI, 
     Shape       from TopoDS
is
    Create returns mutable RevolutionDriver from DNaming;
    ---Purpose: Constructor

    ---Purpose: validation
    --          ==========

    Validate(me; theLog : in out Logbook from TFunction)
    is redefined;
    ---Purpose: Validates labels of a function in <log>.
    --          In regeneration mode this method must be called (by the
    --          solver) even if the function is not executed, to build
    --          the valid label scope.

    ---Purpose: execution of function
    --          ======================

    MustExecute (me; theLog : Logbook from TFunction)
    ---Purpose: Analyse in <log> if the loaded function must be executed
    --          (i.e.arguments are modified) or not.
    --          If the Function label itself is modified, the function must
    --          be executed.
    returns Boolean from Standard
    is redefined;

    Execute (me; theLog : in out Logbook from TFunction)
    ---Purpose: Execute the function and push in <log> the impacted
    --          labels (see method SetImpacted).
    returns Integer from Standard
    is redefined;
 
    LoadNamingDS(me; theResultLabel : Label from TDF; mkRevol : in out MakeRevol from BRepPrimAPI; 
    	    	     Basis : Shape from TopoDS; Context : Shape from TopoDS)  
    is private;      


end RevolutionDriver;
