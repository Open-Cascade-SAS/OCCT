-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Face from StepShape 

inherits TopologicalRepresentationItem from StepShape 

uses

	HArray1OfFaceBound from StepShape, 
	FaceBound from StepShape, 
	HAsciiString from TCollection
is

	Create returns Face;
	---Purpose: Returns a Face


	Init (me : mutable;
	      aName : HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      aName : HAsciiString from TCollection;
	      aBounds : HArray1OfFaceBound from StepShape) is virtual;

	-- Specific Methods for Field Data Access --

	SetBounds(me : mutable; aBounds : HArray1OfFaceBound)
    	is virtual;
	Bounds (me) returns HArray1OfFaceBound
    	is virtual;
	BoundsValue (me; num : Integer) returns FaceBound
    	is virtual;
	NbBounds (me) returns Integer
    	is virtual;

fields

	bounds : HArray1OfFaceBound from StepShape;

end Face;
