-- File:	Geom2dGcc.cdl
-- Created:	Mon Jun 29 14:55:26 1992
-- Author:	Remi GILET
--		<reg@sdsun2>
---Copyright:	 Matra Datavision 1992


package Geom2dGcc 

    	--- Purpose: The Geom2dGcc package describes qualified 2D
    	-- curves used in the construction of constrained geometric
    	-- objects by an algorithm provided by the Geom2dGcc package.
    	-- A qualified 2D curve is a curve with a qualifier which
    	-- specifies whether the solution of a construction
    	-- algorithm using the qualified curve (as an argument):
    	-- -   encloses the curve, or
    	-- -   is enclosed by the curve, or
    	-- -   is built so that both the curve and this solution are external to one another, or
    	-- -   is undefined (all solutions apply).
    	-- These package methods provide simpler functions to construct a qualified curve.
    	-- Note: the interior of a curve is defined as the left-hand
    	-- side of the curve in relation to its orientation.


uses GccEnt,
     GccGeo,
     GccAna,
     GccIter,
     StdFail,
     Geom2dInt,
     Geom2d,
     TColStd,
     TopAbs,	
     Standard,
     Geom2dAdaptor,
     Extrema,
     Adaptor3d,
     Adaptor2d,
     TColgp,
     gp

is

class CurveTool;

class QualifiedCurve;

class Circ2d3Tan;

class Circ2d2TanRad;

class Circ2d2TanOn;

class Circ2dTanOnRad;

class Circ2dTanCen;

class Lin2d2Tan;

class Lin2dTanObl;

class MyQCurve instantiates QualifiedCurv from GccEnt
    	    (Curve  from Geom2dAdaptor);

class MyCurveTool instantiates CurvePGTool from GccGeo
    	    (Curve       from Geom2dAdaptor,
    	     CurveTool   from Geom2dGcc    ,
    	     OffsetCurve from Adaptor3d);
	    
class MyCirc2d2TanOn instantiates Circ2d2TanOn from GccGeo
    	    (Curve                          from Geom2dAdaptor,
	     CurveTool                      from Geom2dGcc,
    	     MyQCurve                       from Geom2dGcc,
             OffsetCurve                    from Adaptor3d,
	     HCurve                         from Geom2dAdaptor,
	     MyCurveTool                    from Geom2dGcc,
	     TheIntConicCurveOfGInter from Geom2dInt);
	     
class MyCirc2d2TanRad instantiates Circ2d2TanRad from GccGeo
    	    (Curve                           from Geom2dAdaptor ,
	     CurveTool                       from Geom2dGcc,
    	     MyQCurve                        from Geom2dGcc,
             OffsetCurve                     from Adaptor3d, 
	     HCurve                         from Geom2dAdaptor,	     
	     MyCurveTool                     from Geom2dGcc,
	     TheIntConicCurveOfGInter  from Geom2dInt,
	     GInter                    from Geom2dInt);

class MyCirc2dTanOnRad instantiates Circ2dTanOnRad from GccGeo
    	    (Curve                           from Geom2dAdaptor ,
	     CurveTool                       from Geom2dGcc,
    	     MyQCurve                        from Geom2dGcc,
	     OffsetCurve                     from Adaptor3d,
	     HCurve                         from Geom2dAdaptor,	     
	     MyCurveTool                     from Geom2dGcc,
	     TheIntConicCurveOfGInter  from Geom2dInt,
	     GInter                    from Geom2dInt);

class MyC2d3Tan instantiates Circ2d3Tan from GccIter	     
    	    (Curve          from Geom2dAdaptor,
	     CurveTool      from Geom2dGcc,
	     MyQCurve       from Geom2dGcc);
	     
class MyCirc2dTanCen instantiates Circ2dTanCen from GccGeo	     
    	    (Curve          from Geom2dAdaptor,
	     CurveTool      from Geom2dGcc,
	     ExtPC2d          from Extrema,
             MyQCurve       from Geom2dGcc);
	     
class MyC2d2TanOn instantiates Circ2d2TanOn from GccIter	     
    	    (Curve          from Geom2dAdaptor,
	     CurveTool      from Geom2dGcc,
	     MyQCurve       from Geom2dGcc);

class MyL2dTanObl instantiates Lin2dTanObl from GccIter	     
    	    (Curve          from Geom2dAdaptor,
	     CurveTool      from Geom2dGcc,
	     MyQCurve       from Geom2dGcc);
	     
class MyL2d2Tan instantiates Lin2d2Tan from GccIter	     
    	    (Curve          from Geom2dAdaptor,
	     CurveTool      from Geom2dGcc,
	     MyQCurve       from Geom2dGcc);

Unqualified(Obj : Curve from Geom2dAdaptor) returns QualifiedCurve;
    	---Purpose: Constructs such a qualified curve that the relative
    	-- position of the solution computed by a construction
    	-- algorithm using the qualified curve to the circle or line is
    	-- not qualified, i.e. all solutions apply.
    	-- Warning
    	-- Obj is an adapted curve, i.e. an object which is an interface between:
    	-- -   the services provided by a 2D curve from the package Geom2d,
    	-- -   and those required on the curve by a computation algorithm.
    	--  The adapted curve is created in the following way:
    	-- Handle(Geom2d_Curve) mycurve = ...
    	-- ;
    	-- Geom2dAdaptor_Curve Obj ( mycurve )
    	-- ;
    	-- The qualified curve is then constructed with this object:
    	-- Geom2dGcc_QualifiedCurve
    	-- myQCurve = Geom2dGcc::Unqualified(Obj);
    
Enclosing(Obj : Curve from Geom2dAdaptor) returns QualifiedCurve;
    	---Purpose: Constructs such a qualified curve that the solution
    	-- computed by a construction algorithm using the qualified
    	-- curve encloses the curve.
    	-- Warning
    	-- Obj is an adapted curve, i.e. an object which is an interface between:
    	-- -   the services provided by a 2D curve from the package Geom2d,
    	-- -   and those required on the curve by a computation algorithm.
    	-- The adapted curve is created in the following way:
    	-- Handle(Geom2d_Curve) mycurve = ...
    	-- ;
    	-- Geom2dAdaptor_Curve Obj ( mycurve )
    	-- ;
    	-- The qualified curve is then constructed with this object:
    	-- Geom2dGcc_QualifiedCurve
    	--              myQCurve = Geom2dGcc::Enclosing(Obj);
  
Enclosed(Obj : Curve from Geom2dAdaptor) returns QualifiedCurve;
    	---Purpose: Constructs such a qualified curve that the solution
    	-- computed by a construction algorithm using the qualified
    	-- curve is enclosed by the curve.
    	-- Warning
    	-- Obj is an adapted curve, i.e. an object which is an interface between:
    	-- -   the services provided by a 2D curve from the package Geom2d,
    	-- -   and those required on the curve by a computation algorithm.
    	-- The adapted curve is created in the following way:
    	-- Handle(Geom2d_Curve) mycurve = ...
    	-- ;
    	-- Geom2dAdaptor_Curve Obj ( mycurve )
    	-- ;
    	-- The qualified curve is then constructed with this object:
    	-- Geom2dGcc_QualifiedCurve
    	--              myQCurve = Geom2dGcc::Enclosed(Obj);
    
Outside(Obj : Curve from Geom2dAdaptor) returns QualifiedCurve;
    	---Purpose: Constructs such a qualified curve that the solution
    	-- computed by a construction algorithm using the qualified
    	-- curve and the curve are external to one another.
    	-- Warning
    	-- Obj is an adapted curve, i.e. an object which is an interface between:
    	-- -   the services provided by a 2D curve from the package Geom2d,
    	-- -   and those required on the curve by a computation algorithm.
    	-- The adapted curve is created in the following way:
    	-- Handle(Geom2d_Curve) mycurve = ...
    	-- ;
    	-- Geom2dAdaptor_Curve Obj ( mycurve )
    	-- ;
    	-- The qualified curve is then constructed with this object:
    	-- Geom2dGcc_QualifiedCurve
    	--              myQCurve = Geom2dGcc::Outside(Obj);
	     
end Geom2dGcc;
