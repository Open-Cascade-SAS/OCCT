-- Created on: 1992-12-15
-- Created by: Jean Louis FRENKEL
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class Root from Prs3d

    	---Purpose: A root class for the standard presentation algorithms
    	-- of the StdPrs package.
    	--          
uses
    Presentation from Prs3d,
    Structure from Graphic3d,
    Group from Graphic3d

is
    CurrentGroup(myclass; Prs3d: Presentation from Prs3d) returns Group from Graphic3d;
    	---Purpose: Returns the current group of primititves inside graphic
    	-- objects in the display.
    	-- A group also contains the attributes whose ranges are
    	-- limited to the primitives in it. 
    
    NewGroup (myclass; Prs3d: Presentation from Prs3d ) returns Group from Graphic3d ;
    	---Purpose: Returns the new group of primitives inside graphic
    	-- objects in the display.
    	-- A group also contains the attributes whose ranges are limited to the primitives in it.
    
end Root from Prs3d;
