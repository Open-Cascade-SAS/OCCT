-- Created on: 1999-05-06
-- Created by: Pavel DURANDIN
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ShapeDivideAngle from ShapeUpgrade inherits ShapeDivide from ShapeUpgrade

	---Purpose: Splits all surfaces of revolution, cylindrical, toroidal, 
    	--          conical, spherical surfaces in the given shape so that 
	--          each resulting segment covers not more than defined number 
	--          of degrees. 

uses
    
    Shape from TopoDS

is
    Create (MaxAngle: Real) returns ShapeDivideAngle from ShapeUpgrade;
    	---Purpose: Empty constructor.
    
    Create (MaxAngle: Real; S: Shape from TopoDS)
    returns ShapeDivideAngle from ShapeUpgrade;
    	---Purpose: Initialize by a Shape.

    InitTool (me: in out; MaxAngle: Real);
     	---Purpose: Resets tool for splitting face with given angle

    SetMaxAngle (me: in out; MaxAngle: Real);
    	---Purpose: Set maximal angle (calls InitTool)
    
    MaxAngle (me) returns Real;
    	---Purpose: Returns maximal angle 
    
end ShapeDivideAngle;
