-- Created on: 1993-03-03
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class Location from PTopLoc inherits Storable

	---Purpose: A Storable  composed local coordinate system. Made
	--          with local   coordinate systems raised   to  power
	--          elevation.
	--          
	--          A Location is either :
	--          
	--          * The Identity.
	--          
	--          * The product  of a Datum3D raised  to a power and
	--          an other Location called the next Location.

uses
    Datum3D      from PTopLoc,
    ItemLocation from PTopLoc

raises
    NoSuchObject from Standard

is
    Create returns Location from PTopLoc;
	---Purpose: Creates an Identity Location.
	---Level: Internal 
	
    Create(D : Datum3D from PTopLoc; 
    	   P : Integer from Standard;
	   N : Location from PTopLoc) 
    returns Location from  PTopLoc;
	---Purpose: Creates a location being the product.
	--          N * D ^ P
	---Level: Internal 
    
    IsIdentity(me) returns Boolean from Standard
	---Purpose: True when the location is an identity.
	---Level: Internal 
    is static;
    
    Datum3D(me) returns Datum3D from PTopLoc
	---Purpose: Returns the first Datum. An error is raised if the
	--          location is an identity.
	---Level: Internal 
    raises NoSuchObject from Standard
    is static;

    Power(me)   returns Integer from Standard
	---Purpose: Returns the power elevation of the first datum. An
	--          error is raised if the location is an identity.
	---Level: Internal 
    raises NoSuchObject from Standard
    is static;
    
    Next(me)    returns Location from PTopLoc
	---Purpose: Returns next Location. An error is raised if the
	--          location is an identity.
	---Level: Internal 
    raises NoSuchObject from Standard
    is static;
    
fields
    myData : ItemLocation from PTopLoc;

end Location;
