-- Created on: 1992-11-18
-- Created by: Christian CAILLET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

generic class SelectList  from IFSelect (Entity as Transient)
    	inherits SelectInList


    ---Purpose : A SelectList kind Selection selects a part of an Entity, as
    --           well as this Entity can be described as an ordered List.
    --           That is to say, it must have two methods :
    --
    --             NbEntities (me) returns Integer;
    --             Entity (me; num : Integer) returns Transient;
    --           
    --           For each class of Entity for which we want to define a
    --           SelectList, we will instanciate this class with the
    --           desired class of Entity as definition parameter : the deferred
    --           methods NbEntities and ListedEntity are now defined to call
    --           the required methods from <Entity>
    --
    --           SelectList works as SelectInList, beeing a sub-class of it

uses AsciiString from TCollection, Transient, EntityIterator, IntParam

raises OutOfRange

is

    Create returns mutable SelectList;
    ---Purpose : Creates a SelectList (with no limit);

    KeepInputEntity (me; iter : in out EntityIterator);
    ---Purpose : Keeps Input Entity, as having required type <Entity>

    NbItems (me; ent : Transient) returns Integer;
    ---Purpose : Returns count of Entities in the list in the Entity <ent>
    --           by calling method NbEntity from parameter class Entity

    ListedEntity (me; num : Integer; ent : Transient)
    	returns Transient  raises OutOfRange;
    ---Purpose : Returns an Entity of the list in the Entity <ent>, by calling
    --           method Entity from parameter class Entity
    --           Error if <ent> has not required type, or if <num> is not in
    --           the right range (1,NbEntities),

    ListLabel (me) returns AsciiString from TCollection;
    ---Purpose : Returns the specific label for the list
    --           then, following cases :
    --           " From .. Until .." or "From .." or "Until .." or "Rank no .."
    --  Warning : it is not possible to give a character constant to instantiate
    --           a generic class, thus "List From Entity" is not adapted :
    --           redefine Label if judged necessary

end SelectList;
