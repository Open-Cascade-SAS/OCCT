-- File:        DocumentUsageConstraint.cdl
-- Created:     Mon Dec  4 12:02:29 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWDocumentUsageConstraint from RWStepBasic

	---Purpose : Read & Write Module for DocumentUsageConstraint

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     DocumentUsageConstraint from StepBasic,
     EntityIterator from Interface

is

	Create returns RWDocumentUsageConstraint;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable DocumentUsageConstraint from StepBasic);

	WriteStep (me; SW : in out StepWriter; ent : DocumentUsageConstraint from StepBasic);

	Share(me; ent : DocumentUsageConstraint from StepBasic; iter : in out EntityIterator);

end RWDocumentUsageConstraint;
