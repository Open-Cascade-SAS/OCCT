-- Created on: 1992-07-20
-- Created by: Arnaud BOUZY
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



deferred class Generator from ExprIntrp inherits TShared from MMgt

	---Purpose: Implements general services for interpretation of 
	--          expressions.

uses NamedExpression from Expr,
    NamedFunction from Expr,
    SequenceOfNamedFunction from ExprIntrp,
    SequenceOfNamedExpression from ExprIntrp,
    AsciiString from TCollection

is

    Initialize;
    
    Use(me : mutable; func : NamedFunction)
    ---Level: Internal 
    is static;

    Use(me : mutable; named : NamedExpression)
    ---Level: Internal 
    is static;
        
    GetNamed(me)
    returns SequenceOfNamedExpression
    ---C++: return const &
    ---Level: Internal 
    is static;
    
    GetFunctions(me)
    returns SequenceOfNamedFunction
    ---C++: return const &
    ---Level: Internal 
    is static;

    GetNamed(me; name : AsciiString)
    ---Purpose: Returns NamedExpression with name <name> already 
    --          interpreted if it exists. Returns a null handle if 
    --          not. 
    ---Level: Advanced
    returns any NamedExpression
    is static;
    
    GetFunction(me; name : AsciiString)
    ---Purpose: Returns NamedFunction with name <name> already 
    --          interpreted if it exists. Returns a null handle if 
    --          not.
    ---Level: Advanced 
    returns any NamedFunction
    is static;
    
fields

    myFunctions : SequenceOfNamedFunction;
    myNamed : SequenceOfNamedExpression;
    
end Generator;
