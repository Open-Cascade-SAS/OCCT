-- Created on: 2005-05-17
-- Created by: Eugeny NAPALKOV <eugeny.napalkov@opencascade.com>
-- Copyright (c) 2005-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class LocationDriver from BinMXCAFDoc inherits ADriver from BinMDF

uses
    MessageDriver    from CDM,
    SRelocationTable from BinObjMgt,
    RRelocationTable from BinObjMgt,
    Persistent       from BinObjMgt,
    Location         from TopLoc,
    Attribute        from TDF,
    LocationSetPtr   from BinTools
is
    Create (theMsgDriver:MessageDriver from CDM)
    returns mutable LocationDriver from BinMXCAFDoc;

    NewEmpty (me)  returns mutable Attribute from TDF
    is redefined;

    Paste(me; theSource     : Persistent from BinObjMgt;
              theTarget     : mutable Attribute from TDF;
              theRelocTable : out RRelocationTable from BinObjMgt)
    returns Boolean from Standard is redefined;

    Paste(me; theSource     : Attribute from TDF;
              theTarget     : in out Persistent from BinObjMgt;
              theRelocTable : out SRelocationTable from BinObjMgt)
    is redefined;
    
    Translate(me; theSource     : Persistent from BinObjMgt;
	               theLoc        : in out Location from TopLoc;
         	       theMap        : out RRelocationTable from BinObjMgt)
    returns Boolean from Standard;
    
    Translate(me; theLoc        : Location from TopLoc;
    	    	       theTarget     : in out Persistent from BinObjMgt;
		       theMap        : out SRelocationTable from BinObjMgt);
    ---Purpose: Translate transient location to storable
    
    SetSharedLocations(me: mutable;
                       theLocations:  in LocationSetPtr  from BinTools);
    ---C++: inline
    
fields
    myLocations : LocationSetPtr   from BinTools;
end;
