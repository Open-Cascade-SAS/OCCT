-- Created on: 1997-07-28
-- Created by: Pierre CHALAMET
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class Texture1D from Graphic3d

inherits TextureMap from Graphic3d

  ---Purpose: This is an abstract class for managing 1D textures.

uses

  TypeOfTexture   from Graphic3d,
  NameOfTexture1D from Graphic3d,
  AsciiString     from TCollection,
  PixMap_Handle   from Image

raises

  OutOfRange from Standard

is

  Initialize (theFileName : AsciiString from TCollection;
              theType     : TypeOfTexture from Graphic3d);

  Initialize (theName : NameOfTexture1D from Graphic3d;
              theType : TypeOfTexture   from Graphic3d);

  Initialize (thePixMap : PixMap_Handle from Image;
              theType   : TypeOfTexture from Graphic3d);

  Name (me) returns NameOfTexture1D from Graphic3d;
  ---Purpose:
  -- Returns the name of the predefined textures or NOT_1D_UNKNOWN
  -- when the name is given as a filename.
  ---Level: Public

  NumberOfTextures (myclass) returns Integer from Standard;
  ---Purpose:
  -- Returns the number of predefined textures.
  ---Level: Public

  TextureName (myclass; aRank: Integer from Standard)
  returns AsciiString from TCollection
  raises OutOfRange from Standard;
  ---Purpose:
  -- Returns the name of the predefined texture of rank <aRank>
  ---Trigger: when <aRank> is < 1 or > NumberOfTextures.
  ---Level: Public

fields

  myName : NameOfTexture1D from Graphic3d;

end Texture1D;
