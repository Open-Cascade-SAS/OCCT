-- Created on: 1998-08-18
-- Created by: Yves FRICAUD
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Association from TopOpeBRepDS inherits TShared from MMgt

	---Purpose: 

uses
    Interference                            from TopOpeBRepDS,
    ListOfInterference                      from TopOpeBRepDS,
    DataMapOfInterferenceListOfInterference from TopOpeBRepDS

is

    Create returns mutable Association from TopOpeBRepDS;
    
    Associate  (me : mutable; I,K : Interference from TopOpeBRepDS) 
    is static;
     
    Associate  (me : mutable; 
    	    	I  : Interference      from TopOpeBRepDS;
    	    	LI : ListOfInterference from TopOpeBRepDS) 
    is static;
    HasAssociation (me ; I : Interference from TopOpeBRepDS)
    returns Boolean from Standard
    is static;
    
    Associated (me : mutable ; I : Interference from TopOpeBRepDS) 
    ---C++: return &
    returns ListOfInterference from TopOpeBRepDS
    is static;
    
    AreAssociated (me; I,K : Interference from TopOpeBRepDS)
    returns Boolean from Standard
    is static;
    
fields

    myMap : DataMapOfInterferenceListOfInterference from TopOpeBRepDS;
    
end Association;
