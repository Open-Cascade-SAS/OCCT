-- File:	StepToTopoDS_MakeTransformed.cdl
-- Created:	Mon Apr 28 14:13:07 1997
-- Author:	Christian CAILLET
--		<cky@heliox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1997


class MakeTransformed  from StepToTopoDS    inherits Root

    ---Purpose : Produces instances by Transformation of a basic item

uses Trsf from gp, Shape from TopoDS,
     TransientProcess from Transfer,
     Axis2Placement3d from StepGeom,
     CartesianTransformationOperator3d from StepGeom,
     MappedItem       from StepRepr

is

    Create returns MakeTransformed;

    Compute (me : in out; Origin, Target : Axis2Placement3d from StepGeom)
    	returns Boolean;
    ---Purpose : Computes a transformation to pass from an Origin placement to
    --           a Target placement. Returns True when done
    --           If not done, the transformation will by Identity

    Compute (me : in out; Operator : CartesianTransformationOperator3d from StepGeom)  returns Boolean;
    ---Purpose : Computes a transformation defined by an operator 3D

    Transformation (me) returns Trsf from gp;
    ---Purpose : Returns the computed transformation (Identity if not yet or
    --           if failed)
    ---C++ : return const &

    Transform      (me; shape : in out Shape from TopoDS) returns Boolean;
    ---Purpose : Applies the computed transformation to a shape
    --           Returns False if the transformation is Identity


    TranslateMappedItem (me : in out; mapit : MappedItem from StepRepr;
    	    	    	 TP : mutable TransientProcess from Transfer)
    	returns Shape;
    ---Purpose : Translates a MappedItem. More precisely
    --           A MappedItem has a MappingSource and a MappingTarget
    --           MappingSource has a MappedRepresentation and a MappingOrigin
    --           MappedRepresentation is the basic item to be instanced
    --           MappingOrigin is the starting placement
    --           MappingTarget is the final placement
    --           
    --           Hence, the transformation from MappingOrigin and MappingTarget
    --           is computed, the MappedRepr. is converted to a Shape, then
    --           transformed as an instance of this Shape

fields

    theTrsf : Trsf from gp;

end MakeTransformed;
