-- Created on: 1991-05-14
-- Created by: Annick PANCHER
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Revised:     Mireille MERCIEN


deferred generic class Compare from TCollection ( Item as any )

	---Purpose: Defines a comparison operator which can be used by
	-- any ordered structure.   The  way to compare items
	-- has  to be described  in  subclasses, which inherit
	-- from instantiations of Compare.

is

    IsLower (me; Left, Right: Item)
	---Level: Public
	---Purpose: returns True if <Left> is lower than <Right>.
    returns Boolean
    is virtual;
    
    IsGreater (me; Left, Right: Item)
	---Level: Public
	---Purpose: returns True if <Left> is greater than <Right>.
    returns Boolean
    is virtual;

    IsEqual(me; Left, Right: Item)
	---Level: Public
	---Purpose: returns True when <Right> and <Left> are equal.
    returns Boolean
    is virtual;
	
end;


