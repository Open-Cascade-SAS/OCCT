-- Created on: 1997-07-28
-- Created by: Pierre CHALAMET
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class TextureMap from Graphic3d

inherits TextureRoot from Graphic3d

  ---Purpose: This is an abstract class for managing texture applyable on polygons.

uses 

  TypeOfTexture from Graphic3d,
  TextureParams from Graphic3d,
  LevelOfTextureAnisotropy from Graphic3d,
  AsciiString   from TCollection

is

  Initialize (theFileName : AsciiString from TCollection;
              theType     : TypeOfTexture from Graphic3d);

  EnableSmooth (me : mutable);
  ---Level: public
  ---Purpose:
  -- enable texture smoothing

  IsSmoothed (me) returns Boolean from Standard;
  ---Level: public
  ---Purpose:
  -- Returns TRUE if the texture is smoothed.

  DisableSmooth (me : mutable);
  ---Level: public
  ---Purpose:
  -- disable texture smoothing

  EnableModulate (me : mutable);
  ---Level: public
  ---Purpose:
  -- enable texture modulate mode.
  -- the image is modulate with the shading of the surface.

  DisableModulate (me : mutable);
  ---Level: public
  ---Purpose:
  -- disable texture modulate mode.
  -- the image is directly decal on the surface.

  IsModulate (me) returns Boolean from Standard;
  ---Level: public
  ---Purpose:
  -- Returns TRUE if the texture is modulate.

  EnableRepeat (me : mutable);
  ---Level: public
  ---Purpose:
  -- use this methods if you want to enable
  -- texture repetition on your objects.

  DisableRepeat (me : mutable);
  ---Level: public
  ---Purpose:
  -- use this methods if you want to disable
  -- texture repetition on your objects.

  IsRepeat (me) returns Boolean from Standard;
  ---Level: public
  ---Purpose:
  -- Returns TRUE if the texture repeat is enable.

  AnisoFilter (me) returns LevelOfTextureAnisotropy from Graphic3d;
  ---Level   : public
  ---Purpose : @return level of anisontropy texture filter.
  -- Default value is Graphic3d_LOTA_OFF.

  SetAnisoFilter (me : mutable;
                  theLevel : LevelOfTextureAnisotropy from Graphic3d);
  ---Level   : public
  ---Purpose : @param theLevel level of anisontropy texture filter.

end TextureMap from Graphic3d;
