-- File     : Prs2d_RadiusIndep.cdl
-- Created  : October 2000
-- Author   : Tanya COOL
---Copyright: Matra Datavision 2000

class RadiusIndep from Prs2d inherits Line from Graphic2d

 ---Purpose: Constructs the primitive Radius

uses

	Drawer	           from Graphic2d,
	GraphicObject      from Graphic2d,
    Pnt2d              from gp,
	ExtendedString     from TCollection, 
    TypeOfRadius       from Prs2d,
    Arrow              from Prs2d,
    Array1OfShortReal  from TShort,
    FStream            from Aspect 
	
raises 

    ConstructionError from Standard
       
is
	Create( aGO           : GraphicObject  from Graphic2d; 
	        anAttachPnt   : Pnt2d          from gp; 
            aCenter       : Pnt2d          from gp;
            aRad          : Real           from Standard; 
            aText         : ExtendedString from TCollection;
            aLength       : Real           from Standard = 10.0;
            aTypeRad      : TypeOfRadius   from Prs2d    = Prs2d_TOR_STANDARD;
            aTxtScale     : Real           from Standard = 1.0) 

	returns mutable RadiusIndep from Prs2d;

    ---Purpose: Creates the radius of the circle <aCenter, aRad> passing through 
    --          the point <anAttachPnt1> on the circle

	----------------------------------------------------
	-- Category: Draw and Pick
	----------------------------------------------------

	Draw( me : mutable; aDrawer: Drawer from Graphic2d )
	is static protected;
	---Level: Internal
	---Purpose: Draws the angle <me>.

    DrawElement( me : mutable; aDrawer: Drawer from Graphic2d;
                 anIndex: Integer from Standard)
        is redefined protected;
    ---Level: Internal
    ---Purpose: Draws element <anIndex> of the radius <me>.

    DrawVertex( me : mutable; aDrawer: Drawer from Graphic2d;
                anIndex: Integer from Standard)
        is redefined protected;
    ---Level: Internal
    ---Purpose: Draws vertex <anIndex> of the radius <me>.

	Pick( me : mutable; X, Y: ShortReal from Standard;
		  aPrecision: ShortReal from Standard;
		  aDrawer: Drawer from Graphic2d)
	returns Boolean from Standard
	is static protected;
	---Level: Internal
	---Purpose: Returns Standard_True if the radius <me> is picked,
	--	    Standard_False if not.
	
    --------------------------------------
	-- Category: Inquire methods
	--------------------------------------
    
    Values( me; 
            anAttPnt, aCenter: out Pnt2d          from gp; 
            aRad             : out Real           from Standard;
            aText            : out ExtendedString from TCollection;
            aLength          : out Real           from Standard;
            aTypeRad         : out TypeOfRadius   from Prs2d;
            aTxtScale        : out Real           from Standard ); 

    ---Level: Internal
    ---Purpose: allows to get the properties of the radius
    
    
    --------------------------------------------
  	-- Category: Modification of the properties
	--------------------------------------------
	
    SetText( me: mutable; aTxt: ExtendedString from TCollection );
	---Level: Public
	---Purpose: Defines the text 

    SetTextScale( me: mutable; aTxtScale: Real from Standard );
	---Level: Public
	---Purpose: Defines the scale factor of text 

    SetTextFont( me: mutable; aTF: Integer from Standard );
    ---Level: Public
	---Purpose: Sets the index of the font of this text to this dimension

    SetFontOfSymb( me: mutable; aFS: Integer from Standard );
    ---Level: Public
	---Purpose: Sets the index of the font of the symbol to this dimension

    DrawSymbol( me: mutable; isDraw: Boolean from Standard );
	---Level: Public
	---Purpose: Sets the flag for drawing additional symbol

    SetSymbolCode( me: mutable; aCode: Integer from Standard );
	---Level: Public
	---Purpose: Sets the ASCII code of the symbol
       
    TextFont( me ) returns Integer from Standard;
    ---Level: Public
	---Purpose: Returns the index of the font of this text of this dimension

    FontOfSymb( me ) returns Integer from Standard;
    ---Level: Public
	---Purpose: Returns the index of the font of the symbol of this dimension

    IsDrawSymbol( me ) returns Boolean from Standard;
    ---Level: Public
	---Purpose: Return true if symbol is drawn, false - in otherwise
	
    SymbolCode( me ) returns Integer from Standard;
    ---Level: Public
	---Purpose: Return ASCII code of the symbol

	Save( me; aFStream: in out FStream from Aspect ) is virtual;
												
fields
 
	myX1           : ShortReal         from Standard;
	myY1           : ShortReal         from Standard;
	myX2           : ShortReal         from Standard;
	myY2           : ShortReal         from Standard;
    myTextScale    : ShortReal         from Standard;
    myText         : ExtendedString    from TCollection;
    myTextX        : ShortReal         from Standard;
    myTextY        : ShortReal         from Standard;
    myTextAng      : ShortReal         from Standard;
    myInside       : Boolean           from Standard;
	myXVert        : Array1OfShortReal from TShort;
	myYVert        : Array1OfShortReal from TShort;
    myIsSymbol     : Boolean           from Standard;
    mySymbCode     : Integer           from Standard;
    myTextFont     : Integer           from Standard;
    mySymbFont     : Integer           from Standard;
    myAttPnt       : Pnt2d             from gp;
    myCenter       : Pnt2d             from gp;
    myRadius       : Real              from Standard;
    myLength       : Real              from Standard;
    myRadType      : TypeOfRadius      from Prs2d;

end RadiusIndep from Prs2d;
