-- Created on: 2002-10-29
-- Created by: Michael SAZONOV
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package BinMDF

        ---Purpose: This package provides classes and methods to
        --          translate a transient DF into a persistent one and
        --          vice versa.
        --          
        --          Driver
        --          
        --          A driver is a tool used to translate a transient
        --          attribute into a persistent one and vice versa.
        --          
        --          Driver Table
        --          
        --          A driver table is an object building links between
        --          object types and object drivers. In the
        --          translation process, a driver table is asked to
        --          give a translation driver for each current object
        --          to be translated.

uses
    TCollection,
    TColStd,
    TDF,
    CDM,
    BinObjMgt

is

    deferred class ADriver; -- Attribute Storage/Retrieve Driver.

    class ReferenceDriver;  -- Driver for reference

    class TagSourceDriver;  -- Driver for TDF_TagSource

    private alias StringIdMap is DataMapOfAsciiStringInteger from TColStd;

    -- Map (Type, ADriver)
    imported TypeADriverMap;
    imported DataMapIteratorOfTypeADriverMap;

    -- Double Map (Type, Integer ID)
    imported TypeIdMap;
    imported DoubleMapIteratorOfTypeIdMap;

    -- Attribute Storage Driver Table.
    class ADriverTable;

    AddDrivers (aDriverTable : ADriverTable  from BinMDF;
                aMsgDrv      : MessageDriver from CDM);
        ---Purpose: Adds the attribute storage drivers to <aDriverTable>.

end BinMDF;
