-- Created on: 1993-12-03
-- Created by: Christophe MARION
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package BRepExtrema

    ---Purpose: This package gives   tools to compute  extrema between
    --          Shapes from BRep.

uses 
    Standard,
    StdFail,
    TopoDS,
    GeomAdaptor,
    BRepAdaptor,
    gp,
    Extrema,
    TColStd,
    TopTools,
    TCollection,
    Bnd
    
is

    ----------------------------------------------------------
    --  Extrema between two Shapes with triangulation.
    ----------------------------------------------------------
    imported Poly;


    ----------------------------------------------------------
    --  Extrema between a Point and an Edge.
    ----------------------------------------------------------
    imported ExtPC;


    ----------------------------------------------------------
    --  Extrema between two Edges.
    ----------------------------------------------------------
    imported ExtCC;


    ----------------------------------------------------------
    --  Extrema between a Point and a Face.
    ----------------------------------------------------------
    imported ExtPF;


    ----------------------------------------------------------
    --  Extrema between an Edge  and a Face.
    ----------------------------------------------------------
    imported ExtCF;


    ----------------------------------------------------------
    --  Extrema between two Faces.
    ----------------------------------------------------------
    imported ExtFF;


    ----------------------------------------------------------
    --  
    ----------------------------------------------------------
    exception UnCompatibleShape inherits DomainError;


    ----------------------------------------------------------
    --  enumeration used to describe the type of the support solution:                                         
    -- 	    IsVertex => The solution is a vertex.
    -- 	    IsOnEdge => The solution belongs to an Edge.
    -- 	    IsInFace => The solution is inside a Face.    
     
    ----------------------------------------------------------
    imported SupportType;


    ----------------------------------------------------------
    -- This  class gives tools  to  compute the minimum distance value
    -- between two shapes and  the corresponding couples of solution points.  
    
    ----------------------------------------------------------
    imported DistShapeShape;


    ----------------------------------------------------------
    --  This class is used to store a solution on a Shape. 
    --  (used only by class DistShapeShape)
    ----------------------------------------------------------
    imported SolutionElem;


    ----------------------------------------------------------
    -- This sequence is used to store all the solution on each Shape.
    ----------------------------------------------------------
    imported SeqOfSolution;

    imported DistanceSS;

end BRepExtrema;
