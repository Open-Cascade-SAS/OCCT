-- Created on: 1992-09-23
-- Created by: Christian CAILLET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class ConnectedComponants  from IFGraph  inherits SubPartsIterator

    	---Purpose : determines Connected Componants in a Graph. They define
    	--           disjoined sets of Entities

uses Graph

is

    Create (agraph : Graph; whole : Boolean) returns ConnectedComponants;
    ---Purpose : creates with a Graph, and will analyse :
    --           whole True  : all the contents of the Model
    --           whole False : sub-parts which will be given later

    Evaluate (me : in out) is redefined;
    ---Purpose : does the computation

    	-- --   Iteration : More-Next-etc... will give the Connected Componants

end ConnectedComponants;
