-- Created on: 1997-07-23
-- Created by: Henri JEANNIN
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package ViewerTest

	---Purpose:

uses
    Draw,
    TCollection,
    TColStd,
    TColgp,
    TopAbs,
    TopTools,
    TopoDS,
    V3d,
    AIS,
    NIS,
    MMgt,
    Quantity

is

    class Tool;
    ---Purpose: to build a context and  set a given context as current
    --          for ViewerTest.



    class EventManager;
    ---Purpose: used to manage mouse event (move,select,shiftselect)
    --          By default the events are transmitted to interactive context.


    class DoubleMapOfInteractiveAndName  instantiates  DoubleMap
    	from  TCollection  (    Transient from Standard,
    	    	    	    	AsciiString  from  TCollection,
    	    	    	    	MapTransientHasher  from  TColStd,
    	    	    	    	AsciiString  from  TCollection);


    -- ----------------------------------------------------------------------
    -- Package methods
    -- ----------------------------------------------------------------------

    Factory (theDI : out Interpretor from Draw);
    ---Purpose: Loads all Draw commands of  V2d & V3d. Used for plugin.

    ---Category: Create the viewer....

    ViewerInit ( thePxLeft,    thePxTop : Integer from Standard = 0;
                thePxWidth, thePxHeight : Integer from Standard = 0;
                theViewName : CString from Standard = "";
                theDisplayName : CString from Standard = "")
    returns AsciiString from TCollection;
    ---Purpose: Creates view with default or custom name
    --          and add this name in map to manage muliple views
    --          implemented in ViewerTest_ViewerCommands.cxx
   
    ---Category: Manage the name of views
    RemoveViewName (theName: AsciiString from TCollection);
    
    InitViewName (theName: AsciiString from TCollection;
                  theView: View from V3d);
    
    GetCurrentViewName returns AsciiString from TCollection;
   
    ---Category: Delete the viewer....
    RemoveView (theViewName:AsciiString from TCollection;
               isContextRemoved:Boolean from Standard= Standard_True);
    ---Purpose: Removes view and clear all maps
    --          with information about its resources if neccessary

    ---Category: Selection in the viewer....

    WClass returns TShared from MMgt is private;
    ---C++:     return const &
    ---Purpose: Returns a window class that implements standard behavior of
    --          all windows of the ViewerTest. This includes usual Open CASCADE
    --          view conventions for mouse buttons (e.g. Ctrl+MB1 for zoom,
    --          Ctrl+MB2 for pan, etc) and keyboard shortcuts.
    --          This method is relevant for MS Windows only and respectively
    --          returns WNT_WClass handle.

    PickShape  (aType      : ShapeEnum from TopAbs;
    	    	MaxPick    : Integer from Standard = 5) returns Shape from TopoDS;
    ---Purpose:  waits until a shape of type <aType> is picked in the AIS Viewer and returns it.
    -- if <aType> == TopAbs_Shape, any shape can be picked...
    -- MaxPick  is the Max number before exiting, if no pick is successfull


    PickShapes (aType      : ShapeEnum from TopAbs;
	        thepicked  : in out HArray1OfShape from TopTools;
    	        MaxPick    : Integer from Standard = 5)
		returns Boolean from Standard;
    ---Purpose: wait until the array is filled with picked shapes.
    --          returns True if the array is filled.
    --          exit if number of unsuccesfull picks =  <MaxPick>

    PickObject(Type      : KindOfInteractive from AIS = AIS_KOI_None;
    	       Signature : Integer from Standard = -1;
    	       MaxPick   : Integer from Standard = 5)
    returns InteractiveObject from AIS;
    ---Purpose: waits until an interactive object of a given Type
    --          and signature is picked (defaut values authorize
    --          selection of any Interactive Object)
    --          exit if number of unsuccesfull picks =  <MaxPick>

    PickObjects(thepicked : in out HArray1OfTransient from TColStd;
    	    	Type      : KindOfInteractive from AIS = AIS_KOI_None;
    	        Signature : Integer from Standard = -1;
    	        MaxPick   : Integer from Standard = 5)
    returns Boolean from Standard;
    ---Purpose: selection of several interactive objects. Number is given
    --          by the size of <thepicked>
    --          exit if number of unsuccesfull picks =  <MaxPick>


    Commands (theCommands : in out Interpretor from Draw);
    AviCommands(theCommands :in out Interpretor from Draw);
    ViewerCommands(theCommands :in out Interpretor from Draw);
    MyCommands (theCommands : in out Interpretor from Draw);   --  My  Own  Com-s
    RelationCommands(theCommands :in out Interpretor from Draw);
    ObjectCommands(theCommands :in out Interpretor from Draw);
    FilletCommands(theCommands :in out Interpretor from Draw);
    VoxelCommands(theCommands :in out Interpretor from Draw);
    OpenGlCommands(theCommands :in out Interpretor from Draw);

    GetMousePosition(xpix,ypix: out Integer from Standard);

    GetViewerFromContext returns Viewer from V3d;

    GetCollectorFromContext returns Viewer from V3d;

    GetAISContext returns InteractiveContext from AIS;
	---C++: return const &
    GetNISContext returns InteractiveContext from NIS;
    ---C++: return &

    SetAISContext (aContext: InteractiveContext from AIS);

    SetNISContext (aContext: InteractiveContext from NIS);

    CurrentView returns View from V3d;
	---C++: return const &
	
    CurrentView (aViou:View from V3d);

    Clear ;

    ---Category: Change behaviour on move,select,... events.

    SetEventManager    (aMgr:EventManager from ViewerTest);
    ---Purpose:      puts  <aMgr>   as     current  eventmanager  (the
    --          move,select,...will be applied to <aMgr>

    UnsetEventManager;
    ---Purpose: removes the last EventManager from the list.

    ResetEventManager;
    ---Purpose: clear the list of EventManagers and
    --          sets the default EventManager as current

    CurrentEventManager returns EventManager from ViewerTest;


    ---Category: privateMethods...


    RemoveSelected;

    StandardModeActivation(Mode  : Integer from Standard);

    GetColorFromName(name: CString from Standard)
    returns NameOfColor from Quantity;

    RedrawAllViews;
    ---Purpose: redraws all defined views.

    SplitParameter (theString : AsciiString from TCollection;
                    theName   : out AsciiString from TCollection;
                    theValue  : out AsciiString from TCollection)
    returns Boolean from Standard;
    ---Purpose: Splits "parameter=value" string into separate
    -- parameter and value strings.
    -- @return TRUE if the string matches pattern "<string>=<empty or string>"

end;
