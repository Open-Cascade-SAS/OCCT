-- Created on: 1998-06-03
-- Created by: data exchange team
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Face from ShapeFix inherits Root from ShapeFix

    ---Purpose: This operator allows to perform various fixes on face
    --          and its wires: fixes provided by ShapeFix_Wire,
    --          fixing orientation of wires, addition of natural bounds,
    --          fixing of missing seam edge,
    --          and detection and removal of null-area wires

uses 

    Surface             from Geom,
    Shape               from TopoDS,
    Face                from TopoDS,
    Wire                from TopoDS,
    BasicMsgRegistrator from ShapeExtend,
    Status              from ShapeExtend,
    Surface             from ShapeAnalysis,
    Wire                from ShapeFix,
    SequenceOfShape     from TopTools,
    WireData            from ShapeExtend,
    Vertex              from TopoDS,
    DataMapOfShapeBox2d from ShapeFix,
    DataMapOfShapeListOfShape from TopTools
is

    Create returns Face from ShapeFix;
        ---Purpose: Creates an empty tool

    Create (face: Face from TopoDS) returns Face from ShapeFix;
        ---Purpose: Creates a tool and loads a face

    ClearModes (me: mutable) is virtual;
        ---Purpose: Sets all modes to default

    Init (me: mutable; face: Face from TopoDS);
        ---Purpose: Loads a whole face already created, with its wires, sense and
        --          location

    Init (me: mutable; surf: Surface from Geom; preci: Real;
    	               fwd: Boolean = Standard_True);
        ---Purpose: Starts the creation of the face
        --          By default it will be FORWARD, or REVERSED if <fwd> is False

    Init (me: mutable; surf: Surface from ShapeAnalysis; preci: Real;
    	               fwd: Boolean = Standard_True);
        ---Purpose: Starts the creation of the face
        --          By default it will be FORWARD, or REVERSED if <fwd> is False

    SetMsgRegistrator (me: mutable; msgreg: BasicMsgRegistrator from ShapeExtend) is redefined;
        ---Purpose: Sets message registrator

    SetPrecision (me: mutable; preci: Real) is redefined;
        ---Purpose: Sets basic precision value (also to FixWireTool)

    SetMinTolerance (me: mutable; mintol: Real) is redefined;
        ---Purpose: Sets minimal allowed tolerance (also to FixWireTool)

    SetMaxTolerance (me: mutable; maxtol: Real) is redefined;
        ---Purpose: Sets maximal allowed tolerance (also to FixWireTool)

    FixWireMode (me: mutable) returns Integer;
        ---C++: return &
        ---C++: inline
        ---Purpose: Returns (modifiable) the mode for applying fixes of 
        --          ShapeFix_Wire, by default True. 

    FixOrientationMode (me: mutable) returns Integer;
        ---C++: return &
        ---C++: inline
        ---Purpose: Returns (modifiable) the fix orientation mode, by default
        --          True. If True, wires oriented to border limited square.

    FixAddNaturalBoundMode (me: mutable) returns Integer;
        ---C++: return &
        ---C++: inline
        ---Purpose: Returns (modifiable) the add natural bound mode.
        --          If true, natural boundary is added on faces that miss them.
        --          Default is False for faces with single wire (they are
        --          handled by FixOrientation in that case) and True for others.

    FixMissingSeamMode (me: mutable) returns Integer;
        ---C++: return &
        ---C++: inline
        ---Purpose: Returns (modifiable) the fix missing seam mode, by default
        --          True. If True, tries to insert seam is missed.

    FixSmallAreaWireMode (me: mutable) returns Integer;
        ---C++: return &
        ---C++: inline
        ---Purpose: Returns (modifiable) the fix small area wire mode, by default
        --          False. If True, drops small wires.
    FixIntersectingWiresMode (me: mutable) returns Integer;
        ---C++: return &
        ---C++: inline
        ---Purpose: Returns (modifiable) the fix intersecting wires mode
        --          by default True.
	
    FixLoopWiresMode (me: mutable) returns Integer;
        ---C++: return &
        ---C++: inline
        ---Purpose: Returns (modifiable) the fix loop wires mode
        --          by default True.
	
    FixSplitFaceMode (me: mutable) returns Integer;
        ---C++: return &
        ---C++: inline
        ---Purpose: Returns (modifiable) the fix split face mode
        --          by default True.
	
    AutoCorrectPrecisionMode (me: mutable) returns Integer;
        ---C++: return &
        ---C++: inline
        ---Purpose: Returns (modifiable) the auto-correct precision mode
        --          by default False.
        
    FixPeriodicDegeneratedMode (me: mutable) returns Integer;
        ---C++: return &
        ---C++: inline
        ---Purpose: Returns (modifiable) the activation flag for periodic
        --          degenerated fix. False by default.
	
    Face (me) returns Face from TopoDS;
        ---C++: inline
        ---Purpose: Returns a face which corresponds to the current state
        --  Warning: The finally produced face may be another one ... but with the
        --          same support

    Result (me) returns Shape from TopoDS;
        ---C++: inline
        ---Purpose: Returns resulting shape (Face or Shell if splitted)
        --          To be used instead of Face() if FixMissingSeam involved

    Add (me: mutable; wire: Wire from TopoDS);
        ---Purpose: Add a wire to current face using BRep_Builder.
        --          Wire is added without taking into account orientation of face
        --          (as if face were FORWARD). 
        ---Warning: Method is retained for compatibility with previous versions.

    Perform (me: mutable) returns Boolean;
        ---Purpose: Performs all the fixes, depending on modes
        -- Function Status returns the status of last call to Perform()
        --          ShapeExtend_OK   : face was OK, nothing done
        --          ShapeExtend_DONE1: some wires are fixed
        --          ShapeExtend_DONE2: orientation of wires fixed
        --          ShapeExtend_DONE3: missing seam added
        --          ShapeExtend_DONE4: small area wire removed
        --          ShapeExtend_DONE5: natural bounds added
        --          ShapeExtend_FAIL1: some fails during fixing wires
        --          ShapeExtend_FAIL2: cannot fix orientation of wires
        --          ShapeExtend_FAIL3: cannot add missing seam
        --          ShapeExtend_FAIL4: cannot remove small area wire

    FixOrientation (me: mutable) returns Boolean;
        ---Purpose: Fixes orientation of wires on the face
        --          It tries to make all wires lie outside all others (according
        --          to orientation) by reversing orientation of some of them. 
        --          If face lying on sphere or torus has single wire and 
        --          AddNaturalBoundMode is True, that wire is not reversed in 
        --          any case (supposing that natural bound will be added).
        --          Returns True if wires were reversed

    FixOrientation (me: mutable; MapWires : in out DataMapOfShapeListOfShape from TopTools)
    returns Boolean;
        ---Purpose: Fixes orientation of wires on the face
        --          It tries to make all wires lie outside all others (according
        --          to orientation) by reversing orientation of some of them. 
        --          If face lying on sphere or torus has single wire and 
        --          AddNaturalBoundMode is True, that wire is not reversed in 
        --          any case (supposing that natural bound will be added).
        --          Returns True if wires were reversed
        --          OutWires return information about out wires + list of
        --          internal wires for each (for performing split face).

    FixAddNaturalBound(me: mutable) returns Boolean;
        ---Purpose: Adds natural boundary on face if it is missing.
        --          Two cases are supported:
        --          - face has no wires
        --          - face lies on geometrically double-closed surface 
        --            (sphere or torus) and none of wires is left-oriented
        --          Returns True if natural boundary was added
    
    FixMissingSeam (me: mutable) returns Boolean;
        ---Purpose: Detects and fixes the special case when face on a closed
        --          surface is given by two wires closed in 3d but with gap in 2d.
        --          In that case it creates a new wire from the two, and adds a 
        --          missing seam edge
        --          Returns True if missing seam was added

    FixSmallAreaWire (me: mutable) returns Boolean;
        ---Purpose: Detects wires with small area (that is less than 
        --          100*Precision::PConfusion(). Removes these wires if they are internal.
        --  Returns : True if at least one small wire removed,
        --    	    False if does nothing.
        
    FixLoopWire(me: mutable; aResWires : out SequenceOfShape from TopTools) returns Boolean;
        ---Purpose: Detects if wire has a loop and fixes this situation by splitting on the few parts.
        --          if wire has a loops and it was splitted Status was set to value ShapeExtend_DONE6.
    	
    SplitEdge (me: mutable; sewd: WireData from ShapeExtend; num: Integer from Standard;
    	    	    	    param: Real from Standard; vert: Vertex from TopoDS;
    	    	    	    preci: Real from Standard; boxes: in out DataMapOfShapeBox2d from ShapeFix)
    returns Boolean from Standard is private;

    SplitEdge (me: mutable; sewd: WireData from ShapeExtend; num: Integer from Standard;
    	    	    	    param1: Real from Standard; param2: Real from Standard;
    	    	    	    vert: Vertex from TopoDS; preci: Real from Standard;
    	    	    	    boxes: in out DataMapOfShapeBox2d from ShapeFix)
    returns Boolean from Standard is private;

    FixIntersectingWires (me: mutable) returns Boolean;
        ---Purpose: Detects and fixes the special case when face has more than one wire
        --          and this wires have intersection point

    FixWiresTwoCoincEdges (me: mutable) returns Boolean;
        ---Purpose: If wire contains two coincidence edges it must be removed
        -- Queries on status after Perform()

    FixSplitFace (me: mutable; MapWires : DataMapOfShapeListOfShape from TopTools)
    returns Boolean;
        ---Purpose: Split face if there are more than one out wire
        --          using inrormation after FixOrientation()
        
    FixPeriodicDegenerated (me: mutable)
    returns Boolean;
        ---Purpose: Fixes topology for a specific case when face is composed
        --          by a single wire belting a periodic surface. In that case
        --          a degenerated edge is reconstructed in the degenerated pole
        --          of the surface. Initial wire gets consistent orientation.
        --          Must be used in couple and before FixMissingSeam routine

    Status (me; status: Status from ShapeExtend) returns Boolean;
        ---Purpose: Returns the status of last call to Perform()
        --          ShapeExtend_OK   : face was OK, nothing done
        --          ShapeExtend_DONE1: some wires are fixed
        --          ShapeExtend_DONE2: orientation of wires fixed
        --          ShapeExtend_DONE3: missing seam added
        --          ShapeExtend_DONE4: small area wire removed
        --          ShapeExtend_DONE5: natural bounds added
        --          ShapeExtend_DONE8: face may be splited
        --          ShapeExtend_FAIL1: some fails during fixing wires
        --          ShapeExtend_FAIL2: cannot fix orientation of wires
        --          ShapeExtend_FAIL3: cannot add missing seam
        --          ShapeExtend_FAIL4: cannot remove small area wire
        ---C++: inline

    FixWireTool (me: mutable) returns Wire from ShapeFix;
        ---Purpose: Returns tool for fixing wires.
        ---C++: inline

fields

    mySurf   : Surface from ShapeAnalysis is protected;
    myFace   : Face from TopoDS is protected;
    myResult : Shape from TopoDS is protected; -- result (shell or face)
    myFixWire: Wire from ShapeFix is protected;
    myFwd    : Boolean is protected;

    myFixWireMode              : Integer;
    myFixOrientationMode       : Integer;
    myFixAddNaturalBoundMode   : Integer;
    myFixMissingSeamMode       : Integer;
    myFixSmallAreaWireMode     : Integer;
    myFixLoopWiresMode         : Integer; -- gka 08.01.2004
    myFixIntersectingWiresMode : Integer; -- skl 23.12.2003
    myFixSplitFaceMode         : Integer; -- skl 03.02.2004
    myAutoCorrectPrecisionMode : Integer; -- skl 26.03.2010
    myFixPeriodicDegenerated   : Integer; -- ssv 29.09.2011
    
    myStatus : Integer is protected;

end Face;
