-- Created on: 1992-11-25
-- Created by: Julia DOROVSKIKH
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


generic class Array1 from XmlObjMgt  (Item as Storable) 

        ---Purpose: The class Array1 represents unidimensionnal 
        -- array of fixed size known at run time. 
        -- The range of the index is user defined.
        --  Warning: Programs clients of such class must be independant
        -- of the range of the first element. Then, a C++ for
        -- loop must be written like this
        --     for (i = A->Lower(); i <= A->Upper(); i++)
uses 
    Element     from XmlObjMgt,
    DOMString   from XmlObjMgt

is
    Create (Low, Up: Integer from Standard) returns Array1;
            ---Purpose: Create an array of lower bound <Low> and 
            -- upper bound <Up>. Range error is raised 
            -- when <Up> is less than <Low>.

    Create (theParent:  Element from XmlObjMgt;
            theName:    DOMString from XmlObjMgt) returns Array1;
            ---Purpose: for restoration from DOM_Element which is child of
            --          theParent:
            --             <theParent ...>
            --                 <theName ...>

    CreateArrayElement (me:in out; theParent: in out Element from XmlObjMgt;
                                   theName  : DOMString from XmlObjMgt);
        ---Purpose: Create DOM_Element representing the array, under 'theParent'

    Element(me) returns Element from XmlObjMgt
                is static;
                ---Purpose:  Returns the DOM element of <me>.
                ---Level: Public
                ---C++: inline
                ---C++: return const &

    Length (me) returns Integer from Standard
                is static;
                ---Purpose:  Returns the number of elements of <me>.
                ---Level: Public
                ---C++: inline

    Lower (me) returns Integer from Standard
                is static;
                ---Purpose: Returns the lower bound.
                ---Level: Public
                ---C++: inline

    Upper (me) returns Integer from Standard
                is static;
                ---Purpose: Returns the upper bound.
                ---Level: Public
                ---C++: inline

    SetValue (me: in out; Index: Integer from Standard;
                          Value: in out Element from XmlObjMgt) 
                is static;
                ---Purpose: Set the <Index>th element of the array to <Value>.
                ---Level: Public

    Value (me; Index: Integer from Standard) returns Element from XmlObjMgt
                is static;
                ---Purpose: Returns the value of <Index>th element of the array.
                ---Level: Public

fields 
    myElement   : Element from XmlObjMgt;
    myFirst     : Integer from Standard;
    myLast      : Integer from Standard;

end Array1;
