-- Created on: 1996-09-04
-- Created by: Christian CAILLET
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DataInfo  from MoniTool

    ---Purpose : Gives informations on an object
    --           Used as template to instantiate Elem, etc
    --           This class is for Transient

uses CString, Transient, Type

is

    Type (myclass; ent : Transient) returns Type;
    ---Purpose : Returns the Type attached to an object
    --           Here, the Dynamic Type of a Transient. Null Type if unknown

    TypeName (myclass; ent : Transient) returns CString;
    ---Purpose : Returns Type Name (string)
    --           Allows to name type of non-handled objects

end DataInfo;
