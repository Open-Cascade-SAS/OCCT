-- Created on: 1991-08-02
-- Created by: Laurent BUCHARD
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.





generic class PolygonTool from IntCurveSurface(
                  ThePoint       as any;
                  ThePolygon     as any;
                  TheBoundingBox as any)

	---Purpose: 

raises  OutOfRange from Standard


is  


    Bounding       (myclass; thePolygon : ThePolygon)
    	    	    returns TheBoundingBox;
    ---Purpose: Give the bounding box of the polygon.
    ---C++: inline 
    ---C++: return const &

    DeflectionOverEstimation
    	    	   (myclass; thePolygon : ThePolygon)
    		   ---C++: inline
		   returns Real from Standard;

    Closed         (myclass; thePolygon : ThePolygon)
    	            ---C++: inline
    	    	    returns Boolean from Standard;

    NbSegments     (myclass; thePolygon : ThePolygon)
                    ---C++: inline
		   returns Integer from Standard;

    BeginOfSeg     (myclass; thePolygon : ThePolygon;
    	    	    Index : in Integer)
		    ---C++: inline
    	    	    returns ThePoint
    	    	    raises OutOfRange from Standard;
                    ---C++: return const &
    ---Purpose: Give the point of range Index in the Polygon. 

    EndOfSeg       (myclass; thePolygon : ThePolygon;
    	    	    Index : in Integer)
		    ---C++: inline
    	    	    returns ThePoint
    	    	    raises OutOfRange from Standard;
		    ---C++: return const &
    ---Purpose: Give the point of range Index in the Polygon. 


    Dump           (myclass; thePolygon : ThePolygon);
		 
end PolygonTool;








