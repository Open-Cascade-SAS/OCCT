-- Created on: 2009-04-06
-- Created by: Sergey ZARITCHNY
-- Copyright (c) 2009-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Axis from TDataXtd inherits Attribute from TDF


	---Purpose: The basis to define an axis attribute.
	--          
	--  Warning: Use TDataXtd_Geometry  attribute  to retrieve  the
	--          gp_Lin of the Axis attribute

uses Attribute       from TDF,
     Label           from TDF,
     GUID            from Standard,
     Line            from Geom,
     Lin             from gp,
     DataSet         from TDF,
     RelocationTable from TDF




is    

   ---Purpose: class methods
    --         =============
    
    GetID(myclass)    
 	---C++: return const & 
    	---Purpose: 	Returns the GUID for an axis. 
    returns GUID from Standard;

    
    Set (myclass ; label : Label from TDF) 
    ---Purpose: Finds or creates an axis attribute defined by the  label.
-- In the case of a creation of an axis, a compatible
-- named shape should already be associated with label.
-- Exceptions
-- Standard_NullObject if no compatible named
-- shape is associated with the label.
    returns Axis from TDataXtd;    

    Set (myclass ; label :  Label from TDF; L : Lin from gp) 
    ---Purpose: Find,  or create,  an Axis  attribute  and set <P>  as
    --          generated in the associated NamedShape.
    returns Axis from TDataXtd;    


    ---Purpose: Axis methods
    --          ============     

    Create
    returns mutable Axis from TDataXtd;  

    ---Category: TDF_Attribute methods
    --           =====================
    
    ID(me)  
    	---C++: return const & 
    returns GUID from Standard;

    Restore(me: mutable; with : Attribute from TDF);

    NewEmpty(me)
    returns mutable Attribute from TDF;

    Paste (me; into : mutable Attribute from TDF;
	       RT   : mutable RelocationTable from TDF);  

    Dump(me; anOS : in out OStream from Standard)
    	returns OStream from Standard
    	is redefined;
	---C++: return &

end Axis;



