-- File:        EvaluatedDegeneratePcurve.cdl
-- Created:     Mon Dec  4 12:02:26 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWEvaluatedDegeneratePcurve from RWStepGeom

	---Purpose : Read & Write Module for EvaluatedDegeneratePcurve

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     EvaluatedDegeneratePcurve from StepGeom,
     EntityIterator from Interface

is

	Create returns RWEvaluatedDegeneratePcurve;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable EvaluatedDegeneratePcurve from StepGeom);

	WriteStep (me; SW : in out StepWriter; ent : EvaluatedDegeneratePcurve from StepGeom);

	Share(me; ent : EvaluatedDegeneratePcurve from StepGeom; iter : in out EntityIterator);

end RWEvaluatedDegeneratePcurve;
