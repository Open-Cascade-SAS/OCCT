-- Created on: 1993-01-14
-- Created by: Isabelle GRIGNON
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

generic class IntCS from IntImp 
    (ThePSurface     as any;
     ThePSurfaceTool as any;
     TheCurve        as any;
     TheCurveTool    as any;
     TheFunction     as any)

    	---Purpose: intersection between a curve and a surface with a close
    	--          point

uses Pnt from gp,
     FunctionSetRoot from math

raises NotDone from StdFail,
       DomainError from Standard    

is

    
    Create( U,V,W       : Real from Standard;
            F           : TheFunction;
	    TolTangency : Real;
    	    MarginCoef  : Real = 0.0)
	    
    	---Purpose: compute the solution point with the close point
    	--          MarginCoef is the coefficient for extension of UV bounds.
    	--          Ex., UFirst -= MarginCoef*(ULast-UFirst)
    	
    returns IntCS from IntImp;
    
    Create( F           : TheFunction;
            TolTangency : Real from Standard)
	    
	    ---Purpose: initialize the parameters to compute the solution

    returns IntCS from IntImp;
    

    Perform(me : in out; U,V,W : Real from Standard;
    	    	    	 Rsnld : in out FunctionSetRoot from math;
    	    	    	 u0,v0,u1,v1,w0,w1 : Real from Standard)
	---Purpose: compute the solution 
	--          it's possible to write to optimize:
	--          IntImp_IntCS inter(S1,C1,Toltangency)
	--          math_FunctionSetRoot rsnld(Inter.function())
	--          while ...{
	--             u=...
	--             v=...
	--             w=...
	--             inter.Perform(u,v,w,rsnld)
	--          }
	--      or
	--          IntImp_IntCS inter(Toltangency)
	--          inter.SetSurface(S);
	--          math_FunctionSetRoot rsnld(Inter.function())
	--          while ...{
	--             C=...  
	--             inter.SetCurve(C);
	--             u=...
	--             v=...
	--             w=...
	--             inter.Perform(u,v,w,rsnld)
	--          }
	--          
    is static;

    IsDone(me) returns Boolean from Standard
        ---Purpose: Returns TRUE if the creation completed without failure.
    is static;

    IsEmpty(me) returns Boolean from Standard
    raises NotDone from StdFail
    is static;
    
    Point(me)
        ---Purpose: returns the intersection point
        --          The exception NotDone is raised if IsDone is false.
    	--          The exception DomainError is raised if IsEmpty is true.

    	returns Pnt from gp
    	---C++: return const &

    	raises NotDone     from StdFail,
	       DomainError from Standard
	
    is static;


    ParameterOnCurve(me) returns Real from Standard
    raises NotDone     from StdFail,
	   DomainError from Standard
	
    is static;
    
    ParameterOnSurface(me;U,V : out Real from Standard)
    raises NotDone     from StdFail,
	   DomainError from Standard
	
    is static;

    Function(me: in out )
    ---Purpose: return the math function which 
    --          is used to compute the intersection
    ---C++: return &
    returns TheFunction
    is static;
    

fields

    done  : Boolean from Standard;
    empty : Boolean from Standard;
    myFunction : TheFunction;
    w     : Real from Standard;
    u     : Real from Standard;
    v     : Real from Standard;
    tol   : Real from Standard;

end IntCS;
