-- Created on: 1999-09-24
-- Created by: Sergey ZARITCHNY
-- Copyright (c) 1999-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Box from QANewBRepNaming  inherits  TopNaming from QANewBRepNaming

    ---Purpose: To load the Box results 

uses MakeBox from BRepPrimAPI,
     Shape   from TopoDS,
     Label   from TDF,
     TypeOfPrimitive3D from QANewBRepNaming

is
 
    Create  returns  Box from QANewBRepNaming;
 
    Create  (ResultLabel :  Label from TDF) 
    returns  Box from QANewBRepNaming;

    Init(me : in out; ResultLabel : Label from TDF);


    Load (me; MakeShape : in out MakeBox from BRepPrimAPI; Type : TypeOfPrimitive3D from QANewBRepNaming);
      ---Purpose : Load  the box in  the data  framework  

    Back (me)   returns Label from TDF;
      ---Purpose : Returns the label of the back face of a box .
    
    Bottom (me) returns Label from TDF;
      ---Purpose : Returns the label of the  bottom face of a box .
    
    Front (me)  returns Label from TDF;
      ---Purpose : Returns the label of the  front face of a box .

    Left (me)   returns Label from TDF;
      ---Purpose : Returns the label of the  left face of a box .

    Right (me)  returns Label from TDF;
      ---Purpose : Returns the  label of the  right face of a box .

    Top (me)    returns Label from TDF;
      ---Purpose : Returns the  label of the  top face of a box . 
    
end Box;
