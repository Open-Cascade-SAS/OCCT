-- File:        RevolvedAreaSolid.cdl
-- Created:     Mon Dec  4 12:02:31 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWRevolvedAreaSolid from RWStepShape

	---Purpose : Read & Write Module for RevolvedAreaSolid

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     RevolvedAreaSolid from StepShape,
     EntityIterator from Interface

is

	Create returns RWRevolvedAreaSolid;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable RevolvedAreaSolid from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : RevolvedAreaSolid from StepShape);

	Share(me; ent : RevolvedAreaSolid from StepShape; iter : in out EntityIterator);

end RWRevolvedAreaSolid;
