-- Created on: 1998-02-18
-- Created by: Jeanine PANCIATICI
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

private  class  InterFunc  from  Adaptor3d  inherits  FunctionWithDerivative  from  math 

         ---Purpose: Used to find the points U(t) = U0 or V(t) = V0 in
         --          order to determine the  Cn discontinuities of  an
         --               Adpator_CurveOnSurface  relativly  to    the
         --          discontinuities of the surface. Used to
         --          find the roots of the functions
	 
uses  
      HCurve2d  from  Adaptor2d
 
raises  ConstructionError

is 
      Create  (C :  HCurve2d  from  Adaptor2d;  FixVal:  Real  from  Standard; 
               Fix:  Integer) 
      returns  InterFunc 
      raises  ConstructionError  from  Standard;  
      ---Purpose:   build the function  U(t)=FixVal   if Fix =1 or 
      --            V(t)=FixVal if Fix=2

    Value(me: in out; X: Real; F: out Real)
        ---Purpose: computes the value <F>of the function for the variable <X>.
    	--         Returns True if the calculation were successfully done, 
    	--          False otherwise.

    returns Boolean;

 
    Derivative(me: in out; X: Real; D: out Real)
         ---Purpose: computes the derivative <D> of the function 
         --          for the variable <X>.
    	--           Returns True if the calculation were successfully done, 
    	--           False otherwise.

    returns Boolean;


    Values(me: in out; X: Real; F, D: out Real)
    	---Purpose: computes the value <F> and the derivative <D> of the 
    	--          function for the variable <X>.
    	--          Returns True if the calculation were successfully done,
    	--          False otherwise.

    returns Boolean;

fields 

    myCurve2d :  HCurve2d    from  Adaptor2d; 
    myFixVal  :  Real  from  Standard;
    myFix    :  Integer     from  Standard; 


    
end InterFunc;
      
