-- Created on: 1997-07-28
-- Created by: Pierre CHALAMET
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class TextureRoot from Graphic3d

inherits TShared from MMgt

  ---Purpose: This is the texture root class enable the dialog with the GraphicDriver allows the loading of texture.

uses

  TextureParams from Graphic3d,
  TypeOfTexture from Graphic3d,
  PixMap        from Image,
  PixMap_Handle from Image,
  Path          from OSD,
  AsciiString   from TCollection

is

  Initialize (theFileName : AsciiString from TCollection;
              theType     : TypeOfTexture from Graphic3d);
  ---Purpose: Creates a texture from a file
  --  Warning: Note that if <FileName> is NULL the texture must be realized
  -- using LoadTexture(image) method.

  Initialize (thePixmap : PixMap_Handle from Image;
              theType   : TypeOfTexture from Graphic3d);
  ---Purpose: Creates a texture from pixmap.
  -- Please note that the implementation expects the image data
  -- to be in Bottom-Up order (see Image_PixMap::IsTopDown()).

  Destroy (me);
  ---C++ : alias ~

  --
  -- public methods
  --

  IsDone (me) returns Boolean from Standard
  is virtual;
  ---Level:   public
  ---Purpose: Checks if a texture class is valid or not.
  -- @return true if the construction of the class is correct

  Path (me) returns Path from OSD;
  ---Level:   public
  ---Purpose:
  -- Returns the full path of the defined texture.
  -- It could be empty path if GetImage() is overridden to load image not from file.
  ---C++: return const &

  Type (me) returns TypeOfTexture from Graphic3d;
  ---Level:   public
  ---Purpose: @return the texture type.

  GetId (me) returns AsciiString from TCollection;
  ---Level:   advanced
  ---Purpose:
  -- This ID will be used to manage resource in graphic driver.
  -- .
  -- Default implementation generates unique ID although inheritors may re-initialize it.
  -- .
  -- Multiple Graphic3d_TextureRoot instancies with same ID
  -- will be treated as single texture with different parameters
  -- to optimize memory usage though this will be more natural
  -- to use same instance of Graphic3d_TextureRoot when possible.
  -- .
  -- Notice that inheritor may set this ID to empty string.
  -- In this case independent graphical resource will be created
  -- for each instance of Graphic3d_AspectFillArea3d where texture will be used.
  -- .
  -- @return texture identifier.
  ---C++: return const &

  GetImage (me) returns PixMap_Handle from Image
  is virtual;
  ---Level   : Public
  ---Purpose :
  -- This method will be called by graphic driver each time when texture resource should be created.
  -- Default constructors allow defining the texture source as path to texture image or directly as pixmap.
  -- If the source is defined as path, then the image will be dynamically loaded when this method is called
  -- (and no copy will be preserved in this class instance).
  -- Inheritors may dynamically generate the image.
  -- Notice, image data should be in Bottom-Up order (see Image_PixMap::IsTopDown())!
  -- @return the image for texture.

  GetParams (me) returns TextureParams from Graphic3d;
  ---Level: public
  ---Purpose: @return low-level texture parameters
  ---C++: return const &

  TexturesFolder (myclass) returns AsciiString from TCollection;
  ---Level   : Public
  ---Purpose :
  -- The path to textures determined from CSF_MDTVTexturesDirectory or CASROOT environment variables.
  -- @return the root folder with default textures.

fields

  myParams : TextureParams from Graphic3d is protected;
  myTexId  : AsciiString from TCollection is protected;
  myPixMap : PixMap_Handle from Image is protected;
  myPath   : Path from OSD is protected;
  myType   : TypeOfTexture from Graphic3d;

end TextureRoot;
