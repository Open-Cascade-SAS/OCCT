-- File:	RWStepBasic_RWProductCategoryRelationship.cdl
-- Created:	Fri Nov 26 16:26:38 1999 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0
-- Copyright:	Matra Datavision 1999

class RWProductCategoryRelationship from RWStepBasic

    ---Purpose: Read & Write tool for ProductCategoryRelationship

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    ProductCategoryRelationship from StepBasic

is
    Create returns RWProductCategoryRelationship from RWStepBasic;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : ProductCategoryRelationship from StepBasic);
	---Purpose: Reads ProductCategoryRelationship

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: ProductCategoryRelationship from StepBasic);
	---Purpose: Writes ProductCategoryRelationship

    Share (me; ent : ProductCategoryRelationship from StepBasic;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWProductCategoryRelationship;
