-- Created by: DAUTRY Philippe
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

--      	---------------------------

---Version:	0.0
--Version	Date		Purpose
--		0.0	Oct 10 1997	Creation


deferred class DeltaOnModification from TDF
    inherits AttributeDelta from TDF

	---Purpose: This class provides default services for an
	--          AttributeDelta on a MODIFICATION action.
	--          
	--          Applying this AttributeDelta means GOING BACK to
	--          the attribute previously registered state.

uses

    Attribute from TDF

-- raises

is

    Initialize(anAttribute: Attribute from TDF)
    	returns DeltaOnModification from TDF;
	---Purpose: Initializes a TDF_DeltaOnModification.

    Apply (me : mutable)
    	is redefined virtual;
    	---Purpose: Applies the delta to the attribute.

end DeltaOnModification;
