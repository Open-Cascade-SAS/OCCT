-- File:	MNaming_NamingRetrievalDriver_1.cdl
-- Created:	Fri Aug 15 17:31:44 2008
-- Author:	Sergey ZARITCHNY <szy@opencascade.com>
---Copyright:	Open CasCade SA 2008

class NamingRetrievalDriver_1 from MNaming inherits ARDriver from MDF

	---Purpose: 

uses RRelocationTable from MDF,
     Attribute        from PDF,
     Attribute        from TDF, 
     MessageDriver    from CDM

is


    Create(theMessageDriver : MessageDriver from CDM)  
    returns mutable NamingRetrievalDriver_1 from MNaming;
    

    VersionNumber(me) returns Integer from Standard;
	---Purpose: Returns the version number from which the driver
	--          is available: 0.

    SourceType(me) returns Type from Standard;
	---Purpose: Returns the type: Naming from PNaming.

    NewEmpty (me)  returns mutable Attribute from TDF;


    Paste(me;
    	  Source     :         Attribute from PDF;
    	  Target     : mutable Attribute from TDF;
    	  RelocTable : RRelocationTable  from MDF);


end NamingRetrievalDriver_1;
