-- Created on: 1992-09-22
-- Created by: Gilles DEBARBOUILLE
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package MAT

uses
    MMgt,
    TCollection,
    TColStd

is
   
    --------------------------------------------------
    --  Classes of exploration of the Bisecting Locus.
    --------------------------------------------------
    enumeration Side is Left,Right end Side;
    	--- Purpose: Definition on the Left and the Right on the Fig.

    class Graph;

    class Arc;

    class Node;

    class BasicElt;

    class Zone;

    imported SequenceOfBasicElt; 
						     
    imported SequenceOfArc;  

    imported DataMapOfIntegerArc;

    imported DataMapIteratorOfDataMapOfIntegerArc;

    imported DataMapOfIntegerBasicElt;

    imported DataMapIteratorOfDataMapOfIntegerBasicElt;
 
    imported DataMapOfIntegerNode;
 
    imported DataMapIteratorOfDataMapOfIntegerNode;
 
 
    --------------------------------------------------- 
    --  Classes used for the computation of the Mat.
    --------------------------------------------------- 

    generic class TList, TListNode;

    class Bisector;
	
    imported DataMapOfIntegerBisector;
	
    imported DataMapIteratorOfDataMapOfIntegerBisector;
				 
    class ListOfBisector instantiates TList from MAT (Bisector from MAT);
    
    class Edge;
    
    class ListOfEdge instantiates TList from MAT (Edge from MAT);
    
end MAT;




