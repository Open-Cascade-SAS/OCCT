-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class AutoDesignGeneralOrgItem from StepAP214 inherits SelectType from StepData

	-- <AutoDesignGeneralOrgItem> is an EXPRESS Select Type construct translation.
	-- it gathers : Product, ProductDefinition, ProductDefinitionFormation, Representation

uses
     AutoDesignDocumentReference from StepAP214,
     ExternallyDefinedRepresentation from StepRepr,
     Product from StepBasic,
     ProductDefinition from StepBasic,
     ProductDefinitionFormation from StepBasic,
     ProductDefinitionRelationship from StepBasic,
     ProductDefinitionWithAssociatedDocuments from StepBasic,
     Representation from StepRepr
is

	Create returns AutoDesignGeneralOrgItem;
	---Purpose : Returns a AutoDesignGeneralOrgItem SelectType

	CaseNum (me; ent : Transient) returns Integer;
	---Purpose: Recognizes a AutoDesignGeneralOrgItem Kind Entity that is :
	-- 1     Product from StepBasic,
	-- 2     ProductDefinition from StepBasic,
	-- 3     ProductDefinitionFormation from StepBasic,
	-- 4     ProductDefinitionRelationship from StepBasic,
	-- 5     ProductDefinitionWithAssociatedDocuments from StepBasic,
	-- 6     Representation from StepRepr
	-- 7     ExternallyDefinedRepresentation from StepRepr,
	-- 8     AutoDesignDocumentReference from StepAP214,
	--        0 else

	Product (me) returns any Product;
	---Purpose : returns Value as a Product (Null if another type)

	ProductDefinition (me) returns any ProductDefinition;
	---Purpose : returns Value as a ProductDefinition (Null if another type)

	ProductDefinitionFormation (me) returns any ProductDefinitionFormation;
	---Purpose : returns Value as a ProductDefinitionFormation (Null if another type)

	ProductDefinitionRelationship (me) returns any ProductDefinitionRelationship;
	---Purpose : returns Value as a ProductDefinitionRelationship (Null if another type)

	ProductDefinitionWithAssociatedDocuments (me) returns any ProductDefinitionWithAssociatedDocuments;
	---Purpose : returns Value as a ProductDefinitionWithAssociatedDocuments (Null if another type)

	Representation (me) returns any Representation;
	---Purpose : returns Value as a Representation (Null if another type)

	ExternallyDefinedRepresentation (me) returns any ExternallyDefinedRepresentation;
	---Purpose : returns Value as a Representation (Null if another type)

    	AutoDesignDocumentReference (me) returns AutoDesignDocumentReference;

end AutoDesignGeneralOrgItem;
