-- File:	PTopoDS_Wire.cdl
-- Created:	Wed May  5 16:55:49 1993
-- Author:	Remi LEQUETTE
--		<rle@sdsun1>
---Copyright:	 Matra Datavision 1993



class Wire from PTopoDS inherits HShape from PTopoDS

is
    Create returns mutable Wire from PTopoDS;
    	---Level: Internal 

end Wire;
