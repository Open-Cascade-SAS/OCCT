-- Created on: 1999-02-26
-- Created by: Christian CAILLET
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SetLabel  from IGESSelect    inherits ModelModifier from IGESSelect

    ---Purpose : Sets/Clears Short Label of Entities, those designated by the
    --           Selection. No Selection means all the file
    --           
    --           May enforce, else it sets only if no label is yet set
    --           Mode : 0 to clear (always enforced)
    --                  1 to set label to DE number (changes it if already set)

uses AsciiString from TCollection,
     IGESModel, CopyTool, ContextModif
 
is

    Create (mode : Integer; enforce : Boolean) returns SetLabel;
    ---Purpose : Creates a SetLabel for IGESEntity
    --           Mode : see Purpose of the class

    Performing (me; ctx : in out ContextModif;
                target  : IGESModel;
                TC      : in out CopyTool);
    ---Purpose : Specific action : Sets or Clears the Label

    Label (me) returns AsciiString from TCollection;
    ---Purpose : Returns a text which is
    --           "Clear Short Label"  or  "Set Label to DE"
    --           With possible additional information " (enforced)"

fields

    themode  : Integer;
    theforce : Boolean;

end SetLabel;
