-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class AutoDesignActualDateAssignment from StepAP214 

inherits DateAssignment from StepBasic 

uses

	HArray1OfAutoDesignDatedItem from StepAP214, 
	AutoDesignDatedItem from StepAP214, 
	Date from StepBasic, 
	DateRole from StepBasic
is

	Create returns mutable AutoDesignActualDateAssignment;
	---Purpose: Returns a AutoDesignActualDateAssignment


	Init (me : mutable;
	      aAssignedDate : mutable Date from StepBasic;
	      aRole : mutable DateRole from StepBasic) is redefined;

	Init (me : mutable;
	      aAssignedDate : mutable Date from StepBasic;
	      aRole : mutable DateRole from StepBasic;
	      aItems : mutable HArray1OfAutoDesignDatedItem from StepAP214) is virtual;

	-- Specific Methods for Field Data Access --

	SetItems(me : mutable; aItems : mutable HArray1OfAutoDesignDatedItem);
	Items (me) returns mutable HArray1OfAutoDesignDatedItem;
	ItemsValue (me; num : Integer) returns AutoDesignDatedItem;
	NbItems (me) returns Integer;

fields

	items : HArray1OfAutoDesignDatedItem from StepAP214; -- a SelectType

end AutoDesignActualDateAssignment;
