-- Created on: 1993-01-11
-- Created by: Christian CAILLET
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SelectIntersection  from IFSelect  inherits SelectCombine

    ---Purpose : A SelectIntersection filters the Entities issued from several
    --           other Selections as Intersection of results : "AND" operator

uses AsciiString from TCollection, EntityIterator, Graph

is

    Create returns SelectIntersection;
    ---Purpose : Creates an empty SelectIntersection

    RootResult (me; G : Graph) returns EntityIterator;
    ---Purpose : Returns the list of selected Entities, which is the common part
    --           of results from all input selections. Uniqueness is guaranteed.

    Label (me) returns AsciiString from TCollection;
    ---Purpose : Returns a text defining the criterium : "Intersection (AND)"

end SelectIntersection;
