-- Created on: 1998-04-02
-- Created by: Christian CAILLET
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class SignLevelNumber  from IGESSelect    inherits Signature  from IFSelect

    ---Purpose : Gives D.E. Level Number under two possible forms :
    --           * for counter : "LEVEL nnnnnnn", " NO LEVEL", " LEVEL LIST"
    --           * for selection : "/nnn/", "/0/", "/1/2/nnn/"
    --           
    --           For matching, giving /nn/ gets any entity attached to level nn
    --           whatever simple or in a level list

uses CString, Transient, AsciiString, InterfaceModel

is

    Create (countmode : Boolean) returns mutable SignLevelNumber;
    ---Purpose : Creates a SignLevelNumber
    --           <countmode> True : values are naturally displayed
    --           <countmode> False: values are separated by slashes
    --             in order to allow selection by signature by Draw or C++

    Value   (me; ent : any Transient; model : InterfaceModel) returns CString;
    ---Purpose : Returns the value (see above)

fields

    thecountmode : Boolean;

end SignLevelNumber;
