-- Created on: 1996-07-05
-- Created by: Jean-Louis Frenkel
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package PTColStd

uses
    Standard,TColStd,TCollection
   ---Category:  reusable class
   --           
is

   class MapPersistentHasher instantiates MapHasher from TCollection(Persistent);

   class DoubleMapOfTransientPersistent  instantiates   
	     DoubleMap from TCollection(Transient from Standard,
      	    	    	    	 Persistent from Standard,
      	    	    	    	 MapTransientHasher from TColStd,
    	    	    	    	 MapPersistentHasher from PTColStd);  

   class TransientPersistentMap instantiates 
   DataMap from TCollection(Transient from Standard,
                            Persistent from Standard,
	       	            MapTransientHasher from TColStd);
    
   class PersistentTransientMap instantiates
   DataMap from TCollection(Persistent from Standard,
                             Transient from Standard,
                             MapPersistentHasher from PTColStd);

end PTColStd;
