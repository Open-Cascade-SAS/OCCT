-- Created on: 1997-09-22
-- Created by: VAUTHIER Jean-Claude
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Chamfer from QANewBRepNaming inherits TopNaming from QANewBRepNaming

    ---Purpose: To load the Chamfer results

uses 
 
    MakeChamfer from BRepFilletAPI,
    Shape       from TopoDS,
    Label       from TDF

is
 
    Create returns Chamfer from QANewBRepNaming; 

    Create(ResultLabel : Label from TDF) 
    returns Chamfer from QANewBRepNaming; 

    Init(me : in out; ResultLabel :  Label from TDF);


    Load (me; part      : in     Shape       from TopoDS;
    	      mkChamfer : in out MakeChamfer from BRepFilletAPI);

    FacesFromEdges (me) 
    ---Purpose: Returns the label of faces generated from edges
    returns Label from TDF;
    
    ModifiedFaces (me)
    ---Purpose: Returns the label of modified faces 
    returns Label from TDF;

    DeletedFaces (me)
    ---Purpose: Returns the label of deleted faces 
    returns Label from TDF;

end Chamfer;
