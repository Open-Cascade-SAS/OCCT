-- File:        RWStepRepr.cdl
-- Created:     Mon Dec  4 12:02:22 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




package RWStepRepr 

uses

	StepData, Interface, TCollection, TColStd, StepRepr

is


--class ReadWriteModule;

--class GeneralModule;

class RWDefinitionalRepresentation;
class RWDescriptiveRepresentationItem;
class RWFunctionallyDefinedTransformation;
class RWGlobalUncertaintyAssignedContext;
class RWGlobalUnitAssignedContext;
class RWItemDefinedTransformation;
--moved to StepBasic: class RWGroup;
--moved to StepBasic: class RWGroupRelationship;
class RWMappedItem;
class RWParametricRepresentationContext;
class RWProductDefinitionShape;
class RWPropertyDefinition;
class RWPropertyDefinitionRepresentation;
--moved to StepAP214: class RWRepItemGroup;
class RWRepresentation;
class RWRepresentationContext;
class RWRepresentationItem;
class RWRepresentationMap;
class RWRepresentationRelationship;

class RWShapeAspect;
class RWShapeAspectRelationship;
class RWShapeAspectTransition;
-- class RWShapeDefinitionRepresentation;  moved to StepShape

    	-- Added from AP214 CC1 to CC2

class RWMakeFromUsageOption;
class RWAssemblyComponentUsage;
class RWQuantifiedAssemblyComponentUsage;
class RWSpecifiedHigherUsageOccurrence;

class RWAssemblyComponentUsageSubstitute;

class RWRepresentationRelationshipWithTransformation;
class RWShapeRepresentationRelationshipWithTransformation;

class RWMaterialDesignation;

-- ABV added for CAX TRJ 2 validation properties
class RWMeasureRepresentationItem;

    -- Added for AP203
    class RWConfigurationDesign;
    class RWConfigurationEffectivity;
    class RWConfigurationItem;
    class RWProductConcept;

    -- Added for Dimensional Tolerancing (CKY 25 APR 2001 for TR7J)
    class RWCompoundRepresentationItem;

	---Package Method ---

--- added for AP209
    class RWDataEnvironment;
    class RWMaterialPropertyRepresentation;
    class RWPropertyDefinitionRelationship;
    class RWMaterialProperty;
    class RWStructuralResponseProperty;
    class RWStructuralResponsePropertyDefinitionRepresentation;

--- added for TR12J (GD&T) 
    class RWCompositeShapeAspect;
    class RWDerivedShapeAspect;
    class RWExtension;
    class RWShapeAspectDerivingRelationship;
    class RWReprItemAndLengthMeasureWithUnit;
    
--	Init;
	---Purpose: enforced the initialisation of the  libraries

end RWStepRepr;
