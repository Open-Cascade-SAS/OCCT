-- Created on: 1998-02-19
-- Created by: s:	Gerard GRAS
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



private class BackgroundGraphicObject from V2d inherits GraphicObject from Graphic2d 

	---Version:

	---Purpose: Creates a 2D background graphic object in a view.
	--	    A graphic object is a primitives manager
	--	    which drawn before all the others graphic objects

	---Keywords:
	---Warning:
	---References:

uses
	View                    from Graphic2d

is
	-------------------------
	-- Category: Constructors
	-------------------------

        Create (aView: View from Graphic2d)
        returns mutable BackgroundGraphicObject from V2d;
        ---Level: Public
        ---Purpose: Creates a graphic object in the view <aView>.
        --          A graphic object manages a sequence of primitives.
        ---Category: Constructors

	-------------------------------------------------
	-- Category: Methods to manage the drawing priority 
	-------------------------------------------------

	MaxPriority (me) returns Integer from Standard is redefined;
	---Level: Public
	---Purpose: Returns the max usable relative priority of the 
	--         "hiding" graphic object. 	

        ----------------------------
        -- Category: Private methods
        ----------------------------

        BasePriority (me) returns Integer from Standard is redefined private;
        ---Level: Internal
        ---Purpose: Returns the min usable absolute priority of the
        --         "hiding" graphic object.  

end BackgroundGraphicObject from V2d;
