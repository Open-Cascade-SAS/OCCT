-- Created on: 1995-10-24
-- Created by: Mister rmi
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Polygon2D from PPoly inherits Persistent from Standard

    	---Purpose: This class represents a 2d polygon.
    	--          
    	--          It is defined by an array of 2d nodes values.
    	--          If the Polygon2D is closed, the point will be
    	--          repeated.


uses HArray1OfPnt2d  from PColgp

is

    Create(Nodes: HArray1OfPnt2d from PColgp;
    	   Defl : Real from Standard) 
    returns mutable Polygon2D from PPoly;
    	---Purpose: Defaults with allocation of nodes.
    
    Deflection(me) returns Real;

    Deflection(me : mutable; Defl : Real from Standard);
    
    NbNodes(me) returns Integer;
    
    Nodes(me) returns HArray1OfPnt2d from PColgp;

    Nodes(me : mutable; Nodes : HArray1OfPnt2d from PColgp);
    
fields

    myDeflection: Real;
    myNodes:      HArray1OfPnt2d from PColgp;

end Polygon2D;
