-- File:	StepFEA_CurveElementLocation.cdl
-- Created:	Thu Dec 12 17:51:04 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class CurveElementLocation from StepFEA
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity CurveElementLocation

uses
    FeaParametricPoint from StepFEA

is
    Create returns CurveElementLocation from StepFEA;
	---Purpose: Empty constructor

    Init (me: mutable; aCoordinate: FeaParametricPoint from StepFEA);
	---Purpose: Initialize all fields (own and inherited)

    Coordinate (me) returns FeaParametricPoint from StepFEA;
	---Purpose: Returns field Coordinate
    SetCoordinate (me: mutable; Coordinate: FeaParametricPoint from StepFEA);
	---Purpose: Set field Coordinate

fields
    theCoordinate: FeaParametricPoint from StepFEA;

end CurveElementLocation;
