-- File:        SurfaceStyleSegmentationCurve.cdl
-- Created:     Mon Dec  4 12:02:32 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWSurfaceStyleSegmentationCurve from RWStepVisual

	---Purpose : Read & Write Module for SurfaceStyleSegmentationCurve

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     SurfaceStyleSegmentationCurve from StepVisual,
     EntityIterator from Interface

is

	Create returns RWSurfaceStyleSegmentationCurve;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable SurfaceStyleSegmentationCurve from StepVisual);

	WriteStep (me; SW : in out StepWriter; ent : SurfaceStyleSegmentationCurve from StepVisual);

	Share(me; ent : SurfaceStyleSegmentationCurve from StepVisual; iter : in out EntityIterator);

end RWSurfaceStyleSegmentationCurve;
