-- Created on: 1998-05-06
-- Created by: Christian CAILLET
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package SWDRAW

    ---Purpose: Provides DRAW interface to the functionalities of Shape Healing
    --          toolkit (SHAPEWORKS Delivery Unit).
    --          
    --          Classes prefixed with Shape* corresponds to the packages of
    --          Shape Healing.

uses  TCollection, TColStd, TopoDS, TopTools, Draw, ShapeProcessAPI

is

    class ShapeTool;
    	---Purpose: Contains commands to activate Topology/Geometry not
    	--          Shape Healing

    class ShapeAnalysis;
    	---Purpose: Contains commands to activate package ShapeAnalysis

    class ShapeBuild;
    	---Purpose: Contains commands to activate package ShapeBuild

    class ShapeConstruct;
    	---Purpose: Contains commands to activate package ShapeConstruct

    class ShapeCustom;
    	---Purpose: Contains commands to activate package ShapeCustom

    class ShapeExtend;
    	---Purpose: Contains commands to activate package ShapeExtend

    class ShapeFix;
    	---Purpose: Contains commands to activate package ShapeFix

    class ShapeUpgrade;
    	---Purpose: Contains commands to activate package ShapeUpgrade

    class ShapeProcess;
    	---Purpose: Contains commands to activate package ShapeProcess
    
    class ShapeProcessAPI;
    	---Purpose: Contains commands to activate package ShapeProcessAPI
	
    class ToVRML;
    	---Purpose: A utility which writes a Shape to VRML format
    	---Remark : It can be placed elsewhere, while it depends on
    	--          only BRepMesh i.e. TOPOLOGY

    Init (theCommands: in out Interpretor from Draw);
    	---Purpose: Loads commands defined in SWDRAW

    GroupName returns CString is private;
    	---Purpose: Returns the name of the DRAW group accumulating the
    	--          commands from the classes prefixed with Shape*.
	--          Returns "Shape Healing".
	
end SWDRAW;
