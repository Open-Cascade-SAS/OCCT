-- Created on: 1995-12-06
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




package BRepCheck 

	---Purpose: This package  provides tools to check the validity
	--          of the BRep.

uses MMgt,
     StdFail,
     TCollection,
     TopAbs,
     Adaptor3d,
     TopoDS,
     BRep,
     TopTools

is

    deferred class Result;   -- inherits TShared from MMgt
    
    class Vertex;            -- inherits Shape
    
    class Edge;              -- inherits Shape
    
    class Wire;              -- inherits Shape
    
    class Face;              -- inherits Shape
    
    class Shell;             -- inherits Shape
    
--    class Solid;             -- inherits Shape

    class Analyzer;


    enumeration Status is
      NoError,
      
      -- for vertices
      InvalidPointOnCurve,
      InvalidPointOnCurveOnSurface,
      InvalidPointOnSurface,
            
      -- for edges
      No3DCurve,
      Multiple3DCurve,
      Invalid3DCurve,
      NoCurveOnSurface,
      InvalidCurveOnSurface,
      InvalidCurveOnClosedSurface,
      InvalidSameRangeFlag,
      InvalidSameParameterFlag,
      InvalidDegeneratedFlag,
      
      FreeEdge,
      InvalidMultiConnexity,
      InvalidRange,
      
      
      -- for wires
      EmptyWire,
      RedundantEdge,
      SelfIntersectingWire, -- on a face

      -- for faces
      NoSurface,
      InvalidWire,
      RedundantWire,
      IntersectingWires,
      InvalidImbricationOfWires,

      -- for shells
      EmptyShell,
      RedundantFace,


      -- for shapes
      UnorientableShape,
      NotClosed,
      NotConnected,
      
      SubshapeNotInShape,
      
      BadOrientation,
      BadOrientationOfSubshape,
      
      InvalidToleranceValue,

      -- for exception
      CheckFail
    
    end Status;


    class ListOfStatus instantiates List from TCollection
        (Status from BRepCheck);
       
    class DataMapOfShapeListOfStatus instantiates DataMap from TCollection 
        (Shape          from TopoDS,
       	 ListOfStatus   from BRepCheck,
         ShapeMapHasher from TopTools);
	
	
    class DataMapOfShapeResult instantiates DataMap from TCollection
    	(Shape          from TopoDS,
       	 Result         from BRepCheck,
         OrientedShapeMapHasher from TopTools);
	 
	 
    -- Package method

    Add(List: in out ListOfStatus from BRepCheck; 
        Stat: Status from BRepCheck);



    Print(Stat: Status from BRepCheck;
          OS: in out OStream from Standard);

    SelfIntersection(W      : Wire from TopoDS;
    	    	   F      : Face from TopoDS;
                   E1 : out Edge from TopoDS;
                   E2 : out Edge from TopoDS)
      returns Boolean from Standard;
      
end BRepCheck;
