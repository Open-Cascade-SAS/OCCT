-- Created on: 1999-11-26
-- Created by: Andrey BETENEV
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0

class ConfigurationDesign from StepRepr
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity ConfigurationDesign

uses
    ConfigurationItem from StepRepr,
    ConfigurationDesignItem from StepRepr

is
    Create returns ConfigurationDesign from StepRepr;
	---Purpose: Empty constructor

    Init (me: mutable; aConfiguration: ConfigurationItem from StepRepr;
                       aDesign: ConfigurationDesignItem from StepRepr);
	---Purpose: Initialize all fields (own and inherited)

    Configuration (me) returns ConfigurationItem from StepRepr;
	---Purpose: Returns field Configuration
    SetConfiguration (me: mutable; Configuration: ConfigurationItem from StepRepr);
	---Purpose: Set field Configuration

    Design (me) returns ConfigurationDesignItem from StepRepr;
	---Purpose: Returns field Design
    SetDesign (me: mutable; Design: ConfigurationDesignItem from StepRepr);
	---Purpose: Set field Design

fields
    theConfiguration: ConfigurationItem from StepRepr;
    theDesign: ConfigurationDesignItem from StepRepr;

end ConfigurationDesign;
