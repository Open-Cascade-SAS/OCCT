-- Created by: Peter KURNEV
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ShrunkRange from IntTools 

 ---Purpose:  
 ---  The class provides the computation of 
 ---  a working (shrunk) range [t1, t2] for 
     ---  the 3D-curve of the edge. 
  
uses
    Box from Bnd, 
    Edge from TopoDS, 
    Vertex from TopoDS, 
    Context  from IntTools

--raises

is 
    Create 
        returns ShrunkRange from IntTools;
    ---C++: alias "Standard_EXPORT virtual ~IntTools_ShrunkRange();"  
    
    SetData (me:out; 
            aE  : Edge from TopoDS;  
            aT1 : Real from Standard;              
            aT2 : Real from Standard;     
            aV1 : Vertex from TopoDS;              
            aV2 : Vertex from TopoDS); 
     
    SetContext(me:out; 
            aCtx: Context from IntTools);  
             
    Context(me) 
        returns Context from IntTools;       
    ---C++: return const &  
    
    SetShrunkRange(me:out; 
         aT1 : Real from Standard;   
         aT2 : Real from Standard);   

    ShrunkRange(me; 
         aT1 :out Real from Standard;   
         aT2 :out Real from Standard); 
  
    BndBox  (me) 
     returns Box from Bnd; 
    ---C++: return const & 
     
    Edge  (me) 
     returns Edge from TopoDS; 
    ---C++: return const &  
      
    Perform(me:out); 
  
    ErrorStatus(me) 
     returns Integer from Standard;  
 ---Purpose:
 --- Returns code of computing shrunk range
 --- completion
 --- 0 - means successful completion
 --- 1 - nothing has been done
 --- 2 - initial range is out of edge's range
 --- 3 - first boundary of initial range is more than
 ---     last boundary
 --- 4 - projection of first vertex failed
 --- 5 - projection of second vertex failed
 --- 6 - shrunk range can not be computed
 ---     shrunk range is setted to initial range
 ---

fields
    myEdge        : Edge from TopoDS is protected; 
    myV1          : Vertex from TopoDS is protected;
    myV2          : Vertex from TopoDS is protected;  
    myT1          : Real from Standard is protected;     
    myT2          : Real from Standard is protected;     
    myTS1         : Real from Standard is protected;     
    myTS2         : Real from Standard is protected;     
    myBndBox      : Box from Bnd is protected;  
    myCtx         : Context from IntTools is protected;
    myErrorStatus : Integer from Standard is protected;   
     
end ShrunkRange;
