-- Created on: 1995-03-08
-- Created by: Laurent BUCHARD
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Class2d from CSLib

uses 
    Pnt2d          from gp,
    Array1OfPnt2d  from TColgp
    
is 

    Create(TP: Array1OfPnt2d from TColgp; aTolu,aTolv:Real from Standard;
           umin,vmin,umax,vmax: Real from Standard)
    returns Class2d     from CSLib;
    
    SiDans(me; P: Pnt2d from gp)
    returns Integer from Standard;
    
    SiDans_OnMode(me; P: Pnt2d from gp; Tol: Real from Standard)
    returns Integer from Standard;
    
    InternalSiDans(me; X,Y: Real from Standard)
    returns Integer from Standard;
    
    InternalSiDansOuOn(me; X,Y: Real from Standard)
    returns Integer from Standard;    

    Copy(me; Other: Class2d from CSLib)
    returns Class2d from CSLib;
    	---C++: return const &
      	---C++: alias operator=
     --Purpose *** Raise if called ***

    Destroy(me: in out);
       	---C++: alias ~
     
    
fields 
    MyPnts2dX: Address  from Standard;
    MyPnts2dY: Address  from Standard;
    Tolu     : Real     from Standard;
    Tolv     : Real     from Standard;
    N        : Integer  from Standard;
    Umin     : Real     from Standard;
    Vmin     : Real     from Standard;
    Umax     : Real     from Standard;
    Vmax     : Real     from Standard;
   
end Class2d from CSLib;


    
    
