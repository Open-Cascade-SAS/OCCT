-- File:	RWStepDimTol_RWGeometricToleranceWithDatumReference.cdl
-- Created:	Wed Jun  4 13:34:35 2003 
-- Author:	Galina KULIKOVA
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWGeometricToleranceWithDatumReference from RWStepDimTol

    ---Purpose: Read & Write tool for GeometricToleranceWithDatumReference

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    GeometricToleranceWithDatumReference from StepDimTol

is
    Create returns RWGeometricToleranceWithDatumReference from RWStepDimTol;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : GeometricToleranceWithDatumReference from StepDimTol);
	---Purpose: Reads GeometricToleranceWithDatumReference

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: GeometricToleranceWithDatumReference from StepDimTol);
	---Purpose: Writes GeometricToleranceWithDatumReference

    Share (me; ent : GeometricToleranceWithDatumReference from StepDimTol;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWGeometricToleranceWithDatumReference;
