-- Created on: 1994-02-14
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

generic class ZerCOnSSParFunc from IntImp 
    (ThePSurface     as any;
     ThePSurfaceTool as any;   --as PSurfaceTool from IntImp(ThePSurface)
     TheCurveOnSurf  as any;
     TheCurveTool    as any     --as COnSCurveTool from IntImp(TheCurve)
    )
    
inherits FunctionSetWithDerivatives from math

      	---Purpose: this function is associated to the intersection between 
      	--          a curve on surface and a surface  .


uses Vector from math,
     Matrix from math,
     Pnt from gp

is
    Create( S1 : ThePSurface;
    	    C  : TheCurveOnSurf;
            S2 : ThePSurface )

	---Purpose: S1 is the surface on which the intersection is searched.
	--          C is a curve on the surface S2.

    	returns ZerCOnSSParFunc from IntImp;
	    

    NbVariables(me) returns Integer from Standard
    is static;
    
    NbEquations(me) returns Integer from Standard
    is static;
    
    Value(me : in out; X : in Vector from math;
    	    	       F : out Vector from math)
    returns Boolean from Standard
    is static;
    
    Derivatives(me : in out;X : in  Vector from math;
    	    	    	    D : out Matrix from math)
    returns Boolean from Standard
    is static;
    
    Values(me : in out;
    	   X  : in Vector from math;
	   F  : out Vector from math; D: out Matrix from math)
    returns Boolean from Standard
    is static;

    Point(me)
    	---C++: return const&
    	returns Pnt from gp
    	is static;
    
    Root(me) returns Real from Standard
    is static;
    
    AuxillarSurface(me)
    	---C++: return const&
    	returns ThePSurface
    	is static;

    AuxillarCurve(me)
    	---C++: return const&
    	returns TheCurveOnSurf
    	is static;
    
fields
     curve    : Address from Standard; --- TheCurveOnSurf;
     surface1 : Address from Standard; --- ThePSurface;
     surface2 : Address from Standard; --- ThePSurface;
     p	      : Pnt from gp;
     f        : Real from Standard;
     
end ZerCOnSSParFunc;
