-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

---Version: 

--  Version	Date         Purpose
--              01/04/93     Creation

class HashAsciiString from PColStd 

---Purpose: Redefines the HashCode for HAsciiString

inherits HOfAsciiString from PColStd

uses

    HAsciiString  from PCollection
    
is

    Create returns HashAsciiString;
    ---Purpose : Empty constructor.

    HashCode (me; MyKey : HAsciiString ; Upper : Integer) 
             returns Integer is redefined;
    ---Purpose : Returns a hashcod value of key bounded by Upper.

    Compare (me; One , Two : HAsciiString) returns Boolean is redefined;
    ---Purpose : Compare two keys and returns a boolean value

end HashAsciiString;

