-- File:        PreDefinedItem.cdl
-- Created:     Mon Dec  4 12:02:29 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWPreDefinedItem from RWStepVisual

	---Purpose : Read & Write Module for PreDefinedItem

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     PreDefinedItem from StepVisual

is

	Create returns RWPreDefinedItem;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable PreDefinedItem from StepVisual);

	WriteStep (me; SW : in out StepWriter; ent : PreDefinedItem from StepVisual);

end RWPreDefinedItem;
