-- Created on: 1992-03-12
-- Created by: Christophe MARION
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

--        <cma@sdsun2> copie quasi exacte de HLRAlgo_Projector

class Projector from Select3D inherits Transient from Standard
    ---Purpose: A framework to define 3D projectors.
    -- Projector provides services for projecting points from
    -- world-coordinates to a viewing plane. Projection could be defined by
    -- corresponding transformation, or coordinate system. The transformation
    -- could be constructed for a view with transposed view transformation
    -- matrix ( that represents view-orientation ), including, for perspective
    -- view, focal distance ( distance from an eye to the view plane ) and
    -- translational part that represents translation of focal point in
    -- view-coordinate space. The Select3D_Projector class recognizes the
    -- predefined set of popular projections: axonometric, top view, front
    -- view and uses more efficient algorithm for projection computations.
    -- User-defined transformation could be also defined in constructor.
    -- Perspective projection consists of two separate parts, that are
    -- composed together during computation: transformation component and
    -- focale distance.

uses
    Real    from Standard,
    Boolean from Standard,
    Trsf    from gp,
    GTrsf   from gp,
    Lin     from gp,
    Pnt     from gp,
    Vec     from gp,
    Ax2     from gp,
    Vec2d   from gp,
    Pnt2d   from gp,
    Box     from Bnd,
    View    from V3d,
    Mat4    from Graphic3d,
    Mat4d   from Graphic3d

raises
    NoSuchObject from Standard

is

    Create (theView : View from V3d) returns Projector from Select3D;
    --- Purpose: Constructs the 3D projector object from the passed view.
    -- The projector captures current model-view and projection transformation
    -- of the passed view.

    Create returns Projector from Select3D;
    --- Purpose: Constructs identity projector.

    Create (theCS : Ax2 from gp)
    ---Purpose: Builds the Projector from the model-view transformation specified
    -- by the passed viewing coordinate system <theCS>. The Projector has
    -- identity projection transformation, is orthogonal.
    -- The viewing coordinate system could be constructed from x direction,
    -- view plane normal direction, and view point location in
    -- world-coordinate space.
    returns Projector from Select3D;

    Create (theCS    : Ax2  from gp;
            theFocus : Real from Standard)
    ---Purpose: Builds the Projector from the model-view transformation specified
    -- by the passed view coordinate system <theCS> and simplified perspective
    -- projection transformation defined by <theFocus> parameter.
    -- The viewing coordinate system could be constructed from x direction,
    -- view plane normal direction, and focal point location in world-coordinate
    -- space. <theFocus> should represent distance of an eye from view plane
    -- in world-coordinate space (focal distance).
    returns Projector from Select3D;

    Create (theViewTrsf : Trsf    from gp;
            theIsPersp  : Boolean from Standard;
            theFocus    : Real    from Standard)
    ---Purpose: Build the Projector from the model-view transformation passed
    -- as <theViewTrsf> and simplified perspective projection transformation
    -- parameters passed as <theIsPersp> and <theFocus>.
    -- In case, when <theViewTrsf> transformation should represent custom view
    -- projection, it could be constructed from two separate components:
    -- transposed view orientation matrix and translation of focal point
    -- in view-coordinate system.
    -- <theViewTrsf> could be built up from x direction, up direction,
    -- view plane normal direction vectors and translation with SetValues(...)
    -- method, where first row arguments (a11, a12, a13, a14)  are x, y, z
    -- component of x direction vector, and x value of reversed translation
    -- vector. Second row arguments, are x y z for up direction and y value of
    -- reversed translation, and the third row defined in the same manner.
    -- This also suits for simple perspective view, where <theFocus> is the focale
    -- distance of an eye from view plane in world-space coordinates.
    -- Note, that in that case amount of perspective distortion (perspective
    -- angle) should be defined through focal distance.
    returns Projector from Select3D;

    Create (theViewTrsf : GTrsf   from gp;
            theIsPersp  : Boolean from Standard;
            theFocus    : Real    from Standard)
    ---Purpose: Builds the Projector from the model-view transformation passed
    -- as <theViewTrsf> and projection transformation for <theIsPersp> and
    -- <theFocus> parameters.
    -- In case, when <theViewTrsf> transformation should represent custom view
    -- projection, it could be constructed from two separate components:
    -- transposed view orientation matrix and translation of a focal point
    -- in view-coordinate system.
    -- This also suits for perspective view, with <theFocus> that could be
    -- equal to distance from an eye to a view plane in 
    -- world-coordinates (focal distance).
    -- The 3x3 transformation matrix is built up from three vectors:
    -- x direction, up direction and view plane normal vectors, where each
    -- vector is a matrix row. Then <theViewTrsf> is constructed from matrix and
    -- reversed translation with methods SetTranslationPart(..) and
    -- SetVectorialPart(..).
    -- Note, that in that case amount of perspective distortion (perspective
    -- angle) should be defined through focal distance.
    returns Projector from Select3D;

    Create (theViewTrsf : Mat4d from Graphic3d;
            theProjTrsf : Mat4d from Graphic3d)
    ---Purpose: Builds the Projector from the passed model-view <theViewTrsf>
    -- and projection <theProjTrsf> transformation matrices.
    returns Projector from Select3D;

    Set (me : mutable;
         theViewTrsf : Trsf    from gp;
         theIsPersp  : Boolean from Standard;
         theFocus    : Real    from Standard);
    ---Purpose: Sets new parameters for the Projector.

    Set (me : mutable;
         theViewTrsf : Mat4d from Graphic3d;
         theProjTrsf : Mat4d from Graphic3d);
    ---Purpose: Sets new parameters for the Projector.

    SetView (me : mutable;
             theView : View from V3d);
    ---Purpose: Sets new parameters for the Projector
    -- captured from the passed view.

    Scaled (me : mutable; theToCheckOptimized : Boolean from Standard = Standard_False)
    ---Purpose: Pre-compute inverse transformation and ensure whether it is possible
    -- to use optimized transformation for the common view-orientation type or not
    -- if <theToCheckOptimized> is TRUE.
    is virtual;

    Perspective (me) returns Boolean
    ---Purpose: Returns True if there is simplified perspective
    -- projection approach is used. Distortion defined by Focus.
    ---C++: inline
    is virtual;

    Focus (me) returns Real from Standard
    ---Purpose: Returns the focal length of simplified perspective
    -- projection approach. Raises program error exception if the
    -- the projection transformation is not specified as simplified
    -- Perspective (for example, custom projection transformation is defined
    -- or the orthogonal Projector is defined).
    ---C++: inline
    is virtual;

    Projection (me) returns Mat4d from Graphic3d;
    ---Purpose: Returns projection transformation. Please note that for
    -- simplified perspective projection approach, defined by Focus, the
    -- returned transformation is identity.
    ---C++: inline
    ---C++: return const &

    Transformation (me) returns GTrsf from gp
    ---Purpose: Returns the view transformation.
    ---C++: inline
    ---C++: return const &
    is virtual;

    InvertedTransformation (me) returns GTrsf from gp
    ---Purpose: Returns the inverted view transformation.
    ---C++: inline
    ---C++: return const &
    is virtual;

    FullTransformation (me) returns Trsf from gp
    ---Purpose: Returns the uniform-scaled view transformation.
    ---C++: inline
    ---C++: return const &
    is virtual;

    Transform (me; theD : in out Vec from gp)
    ---Purpose: Transforms the vector into view-coordinate space.
    ---C++: inline
    is virtual;

    Transform (me; thePnt : in out Pnt from gp)
    ---Purpose: Transforms the point into view-coordinate space.
    ---C++: inline
    is virtual;

    Project (me; theP : Pnt from gp; thePout : out Pnt2d from gp)
    ---Purpose: Transforms the point into view-coordinate space
    -- and applies projection transformation.
    is virtual;

    Project (me; theP : Pnt  from gp; theX, theY, theZ : out Real from Standard)
    ---Purpose: Transforms the point into view-coordinate space
    -- and applies projection transformation.
    is static;

    Project (me; theP     : Pnt   from gp;
                 theD1    : Vec from gp;
                 thePout  : out Pnt2d from gp;
                 theD1out : out Vec2d from gp)
    ---Purpose: Transforms the point and vector passed from its location
    -- into view-coordinate space and applies projection transformation.
    is virtual;

    Shoot (me; theX, theY : Real from Standard) returns Lin from gp
    ---Purpose: Return projection line going through the 2d point <theX, theY>
    is virtual;

    Transform(me; thePnt  : in out Pnt from gp;
                  theTrsf : GTrsf from gp)
    ---C++: inline
    is virtual;

    Transform(me; theLin : in out Lin from gp;
                  theTrsf : GTrsf from gp)
    ---C++: inline
    is virtual;

fields

    myType       : Integer from Standard;
    myPersp      : Boolean from Standard is protected;
    myFocus      : Real    from Standard is protected;
    myGTrsf      : GTrsf   from gp is protected;
    myInvTrsf    : GTrsf   from gp is protected;
    myScaledTrsf : Trsf    from gp is protected;
    myProjTrsf   : Mat4d   from Graphic3d is protected;

end Projector;
