-- File:        LengthMeasureWithUnit.cdl
-- Created:     Mon Dec  4 12:02:27 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWLengthMeasureWithUnit from RWStepBasic

	---Purpose : Read & Write Module for LengthMeasureWithUnit

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     LengthMeasureWithUnit from StepBasic,
     EntityIterator from Interface

is

	Create returns RWLengthMeasureWithUnit;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable LengthMeasureWithUnit from StepBasic);

	WriteStep (me; SW : in out StepWriter; ent : LengthMeasureWithUnit from StepBasic);

	Share(me; ent : LengthMeasureWithUnit from StepBasic; iter : in out EntityIterator);

end RWLengthMeasureWithUnit;
