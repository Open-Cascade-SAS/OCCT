-- File:	IGESGeom_ToolSplineSurface.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolSplineSurface  from IGESGeom

    ---Purpose : Tool to work on a SplineSurface. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses SplineSurface from IGESGeom,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolSplineSurface;
    ---Purpose : Returns a ToolSplineSurface, ready to work


    ReadOwnParams (me; ent : mutable SplineSurface;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : SplineSurface;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : SplineSurface;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a SplineSurface <ent>, from
    --           its specific (own) parameters

    DirChecker (me; ent : SplineSurface) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : SplineSurface;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : SplineSurface; entto : mutable SplineSurface;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : SplineSurface;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolSplineSurface;
