-- Created on: 1992-08-18
-- Created by: Modelistation
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




private class Parameter from Hatch

	---Purpose: Stores an intersection on a line represented by :
	--          
	--          * A Real parameter.
	--          
	--          * A flag True when the parameter starts an interval.
	--          

uses
    Real    from Standard,
    Integer from Standard,
    Boolean from Standard

is
    Create;
    
    Create( Par1  : Real    from Standard;
            Start : Boolean from Standard;
	    Index : Integer from Standard = 0;
	    Par2  : Real    from Standard = 0)
    returns Parameter from Hatch;
    
fields
    myPar1  : Real      from Standard;
    myStart : Boolean   from Standard;
    myIndex : Integer   from Standard;
    myPar2  : Real      from Standard;
    
friends
    class Line    from Hatch,
    class Hatcher from Hatch

end Parameter;
