-- Created on: 1993-07-07
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class ShapeScanner from TopOpeBRep
    
    ---Purpose: Find, among the  subshapes SS of a reference shape
    --          RS, the ones which 3D box interfers with the box of
    --          a shape S (SS and S are of the same type).

uses

    ShapeEnum from TopAbs,
    Shape from TopoDS,
    ListIteratorOfListOfInteger from TColStd,
    ShapeExplorer from TopOpeBRepTool,
    BoxSort from TopOpeBRepTool

is

    Create returns ShapeScanner from TopOpeBRep;
    Clear(me:in out);
    AddBoxesMakeCOB(me:in out;S:Shape;TS:ShapeEnum;TA:ShapeEnum=TopAbs_SHAPE);
    Init(me:in out;E:Shape);
    Init(me:in out;X:in out ShapeExplorer from TopOpeBRepTool);
    More(me) returns Boolean;
    Next(me:in out);
    Current(me) returns Shape;---C++: return const &
    BoxSort(me) returns BoxSort from TopOpeBRepTool;---C++:return const &
    ChangeBoxSort(me:in out) returns BoxSort from TopOpeBRepTool;---C++:return &
    Index(me) returns Integer;
    DumpCurrent(me; OS:in out OStream) returns OStream;---C++: return &
    
fields

    myBoxSort:BoxSort from TopOpeBRepTool;
    myListIterator:ListIteratorOfListOfInteger from TColStd;
    
end ShapeScanner from TopOpeBRep;

