-- File:        IntersectionCurve.cdl
-- Created:     Mon Dec  4 12:02:27 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWIntersectionCurve from RWStepGeom

	---Purpose : Read & Write Module for IntersectionCurve

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     IntersectionCurve from StepGeom,
     EntityIterator from Interface

is

	Create returns RWIntersectionCurve;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable IntersectionCurve from StepGeom);

	WriteStep (me; SW : in out StepWriter; ent : IntersectionCurve from StepGeom);

	Share(me; ent : IntersectionCurve from StepGeom; iter : in out EntityIterator);

end RWIntersectionCurve;
