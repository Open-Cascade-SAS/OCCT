-- File:	BRepFilletAPI_MakeFillet2d.cdl
-- Created:	Thu Aug 31 14:18:16 1995
-- Author:	Remi LEQUETTE
--		<rle@mentox>
---Copyright:	 Matra Datavision 1995



class MakeFillet2d from BRepFilletAPI inherits MakeShape from BRepBuilderAPI

	---Purpose: Describes functions to build fillets and chamfers on the
    	-- vertices of a planar face.
    	-- Fillets and Chamfers on the Vertices of a Planar Face
    	-- A MakeFillet2d object provides a framework for:
    	-- - initializing the construction algorithm with a given face,
    	-- - acquiring the data characterizing the fillets and chamfers,
    	-- -   building the fillets and chamfers, and constructing the
    	--   resulting shape, and
    	-- -   consulting the result.
    	-- Warning
    	-- Only segments of straight lines and arcs of circles are
    	-- treated. BSplines are not processed.
        
uses
    Builder           from ChFi2d,
    ConstructionError from ChFi2d,
    Face              from TopoDS,
    Edge              from TopoDS,
    Vertex            from TopoDS,
    Shape             from TopoDS,
    ShapeModification from BRepBuilderAPI,
    SequenceOfShape   from TopTools,
    ListOfShape       from TopTools

is


    Create returns MakeFillet2d from BRepFilletAPI;
    	---Purpose: Initializes an empty algorithm for computing fillets and
    	--   chamfers. The face on which the fillets and
    	--   chamfers are built is defined using the Init function.
    	-- The vertices on which fillets or chamfers are built are
    	-- defined using the AddFillet or AddChamfer function.
    	-- Warning
    	-- The status of the initialization, as given by the Status
    	-- function, can be one of the following:
    	-- -   ChFi2d_Ready if the initialization is correct,
    	-- -   ChFi2d_NotPlanar if F is not planar,
    	-- -   ChFi2d_NoFace if F is a null face.
        
    Create ( F : Face ) returns MakeFillet2d from BRepFilletAPI;
    	---Purpose: Initializes an algorithm for computing fillets and chamfers on the face F.
    	-- The vertices on which fillets or chamfers are built are
    	-- defined using the AddFillet or AddChamfer function.
    	-- Warning
    	-- The status of the initialization, as given by the Status
    	-- function, can be one of the following:
    	-- -   ChFi2d_Ready if the initialization is correct,
    	-- -   ChFi2d_NotPlanar if F is not planar,
    	-- -   ChFi2d_NoFace if F is a null face.    

    
    Init( me : in out; F : Face );
    	---Purpose: Initializes this algorithm for constructing fillets or
    	-- chamfers with the face F.
    	-- Warning
    	-- The status of the initialization, as given by the Status
    	-- function, can be one of the following:
    	-- -   ChFi2d_Ready if the initialization is correct,
    	-- -   ChFi2d_NotPlanar if F is not planar,
    	-- -   ChFi2d_NoFace if F is a null face.

    Init( me : in out; RefFace, ModFace : Face );
    	---Purpose: This initialize  method allow  to init the builder
    	--          from a  face <RefFace> and  another face <ModFace>
    	--          which derive from  <RefFace>.  This  is usefull to
    	--          modify a fillet or   a chamfer already created  on
    	--          <ModFace> .
    

    AddFillet ( me : in out; V : Vertex; Radius : Real ) returns Edge;
    	---Purpose: Adds a fillet of radius Radius between the two edges
    	-- adjacent to the vertex V on the face modified by this
    	-- algorithm. The two edges do not need to be rectilinear.
    	-- This function returns the fillet and builds the resulting face.
    	-- Warning
    	-- The status of the construction, as given by the Status
    	-- function, can be one of the following:
    	-- - ChFi2d_IsDone if the fillet is built,
    	-- - ChFi2d_ConnexionError if V does not belong to the initial face,
    	-- -   ChFi2d_ComputationError if Radius is too large
    	--   to build a fillet between the two adjacent edges,
    	-- -   ChFi2d_NotAuthorized
    	-- -   if one of the two edges connected to V is a fillet or chamfer, or
    	-- -   if a curve other than a straight line or an arc of a
    	--    circle is used as E, E1 or E2.
    	-- Do not use the returned fillet if the status of the construction is not ChFi2d_IsDone.
    	-- Exceptions
    	-- Standard_NegativeValue if Radius is less than or equal to zero. 


    ModifyFillet ( me : in out; Fillet : Edge; Radius : Real) 
    returns Edge;
    	---Purpose: Assigns the radius Radius to the fillet Fillet already
    	-- built on the face modified by this algorithm.
    	-- This function returns the new fillet and modifies the existing face.
    	-- Warning
    	-- The status of the construction, as given by the Status
    	-- function, can be one of the following:
    	-- -   ChFi2d_IsDone if the new fillet is built,
    	-- -   ChFi2d_ConnexionError if Fillet does not
    	--   belong to the existing face,
    	-- -   ChFi2d_ComputationError if Radius is too
    	--  large to build a fillet between the two adjacent edges.
    	--   Do not use the returned fillet if the status of the
    	-- construction is not ChFi2d_IsDone.
    	-- Exceptions
    	-- Standard_NegativeValue if Radius is less than or equal to zero.    

    RemoveFillet( me : in out; Fillet : Edge)
    returns Vertex;
    	---Purpose: Removes the fillet Fillet already built on the face
    	-- modified by this algorithm.
    	-- This function returns the vertex connecting the two
    	-- adjacent edges of Fillet and modifies the existing face.
    	-- Warning
    	-- -   The returned vertex is only valid if the Status
    	--   function returns ChFi2d_IsDone.
    	-- -   A null vertex is returned if the edge Fillet does not
    	--   belong to the initial face.
  
    
    AddChamfer ( me : in out; E1, E2 : Edge; D1, D2 : Real ) 
    returns Edge;
    	---Purpose: Adds a chamfer on the face modified by this algorithm
    	--    between the two adjacent edges E1 and E2, where
    	--   the extremities of the chamfer are on E1 and E2 at
    	--   distances D1 and D2 respectively
    	--    In cases where the edges are not rectilinear, distances
    	-- are measured using the curvilinear abscissa of the
    	-- edges and the angle is measured with respect to the
    	-- tangent at the corresponding point.
    	-- The angle Ang is given in radians.
    	-- This function returns the chamfer and builds the resulting face.

    AddChamfer ( me : in out; E : Edge; V : Vertex; D, Ang  : Real ) 
    returns Edge;
    	---Purpose: Adds a chamfer on the face modified by this algorithm
    	--   between the two edges connected by the vertex V,
    	--   where E is one of the two edges. The chamfer makes
    	--   an angle Ang with E and one of its extremities is on
    	--   E at distance D from V.
    	--    In cases where the edges are not rectilinear, distances
    	-- are measured using the curvilinear abscissa of the
    	-- edges and the angle is measured with respect to the
    	-- tangent at the corresponding point.
    	-- The angle Ang is given in radians.
    	-- This function returns the chamfer and builds the resulting face. 
    	-- Warning
    	-- The status of the construction, as given by the Status function, can
    	-- be one of the following:
    	-- -          ChFi2d_IsDone if the chamfer is built,
    	-- -  ChFi2d_ParametersError if D1, D2, D or Ang is less than or equal to zero,
    	-- -          ChFi2d_ConnexionError if:
    	-- - the edge E, E1 or E2 does not belong to the initial face, or
    	-- -  the edges E1 and E2 are not adjacent, or
    	-- -  the vertex V is not one of the limit points of the edge E,
    	-- -          ChFi2d_ComputationError if the parameters of the chamfer
    	--   are too large to build a chamfer between the two adjacent edges,
    	-- -          ChFi2d_NotAuthorized if:
    	-- - the edge E1, E2 or one of the two edges connected to V is a fillet or chamfer, or
    	-- - a curve other than a straight line or an arc of a circle is used as E, E1 or E2.
    	-- Do not use the returned chamfer if
    	-- the status of the construction is not ChFi2d_IsDone.
        
    ModifyChamfer ( me : in out; Chamfer : Edge;
    	    	    E1 : Edge; E2 : Edge; D1, D2 : Real)
    returns  Edge;
    	---Purpose: Modifies the chamfer Chamfer on the face modified
    	-- by this algorithm, where:
    	--   E1 and E2 are the two adjacent edges on which
    	--   Chamfer is already built; the extremities of the new
    	--   chamfer are on E1 and E2 at distances D1 and D2 respectively.
        
    
    ModifyChamfer ( me : in out; Chamfer, E : Edge; D, Ang : Real)
    returns  Edge;
    	---Purpose: Modifies the chamfer Chamfer on the face modified
    	-- by this algorithm, where:
    	--   E is one of the two adjacent edges on which
    	--   Chamfer is already built; the new chamfer makes
    	--   an angle Ang with E and one of its extremities is
    	-- on E at distance D from the vertex on which the chamfer is built.
    	--   In cases where the edges are not rectilinear, the
    	-- distances are measured using the curvilinear abscissa
    	-- of the edges and the angle is measured with respect
    	-- to the tangent at the corresponding point.
    	-- The angle Ang is given in radians.
    	-- This function returns the new chamfer and modifies the existing face.
    	-- Warning
    	-- The status of the construction, as given by the Status
    	-- function, can be one of the following:
    	-- -   ChFi2d_IsDone if the chamfer is built,
    	-- -   ChFi2d_ParametersError if D1, D2, D or Ang is less than or equal to zero,
    	-- -   ChFi2d_ConnexionError if:
    	--   -   the edge E, E1, E2 or Chamfer does not belong
    	--    to the existing face, or
    	--   -   the edges E1 and E2 are not adjacent,
    	-- -   ChFi2d_ComputationError if the parameters of
    	--   the chamfer are too large to build a chamfer
    	--   between the two adjacent edges,
    	-- -   ChFi2d_NotAuthorized if E1 or E2 is a fillet or chamfer.
    	-- Do not use the returned chamfer if the status of the
    	-- construction is not ChFi2d_IsDone. 

    RemoveChamfer( me : in out; Chamfer : Edge)
    returns Vertex;
    	---Purpose: Removes the chamfer Chamfer already built on the face
    	-- modified by this algorithm.
    	-- This function returns the vertex connecting the two
    	-- adjacent edges of Chamfer and modifies the existing face.
    	-- Warning
    	-- -   The returned vertex is only valid if the Status
    	--   function returns ChFi2d_IsDone.
    	-- -   A null vertex is returned if the edge Chamfer does
    	--   not belong to the initial face.

    ----------------------------------------------
    -- Results
    ----------------------------------------------
 
    IsModified( me; E : Edge ) returns Boolean;
    	---Purpose:    Returns true if the edge E on the face modified by this
    	-- algorithm is chamfered or filleted.
    	-- Warning
    	-- Returns false if E does not belong to the face modified by this algorithm.
    	---C++:     inline 


    FilletEdges( me ) returns SequenceOfShape; 
    	---Purpose: Returns the table of fillets on the face modified by this algorithm.
    	---C++:     return const &
    	---C++:     inline 
	
    NbFillet( me ) returns Integer;
    	---Purpose: Returns the number of fillets on the face modified by this algorithm.
    	---C++: inline 


    ChamferEdges( me ) returns SequenceOfShape; 
    	---Purpose: Returns the table of chamfers on the face modified by this algorithm.
    	---C++:     return const &
    	---C++:     inline 
	
    NbChamfer( me ) returns Integer;
    	---Purpose: Returns the number of chamfers on the face modified by this algorithm.
    	---C++: inline 

    -------------------------------------------
    -- Methods usefull for historical utilities --
    -------------------------------------------
 
    Modified (me: in out; S : Shape from TopoDS)
    	---Purpose: Returns the list  of shapes modified from the shape
    	--          <S>. 
        ---C++: return const & 
        ---Level: Public
    returns ListOfShape from TopTools
    is redefined virtual;

    NbCurves(me)
    	---Purpose: returns the number of new curves
    	--          after the shape creation.
	---Level: Public
    returns Integer from Standard;



    NewEdges(me: in out; I: Integer from Standard) 
    	---Purpose: Return the Edges created for curve I.
    	---C++:     return const &
	---Level: Public
    returns ListOfShape from TopTools;



    HasDescendant( me; E : Edge) returns Boolean;
    	---C++: inline 
    
    
    DescendantEdge( me; E : Edge) returns Edge;
    	---Purpose: Returns the chamfered or filleted edge built from the
    	-- edge E on the face modified by this algorithm. If E has
    	-- not been modified, this function returns E.
    	-- Exceptions
    	-- Standard_NoSuchObject if the edge E does not
    	-- belong to the initial face.
    	---C++:     return const &
    	---C++:     inline 


    BasisEdge( me; E : Edge) returns Edge;
    	---Purpose: Returns the basis edge on the face modified by this
    	-- algorithm from which the chamfered or filleted edge E is
    	-- built. If E has not been modified, this function returns E.
    	-- Warning
    	-- E is returned if it does not belong to the initial face.
      	---C++:     return const &

    Status(me) returns ConstructionError from ChFi2d;
    	---C++:     inline


    Build(me : in out)
	---Purpose: Update the result and set the Done flag
	---Level: Public
    is redefined;
	

fields

    myMakeChFi2d : Builder from ChFi2d;
    
end MakeFillet2d;
