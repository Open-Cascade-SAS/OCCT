-- Created on: 1992-01-21
-- Created by: GG
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class OrthographicView from V3d

        ---Version:

	---Purpose: Define an orthographic view.
        --          See the methods of the Class View

        ---Keywords: View,Orthographic

        ---Warning:

        ---References:


inherits View from V3d

uses

	Viewer from V3d,
	PerspectiveView from V3d

is

    	Create ( VM : mutable Viewer ) returns mutable OrthographicView; 
	---Level : Public
	---Purpose: Define an orthographic view in the viewer VM.

    	Create ( VM : mutable Viewer ; V : PerspectiveView ) 
					returns mutable OrthographicView; 
	---Level : Public
	---Purpose: Defines an orthographic view from a Perspective view.
	--	    The parameters of the original view are duplicated
	--	    in the resulting view (Projection,Mapping,Context) .
	--	    The view thus created must be activated in a new
	--	    window.

    	Create ( VM : mutable Viewer ; V : OrthographicView ) 
					returns mutable OrthographicView; 
	---Level : Public
	---Purpose: Defines one orthographic view from another.
	--	    The parameters of the original view are duplicated 
	--	    in the resulting view. (Projection,Mapping,Context) .
	--	    The view thus created must be activated in a new window.

        Copy ( me ) returns mutable OrthographicView from V3d is static;
	---Level : Public
end OrthographicView;
