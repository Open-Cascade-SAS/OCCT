-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PresentationSize from StepVisual 

inherits TShared from MMgt

uses

	PresentationSizeAssignmentSelect from StepVisual, 
	PlanarBox from StepVisual
is

	Create returns mutable PresentationSize;
	---Purpose: Returns a PresentationSize

	Init (me : mutable;
	      aUnit : PresentationSizeAssignmentSelect from StepVisual;
	      aSize : mutable PlanarBox from StepVisual) is virtual;

	-- Specific Methods for Field Data Access --

	SetUnit(me : mutable; aUnit : PresentationSizeAssignmentSelect);
	Unit (me) returns PresentationSizeAssignmentSelect;
	SetSize(me : mutable; aSize : mutable PlanarBox);
	Size (me) returns mutable PlanarBox;

fields

	unit : PresentationSizeAssignmentSelect from StepVisual; -- a SelectType
	size : PlanarBox from StepVisual;

end PresentationSize;
