-- Created by: Peter KURNEV
-- Copyright (c) 2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class BuilderAlgo from BRepAlgoAPI
        inherits Algo from BRepAlgoAPI
 ---Purpose: provides the root interface for algorithms

uses
    BaseAllocator from BOPCol,
    PPaveFiller from BOPAlgo,
    PBuilder from BOPAlgo

--raises

is
    Initialize
    returns BuilderAlgo from BRepAlgoAPI;
    ---C++: alias "Standard_EXPORT virtual ~BRepAlgoAPI_BuilderAlgo();"

    Initialize (theAllocator: BaseAllocator from BOPCol)
    returns BuilderAlgo from BRepAlgoAPI;

    SetFuzzyValue(me:out; 
        theFuzz : Real from Standard);
    ---Purpose: Sets the additional tolerance

    FuzzyValue(me)
    returns Real from Standard;
    ---Purpose: Returns the additional tolerance 

fields
    myDSFiller   : PPaveFiller from BOPAlgo  is protected;
    myBuilder    : PBuilder    from BOPAlgo  is protected;
    myFuzzyValue : Real        from Standard is protected;

end BuilderAlgo;
