-- File:	RWStepFEA_RWNodeWithSolutionCoordinateSystem.cdl
-- Created:	Thu Dec 12 17:51:07 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWNodeWithSolutionCoordinateSystem from RWStepFEA

    ---Purpose: Read & Write tool for NodeWithSolutionCoordinateSystem

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    NodeWithSolutionCoordinateSystem from StepFEA

is
    Create returns RWNodeWithSolutionCoordinateSystem from RWStepFEA;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : NodeWithSolutionCoordinateSystem from StepFEA);
	---Purpose: Reads NodeWithSolutionCoordinateSystem

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: NodeWithSolutionCoordinateSystem from StepFEA);
	---Purpose: Writes NodeWithSolutionCoordinateSystem

    Share (me; ent : NodeWithSolutionCoordinateSystem from StepFEA;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWNodeWithSolutionCoordinateSystem;
