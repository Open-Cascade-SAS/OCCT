-- Created on: 1993-01-28
-- Created by: Gilles DEBARBOUILLE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class CompiledMethod from Dynamic

inherits

    MethodDefinition from Dynamic
    ---Purpose: A Dynamic_CompiledMethod adds to the definition of the
    --          Dynamic_Method the C++ mangled name of the function to
    --          be  run. An application using  instances of this class
    --          must bind the C++  name of  the  method with the  true
    --          address in the executable.

uses

    CString from Standard,
    HAsciiString from TCollection,
    AsciiString  from TCollection


is

    Create(aname : CString from Standard;
           afunction : CString from Standard) returns mutable CompiledMethod from Dynamic;
    
    ---Level: Advanced 
    
    ---Purpose: Creates  a compiled method   with <aname> as user name
    --          and <afunction> as C++ mangled name.
    
    Function(me : mutable ; afunction : CString from Standard)
    
    ---Level: Advanced 
    
    ---Purpose: Sets the  C++ mangled name  of the method to the field
    --          <thefunction>.
    
    is static;
    
    Function(me) returns AsciiString from TCollection
    
    ---Level: Advanced 
    
    ---Purpose: Returns the C++ mangled name of the function.
    
    is static;
    
fields

    thefunction : HAsciiString from TCollection;

end CompiledMethod;
