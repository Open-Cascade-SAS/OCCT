-- Created on: 2003-09-29
-- Created by: Alexander SOLOVYOV and Sergey LITONIN
-- Copyright (c) 2003-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class DummySensitiveEntity from MeshVS inherits SensitiveEntity from SelectBasics

	---Purpose: This class allows to create owners to all elements or nodes,
        -- both hidden and shown, but these owners user cannot select "by hands"
        -- in viewer. They means for internal application tasks, for example, receiving
        -- all owners, both for hidden and shown entities.
uses
  EntityOwner   from SelectBasics,
  ListOfBox2d   from SelectBasics,

  Array1OfPnt2d from TColgp,

  Box2d         from Bnd

is
   Create   ( OwnerId : EntityOwner from SelectBasics ) returns mutable DummySensitiveEntity from MeshVS;

   Areas    ( me: mutable;
              aresult: in out ListOfBox2d from SelectBasics ) is redefined;

   Matches  ( me: mutable;
              X, Y, aTol: Real;
              DMin: out Real ) returns Boolean is redefined;

   Matches  ( me: mutable;
              XMin, YMin, XMax, YMax, aTol: Real ) returns Boolean is redefined;

   Matches  ( me: mutable;
              Polyline : Array1OfPnt2d from TColgp;
              aBox     : Box2d from Bnd;
              aTol     : Real    ) returns Boolean is redefined;

   Is3D     ( me ) returns Boolean is redefined;

   NeedsConversion ( me ) returns Boolean is redefined;

   MaxBoxes ( me ) returns Integer is redefined;

end DummySensitiveEntity;
