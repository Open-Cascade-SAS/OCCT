-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.





class Cylinder   from gp   inherits Storable

        --- Purpose :
        --  Describes an infinite cylindrical surface.
        -- A cylinder is defined by its radius and positioned in space
        -- with a coordinate system (a gp_Ax3 object), the "main
        -- Axis" of which is the axis of the cylinder. This coordinate
        -- system is the "local coordinate system" of the cylinder.
        -- Note: when a gp_Cylinder cylinder is converted into a
        -- Geom_CylindricalSurface cylinder, some implicit
        -- properties of its local coordinate system are used explicitly:
        -- -   its origin, "X Direction", "Y Direction" and "main
        -- Direction" are used directly to define the parametric
        -- directions on the cylinder and the origin of the parameters,
        -- -   its implicit orientation (right-handed or left-handed)
        --   gives an orientation (direct or indirect) to the
        --   Geom_CylindricalSurface cylinder.
        -- See Also
        -- gce_MakeCylinder which provides functions for more
        -- complex cylinder constructions
        -- Geom_CylindricalSurface which provides additional
        -- functions for constructing cylinders and works, in
        -- particular, with the parametric equations of cylinders gp_Ax3

uses Ax1  from gp,
     Ax2  from gp, 
     Ax3  from gp, 
     Dir  from gp,
     Pnt  from gp,
     Trsf from gp,
     Vec  from gp

raises ConstructionError from Standard

is

 Create   returns Cylinder;
        ---C++: inline
        --- Purpose : Creates a indefinite cylinder.

  Create (A3 : Ax3; Radius : Real)  returns Cylinder
        ---C++: inline
        --- Purpose : Creates a cylinder of radius Radius, whose axis is the "main
        --  Axis" of A3. A3 is the local coordinate system of the cylinder.   Raises ConstructionErrord if R < 0.0
     raises ConstructionError;

  SetAxis (me : in out; A1 : Ax1)
        ---C++: inline
        --- Purpose : Changes the symmetry axis of the cylinder. Raises ConstructionError if the direction of A1 is parallel to the "XDirection"
        --  of the coordinate system of the cylinder.
     raises ConstructionError
 
     is static;

  SetLocation (me : in out; Loc : Pnt)  is static;
        ---C++:inline
        --- Purpose : Changes the location of the surface.

  SetPosition (me : in out; A3 : Ax3)  is static;
       ---C++:inline
       --- Purpose : Change the local coordinate system of the surface.

  SetRadius (me : in out; R : Real)
        ---C++: inline
        ---Purpose: Modifies the radius of this cylinder.
        -- Exceptions
        -- Standard_ConstructionError if R is negative.
     raises ConstructionError
     is static;

  UReverse (me : in out)
        ---C++:inline
	---Purpose: Reverses the   U   parametrization of   the cylinder
	--          reversing the YAxis.
  is static;

  VReverse (me : in out)
        ---C++:inline
	---Purpose: Reverses the   V   parametrization of   the  plane
	--          reversing the Axis.
  is static;

  Direct (me) returns Boolean from Standard
        ---C++: inline
        ---Purpose: Returns true if the local coordinate system of this cylinder is right-handed.
  is static;

  Axis (me)  returns Ax1  is static;
        ---C++: inline
        --- Purpose : Returns the symmetry axis of the cylinder.
    	---C++: return const&

  Coefficients (me; A1, A2, A3, B1, B2, B3, C1, C2, C3, D : out Real)
     is static;
       --- Purpose :
       --  Computes the coefficients of the implicit equation of the quadric
       --  in the absolute cartesian coordinate system :
       --  A1.X**2 + A2.Y**2 + A3.Z**2 + 2.(B1.X.Y + B2.X.Z + B3.Y.Z) +
       --  2.(C1.X + C2.Y + C3.Z) + D = 0.0

  Location (me) returns Pnt  is static;
        ---C++: inline
        --- Purpose :  Returns the "Location" point of the cylinder.
    	---C++: return const&

  Position (me)  returns Ax3  is static;
        --- Purpose :
        --  Returns the local coordinate system of the cylinder.
        ---C++: inline
        ---C++: return const&

  Radius (me)   returns Real   is static;
        ---C++: inline
        --- Purpose : Returns the radius of the cylinder.

  XAxis (me) returns Ax1  is static;
        ---C++: inline
        --- Purpose : Returns the axis X of the cylinder.

  YAxis (me) returns Ax1  is static;
        ---C++: inline
        --- Purpose : Returns the axis Y of the cylinder.





  Mirror (me : in out; P : Pnt)            is static;

  Mirrored (me; P : Pnt)  returns Cylinder is static;

        --- Purpose :
        --  Performs the symmetrical transformation of a cylinder 
        --  with respect to the point P which is the center of the 
        --  symmetry.
                    


  Mirror (me : in out; A1 : Ax1)              is static;

  Mirrored (me; A1 : Ax1)   returns Cylinder  is static;
        --- Purpose :
        --  Performs the symmetrical transformation of a cylinder with
        --  respect to an axis placement which is the axis of the
        --  symmetry.


 

  Mirror (me : in out; A2 : Ax2)               is static;

  Mirrored (me; A2 : Ax2)    returns Cylinder  is static;

        --- Purpose :
        --  Performs the symmetrical transformation of a cylinder with respect 
        --  to a plane. The axis placement A2 locates the plane of the
        --  of the symmetry : (Location, XDirection, YDirection).

  

  Rotate (me : in out; A1 : Ax1; Ang : Real)           is static;
        ---C++: inline
  Rotated (me; A1 : Ax1; Ang : Real) returns Cylinder  is static;
        ---C++: inline
        --- Purpose :
        --  Rotates a cylinder. A1 is the axis of the rotation.
        --  Ang is the angular value of the rotation in radians.


  Scale (me : in out; P : Pnt; S : Real)            is static;
        ---C++: inline
  Scaled (me; P : Pnt; S : Real)  returns Cylinder  is static;
        ---C++: inline
        --- Purpose : 
        --  Scales a cylinder. S is the scaling value.
        --  The absolute value of S is used to scale the cylinder




  Transform (me : in out; T : Trsf)                 is static;
        ---C++: inline
  Transformed (me; T : Trsf)     returns Cylinder   is static;
        ---C++: inline
        --- Purpose :
        --  Transforms a cylinder with the transformation T from class Trsf.


 
  Translate (me : in out; V : Vec)            is static;
        ---C++: inline
  Translated (me; V : Vec)  returns Cylinder  is static;
        ---C++: inline
        --- Purpose :
        --  Translates a cylinder in the direction of the vector V.
        --  The magnitude of the translation is the vector's magnitude.




  Translate (me : in out; P1, P2 : Pnt)            is static; 
        ---C++: inline
  Translated (me; P1, P2 : Pnt)  returns Cylinder  is static;
        ---C++: inline
        --- Purpose :
        --  Translates a cylinder from the point P1 to the point P2.



fields

  pos    : Ax3;
  radius : Real;

end;
