-- Created on: 2002-02-20
-- Created by: Andrey BETENEV
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ProgressScale from Message 

    ---Purpose: Internal data structure for scale in ProgressIndicator
    --
    --          Basically it defines three things:
    --          - name that can be used for generating user messages
    --          - limits and characteristics of the current scale,
    --            along with derived coefficients to map it into basic scale [0-1]
    --          - methods for conversion of values from current scale
    --            to basic one and back
    --
    --          NOTE: There is no special protection against bad input data
    --          like min > max etc. except cases when it can cause exception

uses
    HAsciiString from TCollection
is

    Create returns ProgressScale from Message;
    	---Purpose: Creates scale ranged from 0 to 100 with step 1

    ---Scope: Access to fields

    SetName(me : out; theName : CString);
    	---C++:inline
    SetName(me : out; theName : HAsciiString from TCollection);
    	---C++:inline
    	---Purpose: Sets scale name
    
    GetName(me) returns HAsciiString from TCollection;
    	---C++:inline
    	---Purpose: Gets scale name
	--          Name may be Null handle if not set

    SetMin(me : out; theMin : Real);
    	---C++:inline
    	---Purpose: Sets minimum value of scale
    
    GetMin(me) returns Real;
    	---C++:inline
    	---Purpose: Gets minimum value of scale

    SetMax(me : out; theMax : Real);
    	---C++:inline
    	---Purpose: Sets minimum value of scale
    
    GetMax(me) returns Real;
    	---C++:inline
    	---Purpose: Gets minimum value of scale

    SetRange (me: out; min, max: Real);
    	---C++: inline
    	---Purpose: Set both min and max
	
    SetStep(me : out; theStep : Real);
    	---C++:inline
    	---Purpose: Sets default step
    
    GetStep(me) returns Real;
    	---C++:inline
    	---Purpose: Gets default step

    SetInfinite(me : out; theInfinite : Boolean = Standard_True);
    	---C++:inline
    	---Purpose: Sets flag for infinite scale
    
    GetInfinite(me) returns Boolean;
    	---C++:inline
    	---Purpose: Gets flag for infinite scale

    SetScale (me: out; min, max, step: Real; theInfinite : Boolean = Standard_True);
    	---C++: inline
    	---Purpose: Set all scale parameters
	
    ---Scope: Mapping to base scale
    
    SetSpan (me: out; first, last: Real);
    	---C++: inline
    	---Purpose: Defines span occupied by the scale on the basis scale
	
    GetFirst (me) returns Real;
    	---C++: inline
    GetLast (me) returns Real;
    	---C++: inline
    	---Purpose: Return information on span occupied by the scale on the base scale
	
    LocalToBase (me; val: Real) returns Real;
    BaseToLocal (me; val: Real) returns Real;
    	---Purpose: Convert value from this scale to base one and back

fields
    
    myName: HAsciiString from TCollection; -- name
    
    myMin, myMax: Real;     -- range of a scale
    myStep : Real;          -- default step
    myInfinite: Boolean;    -- flag for infinite scale

    myFirst, myLast : Real; -- span on base scale

end ProgressScale;
