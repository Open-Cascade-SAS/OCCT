-- Created on: 2009-04-06
-- Created by: Sergey ZARITCHNY
-- Copyright (c) 2009-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Plane from TDataXtd inherits Attribute from TDF

    	
	---Purpose: The basis to define a plane attribute.
    	--  Warning:  Use TDataXtd_Geometry  attribute  to retrieve  the
	--          gp_Pln of the Plane attribute

uses Attribute       from TDF,
     Label           from TDF,
     GUID            from Standard,
     Label           from TDF,
     Plane           from Geom,
     Pln             from gp,
     DataSet         from TDF,
     RelocationTable from TDF

is    

    ---Purpose: class methods
    --          =============
   
    GetID (myclass)    
    	---C++: return const & 
    returns GUID from Standard;
    	---Purpose:
    	-- Returns the GUID for plane attributes.

    Set (myclass ; label : Label from TDF)    
    	---Purpose:  Finds or creates the plane attribute defined by
    	-- the label label.
    	-- Warning
    	-- If you are creating the attribute with this syntax, a
    	-- planar face should already be associated with label.
    returns Plane from TDataXtd;    

    Set (myclass ; label : Label from TDF; P : Pln from gp)
    	---Purpose: Finds,  or creates,  a Plane  attribute  and sets <P>  as
    	--          generated the associated NamedShape.
    returns Plane from TDataXtd;    


    ---Purpose: Plane methods
    --         =============    

    Create
    returns mutable Plane from TDataXtd;  
    
    ---Category: TDF_Attribute methods
    --           =====================
    
    ID (me)  
    	---C++: return const & 
    returns GUID from Standard;

    Restore (me: mutable; With : Attribute from TDF);

    NewEmpty (me)
    returns mutable Attribute from TDF;

    Paste (me; Into : mutable Attribute from TDF;
	       RT   : mutable RelocationTable from TDF);  

    Dump (me; anOS : in out OStream from Standard)
    	returns OStream from Standard
    	is redefined;
	---C++: return &

end Plane;


