-- Created on: 1992-05-27
-- Created by: Remi LEQUETTE
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class TVertex from PBRep inherits TVertex from PTopoDS

	---Purpose: The TVertex from  PBRep inherits  from  the TVertex
	--          from TopoDS. 
	--          
	--          The  TVertex contains a Pnt from gp and a tolerance.
	--            
uses
    Pnt from gp,
    PointRepresentation from PBRep

is
    Create returns mutable TVertex from PBRep;
    	---Level: Internal 

    
    Tolerance(me) returns Real
    is static;
    	---Level: Internal 
    
    Tolerance(me : mutable; T : Real)
    is static;
    	---Level: Internal 

    Pnt(me) returns Pnt from gp
    is static;
    	---Level: Internal 
	
    Pnt(me : mutable; P : Pnt from gp)
    is static;
    	---Level: Internal 

    Points(me) returns PointRepresentation from PBRep
    is static;
    	---Level: Internal 

    Points(me : mutable; P : PointRepresentation from PBRep)
    is static;
    	---Level: Internal 

fields

    myTolerance : Real;
    myPnt       : Pnt from gp;
    myPoints    : PointRepresentation from PBRep;

end TVertex;
