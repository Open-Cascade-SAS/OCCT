-- Created on: 1999-03-24
-- Created by: data exchange team
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class AssemblyLink from STEPSelections inherits TShared from MMgt

	---Purpose: 

uses
    
    NextAssemblyUsageOccurrence from StepRepr,
    ContextDependentShapeRepresentation from StepShape,
    AssemblyComponent from STEPSelections

is

    Create returns mutable AssemblyLink from STEPSelections;
    
    Create(nauo: NextAssemblyUsageOccurrence from StepRepr;
    	   item: Transient from Standard;
	   part: AssemblyComponent from STEPSelections)
    returns mutable AssemblyLink from STEPSelections;
    
    --Methods for setting and obtaining fields
    
    GetNAUO(me) returns NextAssemblyUsageOccurrence from StepRepr;
    	---Purpose:
	---C++: inline
	
    GetItem(me) returns Transient from Standard;
    	---Purpose:
	---C++: inline
	
    GetComponent(me) returns AssemblyComponent from STEPSelections;
    	---Purpose:
	---C++: inline
    
    SetNAUO(me: mutable; nauo: NextAssemblyUsageOccurrence from StepRepr);
    	---Purpose:
	---C++: inline
	
    SetItem(me: mutable; item: Transient from Standard);
    	---Purpose:
	---C++: inline
    
    SetComponent(me: mutable; part: AssemblyComponent from STEPSelections);
	---Purpose:
	---C++: inline

fields

    myNAUO     : NextAssemblyUsageOccurrence from StepRepr;
    myItem     : Transient from Standard;
    myComponent: AssemblyComponent from STEPSelections;

end AssemblyLink;
