-- Created on: 1999-11-26
-- Created by: Andrey BETENEV
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0

class CurveBoundedSurface from StepGeom
inherits BoundedSurface from StepGeom

    ---Purpose: Representation of STEP entity CurveBoundedSurface

uses
    HAsciiString from TCollection,
    Surface from StepGeom,
    HArray1OfSurfaceBoundary from StepGeom

is
    Create returns CurveBoundedSurface from StepGeom;
	---Purpose: Empty constructor

    Init (me: mutable; aRepresentationItem_Name: HAsciiString from TCollection;
                       aBasisSurface: Surface from StepGeom;
                       aBoundaries: HArray1OfSurfaceBoundary from StepGeom;
                       aImplicitOuter: Boolean);
	---Purpose: Initialize all fields (own and inherited)

    BasisSurface (me) returns Surface from StepGeom;
	---Purpose: Returns field BasisSurface
    SetBasisSurface (me: mutable; BasisSurface: Surface from StepGeom);
	---Purpose: Set field BasisSurface

    Boundaries (me) returns HArray1OfSurfaceBoundary from StepGeom;
	---Purpose: Returns field Boundaries
    SetBoundaries (me: mutable; Boundaries: HArray1OfSurfaceBoundary from StepGeom);
	---Purpose: Set field Boundaries

    ImplicitOuter (me) returns Boolean;
	---Purpose: Returns field ImplicitOuter
    SetImplicitOuter (me: mutable; ImplicitOuter: Boolean);
	---Purpose: Set field ImplicitOuter

fields
    theBasisSurface: Surface from StepGeom;
    theBoundaries: HArray1OfSurfaceBoundary from StepGeom;
    theImplicitOuter: Boolean;

end CurveBoundedSurface;
