-- File:        Template.cdl
-- Created:     Mon Dec  4 12:02:32 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWTemplate from RWStepVisual

	---Purpose : Read & Write Module for Template

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     Template from StepVisual,
     EntityIterator from Interface

is

	Create returns RWTemplate;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable Template from StepVisual);

	WriteStep (me; SW : in out StepWriter; ent : Template from StepVisual);

	Share(me; ent : Template from StepVisual; iter : in out EntityIterator);

end RWTemplate;
