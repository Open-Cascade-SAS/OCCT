-- File:	QARoutelous_PresentableObject.cdl
-- Created:	Tue Apr  9 18:33:46 2002
-- Author:	QA Admin
--		<qa@umnox.nnov.matra-dtv.fr>
---Copyright:	 Matra Datavision 2002

class PresentableObject from QARoutelous inherits InteractiveObject from AIS
uses
    Selection from SelectMgr,
    PresentationManager3d from PrsMgr,
    Presentation from Prs3d,
    TypeOfPresentation3d from PrsMgr
is
    
    Create(aTypeOfPresentation3d: TypeOfPresentation3d from PrsMgr = PrsMgr_TOP_AllView) returns mutable PresentableObject from QARoutelous;
    
    ComputeSelection(me:mutable; aSelection :mutable Selection from SelectMgr;
                                 aMode      : Integer) is redefined virtual protected;

    Compute(me:mutable;
    	    aPresentationManager: PresentationManager3d from PrsMgr;
            aPresentation: mutable Presentation from Prs3d;
            aMode: Integer from Standard = 0)
    is redefined virtual protected;
	    
end PresentableObject;
    
