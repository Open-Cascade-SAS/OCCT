-- Created on: 1999-03-10
-- Created by: data exchange team
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DocumentReferenceItem from StepAP214 
inherits SelectType from StepData 


uses
    	Approval from StepBasic,
    	DescriptiveRepresentationItem from StepRepr,
    	MaterialDesignation from StepRepr,
	ProductDefinition from StepBasic,
	ProductDefinitionRelationship from StepBasic,
	PropertyDefinition from StepRepr,
    	Representation from StepRepr,
    	ShapeAspect from StepRepr,
	ShapeAspectRelationship from StepRepr


is
    
    	Create returns DocumentReferenceItem;
	---Purpose : Returns a DocumentReferenceItem SelectType

    	CaseNum (me; ent : Transient) returns Integer ;
	---Purpose: Recognizes a DocumentReferenceItem Kind Entity that is :
    	    	
    	--        1 -> Approval  
	--        2 -> DescriptiveRepresentationItem
    	--        3 -> MaterialDesignation
	--        4 -> ProductDefinition
	--        5 -> ProductDefinitionRelationship
	--        6 -> PropertyDefinition
    	--    	  7 -> 	Representation
    	--    	  8 -> 	ShapeAspect
	--	  9 ->	ShapeAspectRelationship
	--        0 else
	 
    	Approval (me) returns any Approval from StepBasic;
       	---Purpose : returns Value as a Approval (Null if another type)
	
    	DescriptiveRepresentationItem (me) returns any DescriptiveRepresentationItem from StepRepr;
	---Purpose : returns Value as a  (Null if another type)
	
    	MaterialDesignation (me) returns any MaterialDesignation from StepRepr;
	---Purpose : returns Value as a MaterialDesignation (Null if another type)
	
    	ProductDefinition (me) returns any ProductDefinition from StepBasic;
	---Purpose : returns Value as a ProductDefinition (Null if another type)

    	ProductDefinitionRelationship (me) returns any ProductDefinitionRelationship from StepBasic; 
	---Purpose : returns Value as aProductDefinitionRelationship (Null if another type)

    	PropertyDefinition (me) returns any PropertyDefinition from StepRepr;
	---Purpose : returns Value as a PropertyDefinition (Null if another type)
	
    	Representation(me) returns any Representation from StepRepr;
	---Purpose : returns Value as a Representation (Null if another type)
	
	ShapeAspect(me) returns any ShapeAspect  from StepRepr;
	---Purpose : returns Value as a ShapeAspect (Null if another type)
	
	ShapeAspectRelationship(me) returns any ShapeAspectRelationship from StepRepr;
	---Purpose : returns Value as a ShapeAspectRelationship (Null if another type) 


end DocumentReferenceItem;
