-- Created on: 2007-08-22
-- Created by: Sergey ZARITCHNY
-- Copyright (c) 2007-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class AsciiString from PDataStd inherits Attribute from PDF

	---Purpose: Persistance attribute of  TDataStd_AsciiString

uses  HAsciiString from PCollection

is
    Create returns mutable  AsciiString from  PDataStd;
    
    
    Create (V : HAsciiString from PCollection) 
    returns mutable  AsciiString from PDataStd;
    
    
    Get (me) returns HAsciiString from PCollection;
    
    
    Set (me : mutable; V : HAsciiString from PCollection);
    
fields

    myValue : HAsciiString from PCollection;


end AsciiString;
