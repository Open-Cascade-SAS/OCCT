-- Created on: 1997-08-04
-- Created by: VAUTHIER Jean-Claude
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class TagSource from TDF inherits Attribute from TDF

	---Purpose: This attribute manage   a tag provider   to create
	--          child labels of a given one.

uses GUID            from Standard,
     Attribute       from TDF,
     Label           from TDF,
     RelocationTable from TDF
     

is

    ---Purpose: class methods
    --          =============

    
    GetID (myclass)   
    	---C++: return const &  
    returns GUID from Standard;

    Set (myclass; label : Label from TDF)   
    ---Purpose: Find, or create, a  TagSource attribute. the TagSource
    --          attribute is returned.
    returns TagSource from TDF;
    
    NewChild (myclass; L : Label from TDF)
    ---Purpose: Find (or create) a  tagSource attribute located at <L>
    --          and make a new child label.
    returns Label from TDF;
    
    ---Purpose: TagSource methods
    --          =================

    Create
    returns mutable TagSource from TDF;
    
    NewTag (me : mutable)
    returns Integer from Standard;

    NewChild (me : mutable)
    returns Label from TDF;

    Get (me) returns Integer from Standard;

    Set (me : mutable; T : Integer from Standard);
    
    ---Purpose: TDF_Attribute methods
    --          =====================

    ID (me)
    	---C++: return const & 
    returns GUID from Standard;

    Restore (me: mutable; with : Attribute from TDF);


    NewEmpty (me)
    returns mutable Attribute from TDF;


    Paste (me; Into : mutable Attribute from TDF;
	       RT   : mutable RelocationTable from TDF);    

fields
    
    myTag : Integer from Standard;
    
end TagSource;

