-- Created on: 1996-03-05
-- Created by: Joelle CHAUVET
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class MakeApprox from GeomPlate
---Purpose:
-- Allows you to convert a GeomPlate surface into a BSpline.
uses

    Surface        from GeomPlate,
    BSplineSurface from Geom, 
    Shape          from GeomAbs,
    Criterion      from AdvApp2Var


is
    Create(SurfPlate: Surface from GeomPlate;
    	   PlateCrit: Criterion from AdvApp2Var;
    	   Tol3d: Real;
    	   Nbmax: Integer; 
    	   dgmax: Integer; 
     	   Continuity:  Shape  from  GeomAbs  =  GeomAbs_C1;
	   EnlargeCoeff : Real from Standard = 1.1)
    returns MakeApprox;
    ---Purpose:  Converts SurfPlate into a Geom_BSplineSurface with
    --  n Bezier pieces (n<=Nbmax) of degree <= dgmax 
    --  and an approximation error < Tol3d if possible
    --  the criterion CritPlate is satisfied if possible
    
    Create(SurfPlate: Surface from GeomPlate;
    	   Tol3d: Real;
    	   Nbmax: Integer; 
    	   dgmax: Integer;
    	   dmax : Real;
    	   CritOrder: Integer = 0; 
           Continuity:  Shape  from  GeomAbs  =  GeomAbs_C1;
	   EnlargeCoeff : Real from Standard = 1.1)
    returns MakeApprox;
    ---Purpose:  Converts SurfPlate into a Geom_BSplineSurface with
    --  n Bezier pieces (n<=Nbmax) of degree <= dgmax 
    --  and an approximation error < Tol3d if possible
    --  if CritOrder = -1 , no criterion is used
    --  if CritOrder = 0 , a PlateG0Criterion is used with max value > 10*dmax
    --  if CritOrder = 1 , a PlateG1Criterion is used with max value > 10*dmax
    --  WARNING : for CritOrder = 0 or 1, only the constraints points of SurfPlate
    --            are used to evaluate the value of the criterion
    
    Surface(me) returns BSplineSurface from Geom;
    ---Purpose: Returns the BSpline surface extracted from the
    --          GeomPlate_MakeApprox object.   
    
    ApproxError(me) returns Real;
    ---Purpose: Returns the error in computation of the approximation
    --          surface. This is the distance between the entire target
    --          BSpline surface and the entire original surface
    --          generated by BuildPlateSurface and converted by GeomPlate_Surface.    
    CriterionError(me) returns Real;
    ---Purpose: Returns the criterion error in computation of the
    --          approximation surface. This is estimated relative to the
    --          curve and point constraints only.
fields

    myPlate : Surface from GeomPlate;
    mySurface : BSplineSurface from Geom;
    myAppError,myCritError : Real;

end;
