-- Created on: 1995-04-24
-- Created by: Modelistation
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class ChamfSpine from ChFiDS inherits Spine from ChFiDS 

	---Purpose:  Provides  data specific to chamfers 
	--         distances on  each  of faces.
uses
  ChamfMethod from ChFiDS           
 
is
    Create  returns  mutable ChamfSpine from ChFiDS;
    Create (Tol : Real from Standard) returns  mutable ChamfSpine from ChFiDS;
    
    SetDist (me : mutable; Dis : Real from Standard) is static;

    GetDist (me; Dis : in out Real from Standard) is static;    
    
    SetDists (me : mutable; Dis1, Dis2 : Real from Standard) is static;

    Dists (me; Dis1, Dis2 : in out Real from Standard) is static;

    GetDistAngle (me; 
                  Dis, Angle : in out Real from Standard;
                  DisOnF1    : in out Boolean from Standard) is static;
    
    SetDistAngle(me : mutable;
               	 Dis, Angle : Real from Standard;
                 DisOnF1    : Boolean from Standard) is static;

              
    IsChamfer(me) returns ChamfMethod from ChFiDS is static;
    	---Purpose: Return the method of chamfers used 


fields
    d1     : Real        from Standard;
    d2     : Real        from Standard;
    dison1 : Boolean     from Standard;
    angle  : Real        from Standard;
    mChamf : ChamfMethod from ChFiDS;
end ChamfSpine;



