-- Created on: 1998-09-03
-- Created by: Julia GERASIMOVA
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



private class FaceAndOrder from BRepFill

	---Purpose: A structure containing Face and Order of constraint

uses
    Face from TopoDS, 
    Shape from GeomAbs
is
    Create returns FaceAndOrder from BRepFill;
    
    Create( aFace   : Face from TopoDS; 
    	    anOrder : Shape from GeomAbs )
    returns FaceAndOrder from BRepFill;

    --Face(me : in out) returns Face from TopoDS;
    -- ---C++: return &
    --Order(me : in out) returns Integer from Standard;
    -- ---C++: return &

fields

    myFace  : Face from TopoDS;
    myOrder : Shape from GeomAbs;

friends
    class Filling from BRepFill

end FaceAndOrder;
