-- Created on: 1992-09-28
-- Created by: Remi GILET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MakeTranslation

from GC

    	---Purpose: This class mplements elementary construction algorithms for a
    	-- translation in 3D space. The result is a
    	-- Geom_Transformation transformation.
    	-- A MakeTranslation object provides a framework for:
    	-- -   defining the construction of the transformation,
    	-- -   implementing the construction algorithm, and
    	-- -   consulting the result.

uses Pnt            from gp,
     Transformation from Geom,
     Vec            from gp,
     Real           from Standard
     
is

Create(Vect : Vec from gp) returns MakeTranslation;
    	---Purpose: Constructs a translation along the vector " Vect "        
Create(Point1 : Pnt from gp;
       Point2 : Pnt from gp) returns MakeTranslation;
    	---Purpose: Constructs a translation along the vector (Point1,Point2)
    	--  defined from the point Point1 to the point Point2.
    
Value(me) returns Transformation from Geom
    is static;
    	---Purpose:  Returns the constructed transformation.
    	---C++: return const&

Operator(me) returns Transformation from Geom
    is static;
    	---C++: return const&
    	---C++: alias "Standard_EXPORT operator Handle_Geom_Transformation() const;"

fields

    TheTranslation : Transformation from Geom;

end MakeTranslation;

