-- Created on: 1992-09-28
-- Created by: Remi GILET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class MakePlane from GC inherits Root from GC

    ---Purpose : This class implements the following algorithms used 
    --           to create a Plane from gp.
    --           * Create a Plane parallel to another and passing 
    --             through a point.
    --           * Create a Plane passing through 3 points.
    --           * Create a Plane by its normal
    --           A MakePlane object provides a framework for:
    --           -   defining the construction of the plane,
    --           -   implementing the construction algorithm, and
    --           -   consulting the results. In particular, the Value
    --           function returns the constructed plane.
        
uses Pnt       from gp,
     Pln       from gp,
     Ax2       from gp,
     Dir       from gp,
     Plane     from Geom,
     Ax1       from gp,
     Real      from Standard

raises NotDone from StdFail

is

Create (A2 : Ax2)    returns MakePlane;
    --- Purpose :
    --  Creates a plane located in 3D space with an axis placement
    --  two axis.  The "ZDirection" of "A2" is the direction normal
    --  to the plane.  The "Location" point of "A2" is the origin of
    --  the plane. The "XDirection" and "YDirection" of "A2" define
    --  the directions of the U isoparametric and V isoparametric
    --  curves.

Create (Pl : Pln from gp) returns MakePlane;
    --- Purpose :
    --  Creates a plane from a non persistent plane from package gp.

Create (P : Pnt from gp; 
    	V : Dir from gp) returns MakePlane;
    --- Purpose :
    --  P is the "Location" point or origin of the plane.
    --  V is the direction normal to the plane.

Create (A, B, C ,D : Real from Standard) returns MakePlane;
    --- Purpose :
    --  Creates a plane from its cartesian equation :
    --  Ax + By + Cz + D = 0.0
    --  Status is "BadEquation" if Sqrt (A*A + B*B + C*C) 
    --  <= Resolution from gp

Create(Pln    :     Pln from gp;
       Point  :     Pnt from gp) returns MakePlane;
    ---Purpose : Make a Plane from Geom <ThePlane> parallel to another 
    --           Pln <Pln> and passing through a Pnt <Point>.

Create(Pln  : Pln  from gp      ;
       Dist : Real from Standard) returns MakePlane;
    ---Purpose : Make a Plane from Geom <ThePlane> parallel to another 
    --           Pln <Pln> at the distance <Dist> which can be greater 
    --           or lower than zero.
    --           In the first case the result is at the distance 
    --           <Dist> to the plane <Pln> in the direction of the 
    --           normal to <Pln>.
    --           Otherwize it is in the oposite direction.

Create(P1     :     Pnt from gp;
       P2     :     Pnt from gp;
       P3     :     Pnt from gp) returns MakePlane;
    ---Purpose : Make a Plane from Geom <ThePlane> passing through 3
    --           Pnt <P1>,<P2>,<P3>.
    --           It returns false if <P1> <P2> <P3> are confused.

Create(Axis : Ax1 from gp) returns MakePlane;
    ---Purpose: Make a Plane  passing through the location of <Axis>and 
    --          normal to the Direction of <Axis>.

Value(me) returns Plane from Geom
    raises NotDone
    is static;
    ---Purpose: Returns the constructed plane.
    -- Exceptions StdFail_NotDone if no plane is constructed.
    ---C++: return const&

Operator(me) returns Plane from Geom
    is static;
    ---C++: return const&
    ---C++: alias "Standard_EXPORT operator Handle_Geom_Plane() const;"

fields

    ThePlane : Plane from Geom;
    --The solution from Geom.
    
end MakePlane;

