-- Created on: 2004-09-03
-- Created by: Oleg FEDYAEV
-- Copyright (c) 2004-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class CheckResult from BOPAlgo
    ---Purpose: contains information about faulty shapes and faulty types
    ---         can't be processed by Boolean Operations

uses

    Shape       from TopoDS, 
    CheckStatus from BOPAlgo,
    ListOfShape from BOPCol
    
is

    Create
    returns CheckResult;
    ---Purpose: empty constructor
    
    SetShape1(me: in out; TheShape : Shape from TopoDS);
    ---Purpose: sets ancestor shape (object) for faulty sub-shapes
    
    AddFaultyShape1(me: in out; TheShape: Shape from TopoDS);
    ---Purpose: adds faulty sub-shapes from object to a list
    
    SetShape2(me: in out; TheShape: Shape from TopoDS);
    ---Purpose: sets ancestor shape (tool) for faulty sub-shapes
    
    AddFaultyShape2(me: in out; TheShape: Shape from TopoDS);
    ---Purpose: adds faulty sub-shapes from tool to a list
    
    GetShape1(me)
    returns Shape from TopoDS;
    ---C++: return const&
    ---Purpose: returns ancestor shape (object) for faulties

    GetShape2(me)
    returns Shape from TopoDS;
    ---C++: return const&
    ---Purpose: returns ancestor shape (tool) for faulties

    GetFaultyShapes1(me)
    returns ListOfShape from BOPCol;
    ---C++: return const&
    ---Purpose: returns list of faulty shapes for object

    GetFaultyShapes2(me)
    returns ListOfShape from BOPCol;
    ---C++: return const&
    ---Purpose: returns list of faulty shapes for tool

    SetCheckStatus(me: in out; TheStatus: CheckStatus from BOPAlgo);
    ---Purpose: set status of faulty
    
    GetCheckStatus(me)
    returns CheckStatus from BOPAlgo;
    ---Purpose: gets status of faulty
  
fields

    myShape1 : Shape from TopoDS;
    myShape2 : Shape from TopoDS;
    myStatus : CheckStatus from BOPAlgo;
    myFaulty1 : ListOfShape from BOPCol;
    myFaulty2 : ListOfShape from BOPCol;

end CheckResult;
