-- Created on: 1993-01-09
-- Created by: CKY / Contract Toubro-Larsen ( Anand NATRAJAN )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class AssocGroupType from IGESBasic  inherits IGESEntity

        ---Purpose: defines AssocGroupType, Type <406> Form <23>
        --          in package IGESBasic
        --          Used to assign an unambiguous identification to a Group
        --          Associativity.

uses

        HAsciiString from TCollection

is

        Create returns mutable AssocGroupType;

        -- Specific Methods pertaining to the class

        Init (me : mutable; nbDataFields, aType : Integer; 
              aName : HAsciiString );
        ---Purpose : This method is used to set the fields of the class
        --           AssocGroupType
        --       - nbDataFields : number of parameter data fields = 2
        --       - aType        : type of attached associativity
        --       - aName        : identifier of associativity of type AType

        NbData (me) returns Integer;
        ---Purpose : returns the number of parameter data fields, always = 2

        AssocType (me) returns Integer;
        ---Purpose : returns the type of attached associativity

        Name (me) returns HAsciiString from TCollection;
        ---Purpose : returns identifier of instance of specified associativity

fields

--
-- Class    : IGESBasic_AssocGroupType
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class AssocGroupType.
--
-- Reminder : A AssocGroupType instance is defined by :
--            - the number of parameter data fields, always = 2
--            - the type of attached associativity
--            - the identifier of instance of specified associativity

        theNbData : Integer;
        theType   : Integer;
        theName   : HAsciiString from TCollection;

end AssocGroupType;
