-- Created on: 1995-06-13
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class LocalOperation from BRepFeat inherits Builder from BRepFeat

	---Purpose: One of the most significant
	-- aspects of BRepFeat functionality is the use of local operations as
	-- opposed to global ones. In a global operation, you would first
	-- construct a form of the type you wanted in your final feature, and
	-- then remove matter so that it could fit into your initial basis
	-- object. In a local operation, however, you specify the domain
	-- of the feature construction with aspects of the shape on which the
	-- feature is being created. These semantics are expressed in terms
	-- of a member shape of the basis shape from which - or up to which
	-- - matter will be added or removed. As a result, local
	-- operations make calculations simpler and faster than global operations.
	-- In BRepFeat, the semantics of local operations define features
	-- constructed from a contour or a part of the basis shape referred to as the tool.

uses 
    Shape       from TopoDS,
    ListOfShape from TopTools

raises
    NotDone           from StdFail,
    ConstructionError from Standard

is

    Create
	---Purpose: Builds the framework to store the topological shape
	-- which is to be created by the local operation.
	-- Initializes the empty constructor.
      	returns LocalOperation from BRepFeat;
        ---C++: inline	

	 
    Create(S: Shape from TopoDS)
	---C++: inline
	---Purpose: Builds the framework to store the topological shape
	-- which is to be created by the local operation.
	-- Initializes shape S for a local operation.
	-- The exception ConstructionError is raised if <S> is a null shape.
	returns LocalOperation from BRepFeat
	raises ConstructionError from Standard;


    Create(S1,S2: Shape from TopoDS)
	---C++: inline
	---Purpose: Builds the framework to store the topological shape
	-- which is to be created by the local operation.
	-- Initializes S1 and S2 for a local operation.
	-- The exception ConstructionError is raised if <S> is a null shape.
    	returns LocalOperation from BRepFeat
	raises ConstructionError from Standard;

--  Init(me: in out; S: Shape from TopoDS) is inherited from BRepFeat_Builder.

--  Init(me: in out; S,T: Shape from TopoDS) is inherited from BRepFeat_Builder.


    Perform(me: in out; T    : Shape from TopoDS;
                        L    : ListOfShape from TopTools;
                        Fuse : Boolean from Standard)
	---Purpose: Performs the local operation on the formerly given
	--          shape,  with the tool <T>.  <L>  defines  a set of
	--          faces  of  the shape.  The list  may not be empty.
	--          The boolean <Fuse> gives the type of operation. If
	--          set to  Standard_True, the operation  is a fusion.
	--          If  set  to Standard_False,   the operation   is a
	--          cutting one.
	--          
	--          The Perform process stops just before constructing
	--          any result in order to authorize  the selection of
	--          parts of the tool.  After a call to Perform, it is
	--          possible   to call     BuilPartsOfTool,       then
	--          RemovePart/ActivatePart to select valid parts, and
	--          it  is necessary to  call PerformResult to get any
	--          result. 
	---C++: inline

	raises ConstructionError from Standard
	--- The exception is raised if <T> is null or same as the shape.
    	is static;



    Perform(me: in out; LShape : ListOfShape from TopTools;
                        LTool  : ListOfShape from TopTools;
                        Fuse   : Boolean from Standard)

	---Purpose: Performs the local operation on the formerly given
	--          shape and tool.  <LShape>  defines a set  of faces
	--          of the shape, <LTool> a set of  faces of the tool.
	--          The boolean  <Fuse> gives the  type of  operation.
	--          If  set  to   Standard_True,  the operation  is  a
	--          fusion.   If  set to Standard_False, the operation
	--          is a cutting one.  If <LShape> (resp.  <LTool>) is
	--          empty, the whole shape (resp.  tool) is used. 
	--          
	--          The Perform process stops just before constructing
	--          any result in  order to authorize the selection of
	--          parts of the tool.  After a call to Perform, it is
	--          possible     to   call     BuilPartsOfTool,   then
	--          RemovePart/ActivatePart to select valid parts, and
	--          it is necessary  to call PerformResult to  get any
	--          result.  
	---C++: inline

	raises ConstructionError from Standard
	--- The exception is raised if <T> is a null shape.
    	is static;



    BuildPartsOfTool(me: in out)
	---Purpose: Constructs the primitive which serves as the tool for the
    	-- feature construction. Gives faces concerned by the
    	-- construction and builds by performing one of the
    	-- Boolean operations on the two intersecting shapes.
    	--    Raises NotDone from StdFail if no call to Perform has been done.
    		---C++: inline
    	    	raises NotDone from StdFail
	    	is static;
    

    PartsOfTool(me)
	---Purpose: Returns  the list of  the  parts of tool.  Each of
	--          these parts is a TopoDS_Shell.
    	-- Raises NotDone  if no  call to BuildPartsOfTool has been done. 
    returns ListOfShape from TopTools
	---C++: return const&
	---C++: inline
    	raises NotDone from StdFail
	
	is static;


    RemovePart(me: in out; S: Shape from TopoDS)
	---Purpose: Removes <S> from the list of valid parts of tool.
	-- Raises NotDone  if no  call to BuildPartsOfTool has
	-- been done. 
    		---C++: inline
    	    	raises NotDone from StdFail
	    	is static;


    ActivatePart(me: in out; S: Shape from TopoDS)
	---Purpose: By default, all tool parts are valid for the local operation.
    	--        This method removes <S>  from  the list  of  invalid parts  of
	--          tool. By default, all parts  of tool are valid for
	--          the local operation.
	---C++: inline
    	raises NotDone from StdFail
	-- The exception is raised if no  call to BuildPartsOfTool has
	-- been done. 
    	is static;
	
--- Redefinition of BRepBuilderAPI_MakeShape methods
--  
--  

    Build(me: in out)
	---Purpose: Builds the    resulting shape  (redefined     from
	--          MakeShape). Invalidates the  given parts  of tools
	--          if  any,   and performs the  result   of the local
	--          operation.

    	is redefined;

end LocalOperation;
