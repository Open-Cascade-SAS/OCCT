-- File:        PlanarBox.cdl
-- Created:     Mon Dec  4 12:02:28 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWPlanarBox from RWStepVisual

	---Purpose : Read & Write Module for PlanarBox

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     PlanarBox from StepVisual,
     EntityIterator from Interface

is

	Create returns RWPlanarBox;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable PlanarBox from StepVisual);

	WriteStep (me; SW : in out StepWriter; ent : PlanarBox from StepVisual);

	Share(me; ent : PlanarBox from StepVisual; iter : in out EntityIterator);

end RWPlanarBox;
