-- File:        CameraImage.cdl
-- Created:     Mon Dec  4 12:02:24 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWCameraImage from RWStepVisual

	---Purpose : Read & Write Module for CameraImage

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     CameraImage from StepVisual,
     EntityIterator from Interface

is

	Create returns RWCameraImage;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable CameraImage from StepVisual);

	WriteStep (me; SW : in out StepWriter; ent : CameraImage from StepVisual);

	Share(me; ent : CameraImage from StepVisual; iter : in out EntityIterator);

end RWCameraImage;
