-- Created on: 1993-07-05
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Update:      Frederic MAUPAS



deferred class CurveRepresentation from PBRep inherits Persistent

	---Purpose: Root class for the curve representations.

uses
    Location from PTopLoc


is

    Initialize(L : Location from PTopLoc);
    	---Level: Internal 

    Location(me) returns Location from PTopLoc
    is static;
    	---Level: Internal 
    
    Next(me) returns CurveRepresentation from PBRep
    is static;
    	---Level: Internal 
		
    Next(me : mutable; N :  CurveRepresentation from PBRep)
    is static;
    	---Level: Internal 

    ------------------------------------------------------
    -- What kind of representation : used to speed Mapping
    ------------------------------------------------------

    IsCurve3D(me)               returns Boolean
	 ---Purpose: A 3D curve representation.
    is virtual;

    IsCurveOnSurface(me)        returns Boolean
	---Purpose: A curve in the parametric space of a surface.
    is virtual;

    IsRegularity(me)            returns Boolean
	---Purpose: A continuity between two surfaces.
    is virtual;
    
    IsCurveOnClosedSurface(me)  returns Boolean
	---Purpose: A curve with two parametric   curves  on the  same
	--          surface. 
    is virtual;

    IsGCurve(me) returns Boolean from Standard
    	---Purpose:
    is virtual;
    
    IsPolygon3D(me) returns Boolean
	---Purpose: 
    is virtual;
    
    IsPolygonOnTriangulation(me) returns Boolean
	---Purpose: 
    is virtual;

    IsPolygonOnClosedTriangulation(me) returns Boolean
	---Purpose: 
    is virtual;

    IsPolygonOnSurface(me) returns Boolean
	---Purpose: 
    is virtual;

    IsPolygonOnClosedSurface(me) returns Boolean
	---Purpose: 
    is virtual;
    
    
fields
    
    myLocation : Location from PTopLoc;
    myNext     : CurveRepresentation from PBRep;

end CurveRepresentation;
