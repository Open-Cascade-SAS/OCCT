-- Created on: 2000-09-29
-- Created by: Pavel TELKOV
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class GraphNode from PXCAFDoc inherits Attribute from PDF

	---Purpose: 

uses
    Attribute         from PDF,
    GUID              from Standard,
    GraphNodeSequence from PXCAFDoc

is
    Create returns mutable GraphNode from PXCAFDoc;
    
    SetFather (me : mutable;F : GraphNode from PXCAFDoc)
    returns Integer from Standard;

    SetChild (me : mutable;Ch : GraphNode from PXCAFDoc)
    returns Integer from Standard;
    
    GetFather (me ; Findex : Integer from Standard)
    returns GraphNode from PXCAFDoc;
	
    GetChild (me ; Chindex : Integer from Standard)
    returns GraphNode from PXCAFDoc;
    
    FatherIndex (me ; F : GraphNode from PXCAFDoc)
    returns Integer from Standard;
    
    ChildIndex (me ; Ch : GraphNode from PXCAFDoc)
    returns Integer from Standard;

    NbFathers (me) returns Integer from Standard;

    NbChildren (me) returns Integer from Standard;

    SetGraphID(me : mutable; GUID : GUID from Standard);

    GetGraphID(me) returns GUID from Standard;

fields

	myFathers  : GraphNodeSequence from PXCAFDoc;
	myChildren : GraphNodeSequence from PXCAFDoc;
    	myGraphID  : GUID              from Standard;
	
end GraphNode;
