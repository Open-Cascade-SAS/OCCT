-- Created on: 1993-03-23
-- Created by: BBL
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


deferred class ColorMap from Aspect inherits TShared from MMgt

	---Version: 0.0

	---Purpose: This class defines a ColorMap object.
	---Keywords:
	---Warning:
	---References:
uses
	Color			from Quantity,
	TypeOfColorMap 		from Aspect,
	ColorMapEntry 		from Aspect,
	SequenceOfColorMapEntry from Aspect

raises
	BadAccess 	from Aspect

is

	Initialize( type : TypeOfColorMap from Aspect );

	Type( me )
	returns TypeOfColorMap from Aspect is static;
	---Level: Public

	Size( me ) returns Integer from Standard is static;
	---Level: Public
	---Purpose: Returns the Allocated colormap Size

	Index( me ; aColormapIndex : Integer ) returns Integer from Standard
	---Level: Public
	---Purpose: Returns the ColorMapEntry.Index of the ColorMap  
	--	    at rank <aColormapIndex> .
	raises BadAccess from Aspect is static;
	---Trigger: Raises BadAccess if the index less than 1 or
	--	    greater than Size.

	Dump( me ) ;
	---Level: Internal

	Entry ( me ; AColorMapIndex : Integer from Standard )
	returns ColorMapEntry from Aspect
	---Level: Public
    	---Purpose: Return the value of the <Index>th element of
	--	    the ColorMap
	raises BadAccess from Aspect is static;
	---Trigger: Raises BadAccess if the index less than 1 or
	--	    greater than Size.
    	---C++: return const &

	FindColorMapIndex ( me ;
		AColorMapEntryIndex : Integer from Standard )
		returns Integer from Standard
	---Level: Public
	---Purpose: Returns the index in the ColorMap of the 
	--	    ColorMapEntry.Index() equal to <AnEntryIndex>.
		raises BadAccess from Aspect is deferred ;
	---Trigger: Raises BadAccess if the index is not defined in the
	--	    ColorMap.

	FindEntry ( me ; AColorMapEntryIndex : Integer from Standard )
		returns ColorMapEntry from Aspect
	---Level: Public
	---Purpose: Returns the ColorMapEntry with ColorMapEntry.Index()
	--	    equal to <AnEntryIndex>.
		raises BadAccess from Aspect is deferred ;
	---Trigger: Raises BadAccess if the index is not defined in the
	--	    ColorMap.
    	---C++: return const &

	NearestColorMapIndex( me ; aColor : Color from Quantity )
		returns Integer from Standard is deferred ;
	---Level: Public
	---Purpose: Returns the index in the ColorMap of the
	--	    nearest matching ColorMapEntry 

	NearestEntry( me ; aColor : Color from Quantity )
		returns ColorMapEntry from Aspect is deferred ;
	---Level: Public
	---Purpose: Returns the nearest ColorMapEntry that match aColor .
    	---C++: return const &

        AddEntry (me : mutable; aColor : Color from Quantity)
             	returns Integer from Standard is deferred;
        ---Level: Public
        ---Purpose: Search an identical color entry in the color map <me>
        -- and returns the ColorMapEntry Index if exist.
        -- Or add a new entry and returns the computed ColorMapEntry index used.

fields

	mytype		: TypeOfColorMap	  from Aspect;
	mydata		: SequenceOfColorMapEntry from Aspect is protected;

end ColorMap ;
