-- File:	math_ComputeKronrodPointsAndWeights.cdl
-- Created:	Wed Dec 21 18:07:18 2005
-- Author:	Julia GERASIMOVA
--		<jgv@clubox>
---Copyright:	 Matra Datavision 2005

class ComputeKronrodPointsAndWeights from math 

uses 
 
    Vector from math, 
    HArray1OfReal from TColStd

is 
    Create(Number : Integer from Standard) 
    returns ComputeKronrodPointsAndWeights; 

    IsDone(me) 
    returns Boolean from Standard;

    Points(me) 
    returns Vector from math;

    Weights(me)
    returns Vector from math;

fields 
 
    myPoints  : HArray1OfReal from TColStd;
    myWeights : HArray1OfReal from TColStd; 
    myIsDone  : Boolean from Standard;
     
end ComputeKronrodPointsAndWeights;
