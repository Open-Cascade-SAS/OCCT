-- Created on: 1995-01-23
-- Created by: Mister rmi
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class SensitiveEntity from SelectBasics inherits TShared from MMgt

  ---Purpose: root class; the inheriting classes will be able to give
  --          sensitive Areas for the dynamic selection algorithms

uses 
    EntityOwner,
    BndBox3d from Select3D,
    PickResult,
    SelectingVolumeManager

is


    Initialize (theOwnerId       : EntityOwner;
                theSensFactor    : Real from Standard = 2.0);

    Set (me : mutable;
         theOwnerId : EntityOwner)
      is virtual;
    ---Level: Public
    ---Purpose: Sets owner of the entity


    OwnerId (me)
      returns any EntityOwner
      is static;
    ---Level: Public 
    ---C++: return const&
    ---Purpose: Returns pointer to owner of the entity


    Matches (me           : mutable;
            theMgr        : out SelectingVolumeManager from SelectBasics;
            thePickResult : out PickResult from SelectBasics)
    returns Boolean is deferred;
    ---Level: Public
    ---Purpose: Checks whether the sensitive entity is overlapped by
    --          current selecting volume

    SetSensitivityFactor (me : mutable;
                          theSensFactor :Real from Standard);
    ---C++: inline
    ---Purpose: Allows to manage the sensitivity of the entity

    SensitivityFactor (me)
      returns Real from Standard;
    ---C++: inline
    ---Purpose: allows a better sensitivity for
    --          a specific entity in selection algorithms
    --          useful for small sized entities.

    NbSubElements (me : mutable) returns Integer from Standard
    is deferred;
    ---Purpose: Returns the number of sub-entities or elements in
    --          sensitive entity. Is used to determine if entity is
    --          complex and needs to pre-build BVH at the creation of
    --          sensitive entity step or is light-weighted so the tree
    --          can be build on demand with unnoticeable delay

    BoundingBox (me : mutable) returns BndBox3d from Select3D is deferred;
    ---Purpose: Returns bounding box of sensitive entity

    BVH (me : mutable) is deferred;
    ---Purpose: Builds BVH tree for sensitive if it is needed

    Clear (me : mutable) is deferred;
    ---Purpose: Clears up all the resources and memory allocated


fields
    
    myOwnerId       : EntityOwner from SelectBasics is protected;
    mySFactor       : Real from Standard;
end SensitiveEntity;
