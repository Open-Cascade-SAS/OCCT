-- Created on: 1997-11-17
-- Created by: Jean-Louis Frenkel
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


deferred class MetaDataDriver from CDF inherits Transient from Standard


uses
    Document from CDM, MetaData from CDM,
    ExtendedString from TCollection,
    ReferenceIterator from PCDM
    
raises 
    NotImplemented from Standard
is

    Initialize;

    ---Category: virtual methods

    HasVersionCapability(me: mutable)
    ---Purpose: returns true if the MetaDataDriver can manage different
    --          versions of a Data.
    --          By default, returns Standard_False.
    returns Boolean from Standard
    is virtual;

    CreateDependsOn(me: mutable; aFirstData: MetaData from CDM;
                                aSecondData: MetaData from CDM)
    ---Purpose: Creates a "Depends On"  relation between two Datas.
    --          By default does nothing
    is virtual;
    
    CreateReference(me: mutable; aFrom, aTo: MetaData from CDM; aReferenceIdentifier: Integer from Standard; aToDocumentVersion: Integer from Standard)
    is virtual;
    
    HasVersion(me: mutable; aFolder, aName: ExtendedString from TCollection)
    returns Boolean from Standard
    ---Purpose: by default return Standard_True.
    is virtual;
    
    BuildFileName(me: mutable; aDocument: Document from CDM)
    returns ExtendedString from TCollection
    is deferred;

    SetName(me: mutable; aDocument: Document from CDM; aName: ExtendedString from TCollection)
    returns ExtendedString from TCollection
    is virtual;
    ---Purpose: this methods  is usefull if the name  of an  object --
    --           depends on  the metadatadriver. For  example a Driver
    --           -- based  on the operating  system can choose to  add
    --           the extension of file to create to the object.
    
---Category: Deferred methods

    ---Overview: inquiring can be made either using a folder, a name and eventually
    --           a version 
    --           or a path which is the concatenation of a folder, a name  and eventually
    --           a version.
    Find(me: mutable; aFolder, aName, aVersion: ExtendedString from TCollection)
    returns Boolean from Standard
    ---Purpose: should indicate whether meta-data exist in the DBMS corresponding 
    --          to the Data.
    --          aVersion may be NULL;
    is deferred;
    
    HasReadPermission(me: mutable; aFolder, aName, aVersion: ExtendedString from TCollection)
    returns Boolean from Standard
    is deferred;
    
    MetaData(me: mutable; aFolder, aName, aVersion: ExtendedString from TCollection)
    returns MetaData from CDM
    ---Purpose: should return the MetaData stored in the DBMS with the meta-data
    --          corresponding to the Data. If the MetaDataDriver has version management capabilities
    --          the version has to be set in the returned MetaData.
    --          aVersion may be NULL
    --          MetaData is called by GetMetaData
    --          If the version is  set to NULL, MetaData should return
    --          the last version of the metadata 
    is deferred;
    
    LastVersion(me: mutable; aMetaData: MetaData from CDM)
    returns MetaData from CDM
    is virtual;
    ---Purpose: by default returns aMetaDATA
	    
--    MetaData(me: mutable; aPath: ExtendedString from TCollection)
--    returns MetaData from CDM
    ---Purpose: should return the MetaData stored in the DBMS with the meta-data
    --          corresponding to the path. If the MetaDataDriver has version management capabilities
    --          the version has to be set in the returned MetaData.
    --          MetaData is called by GetMetaData
    --          If the version is not included in the path , MetaData should return
    --          the last version of the metadata 
--    is deferred;
    


    
    CreateMetaData(me: mutable; aDocument: Document from CDM;
    	         aFileName: ExtendedString from TCollection)
    ---Purpose:  should create meta-data corresponding to aData and maintaining a meta-link
    --           between these meta-data and aFileName
    --           CreateMetaData is called by CreateData
    returns  MetaData from CDM
    ---Purpose: If the metadata-driver 
    --          has version capabilities, version must be set in the returned Data.
    is deferred;
    
    FindFolder(me: mutable; aFolder: ExtendedString from TCollection)
    returns Boolean from Standard
    is deferred;

   DefaultFolder(me: mutable) returns ExtendedString from TCollection
   is deferred;
   
   
---Category:  methods about references.

    ReferenceIterator(me: mutable)
    returns ReferenceIterator from PCDM
    is virtual;
    

    Find(me: mutable; aFolder, aName: ExtendedString from TCollection)
    returns Boolean from Standard;
    ---Purpose: calls Find with an empty version

    MetaData(me: mutable; aFolder, aName: ExtendedString from TCollection)
    returns MetaData from CDM;
    ---Purpose: calls MetaData with an empty version
    

end MetaDataDriver from CDF;
