-- Created on: 1999-02-26
-- Created by: Christian CAILLET
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SelectPCurves  from IGESSelect    inherits SelectExplore

    ---Purpose : This Selection returns the pcurves which lie on a face
    --           In two modes : global (i.e. a CompositeCurve is not explored)
    --           or basic (all the basic curves are listed)

uses AsciiString from TCollection, Transient, EntityIterator, Graph

is

    Create (basic : Boolean) returns mutable SelectPCurves;
    ---Purpose : Creates a SelectPCurves
    --           basic True  : lists all the components of pcurves
    --           basic False : lists the uppest level definitions
    --             (i.e. stops at CompositeCurve)

    Explore (me; level : Integer; ent : Transient; G : Graph;
    	     explored : in out EntityIterator)
    	returns Boolean;
    ---Purpose : Explores an entity, to take its contained PCurves
    --           An independant curve is IGNORED : only faces are explored

    ExploreLabel (me) returns AsciiString from TCollection;
    ---Purpose : Returns a text defining the criterium : "Basic PCurves" or
    --           "Global PCurves"

fields

    thebasic : Boolean;

end SelectPCurves;
