-- Created by: Peter KURNEV
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class ShrunkRange from BOPInt 

	---Purpose:  
	---  The class provides the computation of 
	---  a working (shrunk) range [t1, t2] for 
    	---  the 3D-curve of the edge. 
	 
uses
    Box from Bnd, 
    Edge from TopoDS, 
    Vertex from TopoDS, 
    Context  from BOPInt

--raises

is 
    Create 
    	returns ShrunkRange from BOPInt;

    SetData (me:out; 
    	    aE  : Edge from TopoDS;  
    	    aT1 : Real from Standard;              
	    aT2 : Real from Standard;     
	    aV1 : Vertex from TopoDS;              
	    aV2 : Vertex from TopoDS; 
    	    ICtx: Context from BOPInt);   

    SetShrunkRange(me:out; 
    	    aT1 : Real from Standard;   
    	    aT2 : Real from Standard);   

    ShrunkRange(me; 
    	    aT1 :out Real from Standard;   
    	    aT2 :out Real from Standard); 
  
    BndBox  (me) 
    	returns Box from Bnd; 
    ---C++: return const & 
     
    Edge  (me) 
    	returns Edge from TopoDS; 
    ---C++: return const &	 
	     
    Perform(me:out); 
	 
    ErrorStatus(me) 
    	returns Integer from Standard;  
	---Purpose:
	--- Returns code of computing shrunk range
	--- completion
	--- 0 - means successful completion
	--- 1 - nothing has been done
	--- 2 - initial range is out of edge's range
	--- 3 - first boundary of initial range is more than
	---     last boundary
	--- 4 - projection of first vertex failed
	--- 5 - projection of second vertex failed
	--- 6 - shrunk range can not be computed
	---     shrunk range is setted to initial range
	---

fields
    myEdge        : Edge from TopoDS is protected; 
    myV1          : Vertex from TopoDS is protected;
    myV2          : Vertex from TopoDS is protected;  
    myT1          : Real from Standard is protected;     
    myT2          : Real from Standard is protected;     
    myTS1         : Real from Standard is protected;     
    myTS2         : Real from Standard is protected;     
    myBndBox      : Box from Bnd is protected;  
    myCtx         : Context from BOPInt is protected;
    myErrorStatus : Integer from Standard is protected;   
     
end ShrunkRange;
