-- Created on: 1993-10-14
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Common from BRepAlgoAPI inherits BooleanOperation from BRepAlgoAPI

	---Purpose: The class Common provides a
    	-- Boolean common operation on a pair of arguments (Boolean Intersection).
    	--  The class Common provides a framework for:
    	-- -           Defining the construction of a common shape;
    	-- -           Implementing the   building algorithm
    	-- -           Consulting the result.

uses
    Shape from TopoDS, 
    PaveFiller from BOPAlgo

is
    Create (S1,S2 : Shape from TopoDS)  
    	returns Common from BRepAlgoAPI;  
	---Purpose: Constructs a common part for shapes aS1 and aS2 .
 
    Create (S1,S2 : Shape from TopoDS; 
    	    aDSF:PaveFiller from BOPAlgo)  
    	returns Common from BRepAlgoAPI;
end Common;
--- Purpose: Constructs a common part for shapes aS1 and aS2 using aDSFiller
