-- Created on: 1991-07-16
-- Created by: Christophe MARION
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




deferred class Drawable from DrawTrSurf inherits Drawable3D from Draw

	---Purpose: this  class adds   to   the Drawable3D methods  to
	--          display Curves and Curves on Surface.
	--          
	--          The discretisation,  number  of points on a Curve,
	--          is stored in this class.

uses
    Display        from Draw,
    Curve          from Adaptor3d,
    Curve2d        from Adaptor2d,
    IsoCurve       from Adaptor3d,
    IsoType        from GeomAbs

is
    Initialize(discret : Integer; deflection : Real = 0.01; DrawMode : Integer = 0);
	---Purpose: set the number of points on a curve at creation.
	
    DrawCurve2dOn(me;
                C : in out Curve2d from Adaptor2d;
    	        D : in out Display from Draw);
	---Purpose: Draw a polygon of the curve on the Display
	
    DrawCurveOn(me;
                C : in out Curve from Adaptor3d;
    	        D : in out Display from Draw);
	---Purpose: Draw a polygon of the curve on the Display
	
    DrawIsoCurveOn(me;
                C : in out IsoCurve from Adaptor3d;
		T : IsoType from GeomAbs;
		P, F, L : Real;
    	        D : in out Display from Draw);
	---Purpose: Load C  with the specified iso  and Draw a polygon
	--          of the curve on the Display
	
    DrawOn(me; dis : in out Display from Draw)
	---Purpose: this is defined only to tell C++ not to complain
	--          about inheriting a pure virtual method.
    is deferred;

   
    SetDiscretisation (me : mutable; Discret : Integer);
        ---C++: inline
    
    GetDiscretisation (me) returns Integer;
        ---C++: inline
    
    SetDeflection (me : mutable; Deflection : Real);
        ---C++: inline
    
    GetDeflection (me) returns Real;
        ---C++: inline

    SetDrawMode (me : mutable; DrawMode : Integer);
        ---C++: inline
    
    GetDrawMode (me) returns Integer;
        ---C++: inline

        

    
fields
    myDrawMode   : Integer;
       --- Purpose : 0 parametre constant, 1 fleche constante
    myDiscret    : Integer;
    myDeflection : Real;

end Drawable;

