-- Created on: 1993-06-18
-- Created by: Didier PIFFAULT
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ComparatorOfVertexOfDelaun from BRepMesh

  ---Purpose: Sort two point in a given direction.


  uses  Boolean from Standard,
        Vertex from BRepMesh,
        XY from gp


  is      Create (theDir : XY from gp) 
            returns ComparatorOfVertexOfDelaun;


          IsLower (me; Left, Right: Vertex from BRepMesh)
          ---Purpose: returns True if <Left> is lower than <Right>
          returns Boolean from Standard;

          IsGreater (me; Left, Right: Vertex from BRepMesh)
          ---Purpose: returns True if <Left> is greater than <Right>
          returns Boolean from Standard;

          IsEqual(me; Left, Right: Vertex from BRepMesh)
          ---Purpose: returns True when <Right> and <Left> are equal.
          returns Boolean from Standard;


fields  DirectionOfSort : XY from gp;
        Tolerance       : Real from Standard;

end ComparatorOfVertexOfDelaun;
