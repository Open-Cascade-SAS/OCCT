-- Created on: 1995-05-04
-- Created by: Dieter THIEMANN
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MakeHyperbola from GeomToStep inherits Root from GeomToStep

    ---Purpose: This class implements the mapping between the class
    --          Hyperbola from Geom and the class Hyperbola from
    --          StepGeom which describes a Hyperbola from ProSTEP


uses Hyperbola from Geom,
     Hyperbola from Geom2d,
     Hyperbola from StepGeom
     
raises NotDone from StdFail

is

Create ( C : Hyperbola from Geom2d) returns MakeHyperbola;

Create ( C : Hyperbola from Geom) returns MakeHyperbola;


Value (me) returns Hyperbola from StepGeom
    raises NotDone
    is static;
    ---C++: return const&


fields

    theHyperbola : Hyperbola from StepGeom;
    	-- The solution from StepGeom

end MakeHyperbola;
