-- Created on: 1994-08-26
-- Created by: Frederic MAUPAS
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MakeConic2d from StepToGeom

    ---Purpose: This class implements the mapping between classes 
    --          Conic from StepGeom
    --          which describes a Conic from prostep and Conic from Geom2d.
    --          As Conic is an abstract class
    --          this class is an access to the sub-class required.
  
uses Conic from Geom2d,
     Conic from StepGeom
     
is 

    Convert ( myclass; SC : Conic from StepGeom;
                       CC : out Conic from Geom2d )
    returns Boolean from Standard;

end MakeConic2d;
