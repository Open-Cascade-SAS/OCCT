-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PresentationSizeAssignmentSelect from StepVisual inherits SelectType from StepData

	-- <PresentationSizeAssignmentSelect> is an EXPRESS Select Type construct translation.
	-- it gathers : PresentationView, PresentationArea, AreaInSet

uses

	PresentationView,
	PresentationArea,
	AreaInSet
is

	Create returns PresentationSizeAssignmentSelect;
	---Purpose : Returns a PresentationSizeAssignmentSelect SelectType

	CaseNum (me; ent : Transient) returns Integer;
	---Purpose: Recognizes a PresentationSizeAssignmentSelect Kind Entity that is :
	--        1 -> PresentationView
	--        2 -> PresentationArea
	--        3 -> AreaInSet
	--        0 else

	PresentationView (me) returns any PresentationView;
	---Purpose : returns Value as a PresentationView (Null if another type)

	PresentationArea (me) returns any PresentationArea;
	---Purpose : returns Value as a PresentationArea (Null if another type)

	AreaInSet (me) returns any AreaInSet;
	---Purpose : returns Value as a AreaInSet (Null if another type)


end PresentationSizeAssignmentSelect;

