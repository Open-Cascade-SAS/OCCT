-- Created on: 2002-02-01
-- Created by: QA Admin
-- Copyright (c) 2002-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


package QADraw
    uses Draw,
         TCollection
is
    
    class DataMapOfAsciiStringOfAddress instantiates 
		    DataMap from TCollection(AsciiString from TCollection,
					     Address from Standard,
					     AsciiString from TCollection);

    CommonCommands(DI : in out Interpretor from Draw);
    ---Purpose: Define specicial commands for AIS.

    AdditionalCommands(DI : in out Interpretor from Draw);
    
    Factory (DI : out Interpretor from Draw);
    ---Purpose: Loads all QA Draw commands. Used for plugin.

end;
    
