-- Created on: 2006-08-08
-- Created by: Galina KULIKOVA
-- Copyright (c) 2006-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ShapeDivideArea from ShapeUpgrade  inherits ShapeDivide from ShapeUpgrade

	---Purpose: Divides faces from sprcified shape  by max area criterium.

uses

    Shape from TopoDS,
    FaceDivide from ShapeUpgrade

is
     Create returns ShapeDivideArea from ShapeUpgrade;
    	---Purpose:
    
    Create (S: Shape from TopoDS)
    returns ShapeDivideArea from ShapeUpgrade;
    	---Purpose: Initialize by a Shape.
	
    GetSplitFaceTool (me) returns FaceDivide from ShapeUpgrade
    is redefined protected;
    	---Purpose: Returns the tool for splitting faces. 
	

     MaxArea(me: in out) returns Real;
    ---C++: inline
    ---C++: return &
    ---Purpose:Set max area allowed for faces 	

    
fields

    myMaxArea : Real;

end ShapeDivideArea;
