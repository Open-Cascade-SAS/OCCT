-- Created on: 1991-09-05
-- Created by: J.P. TIRAUlt
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

--              C. LEYNADIER 

package Standard

    ---Purpose: 
    --   The package Standard provides the minimum services necessary 
    --   for other toolkits to handle persistent and transient objects. 
    --   It is the Standard run-time encapsulation of the CAS.CADE 
    --   database, that is, it defines a single programming interface 
    --   for creating and accessing persistent objects manipulated by 
    --   handles.


is
    enumeration InternalType is
    	    	Void,          -- TYPUND     0x00000000  /* Undefined    */
		Char,          -- TYPIT1     0x00010001  /* Byte         */
		ExtChar,       -- TYPIT2     0x00020001  /* Integer*2    */
		LongInt,       -- TYPIT4     0x00040001  /* Integer*4    */
		Bool,          -- TYPLO4     0x00040002  /* Logical*4    */
		Float,         -- TYPRE4     0x00040004  /* Real*4       */
		LongDouble,    -- TYPRE8     0x00080004  /* Real*8       */
		String,        -- TYPCHR     0x00000010  /* Character    */
		EString,       -- TYPCHREXT  0x00000011  /* Character    */
		EntryAddress,  -- TYPENT     0x00040020	 /* Function address */
		DataAddress,   -- TYPDAD     0x00040080  /* Data address */
		EngineHandle,  -- TYPHDLE    0x00004000  /* Handle       */
		Long64,        -- TYPIT8     0x00080001  /* Integer*8    */
		Array;         -- TYPARR     0x00008000  /* Tableau      */

    enumeration WayOfLife is IsNothing, IsAddress, IsTransient, IsPersistent, IsNotLoaded;
    enumeration KindOfType is IsUnKnown, IsClass, IsEnumeration, IsPrimitive, IsImported, IsPackage;
    enumeration HandlerStatus is HandlerVoid, HandlerJumped, HandlerProcessed;

    imported IStream;
    imported OStream;
    imported SStream;
    imported UUID;
    imported JmpBuf;
    imported ThreadId;

    primitive CString;
    primitive ExtString;
    primitive Address;
    primitive Size;
    primitive PByte;
    primitive PCharacter;
    primitive PExtCharacter;

    primitive Utf8Char;
    primitive Utf16Char;
    primitive Utf32Char;
    primitive WideChar;

    deferred class ErrorHandlerCallback;
    class ErrorHandler;
    
    class AncestorIterator;
    
    primitive Boolean;
    primitive Character;
    primitive ExtCharacter;
    primitive Integer;
    primitive Byte;
    primitive Real;
    primitive ShortReal;
    primitive Time;
    primitive OId;
    
    class GUID;

    deferred class Persistent ;

    deferred class Transient ;
   	    class Type; -- inherits Transient
    	    class Failure; --  inherits Transient
    	    	exception AbortiveTransaction inherits Failure;
	        exception DomainError inherits Failure;
    	    	    exception ConstructionError inherits DomainError;
    	    	    exception NullObject inherits DomainError;
		    exception NoSuchObject inherits DomainError;
		    exception NoMoreObject inherits DomainError;
		    exception ImmutableObject inherits DomainError;
		    exception TypeMismatch inherits DomainError;
		    exception MultiplyDefined inherits DomainError;
		    exception DimensionError inherits DomainError;
			exception DimensionMismatch inherits DimensionError;
		    exception RangeError inherits DomainError;
			exception OutOfRange inherits RangeError;
			exception NullValue inherits RangeError;
			exception NegativeValue inherits RangeError;
    	    	exception NumericError inherits Failure;
    	    	    exception Underflow inherits NumericError;
    	    	    exception Overflow inherits NumericError;
    	    	    exception DivideByZero inherits NumericError;
    	    	exception ProgramError inherits Failure;
    	    	    exception NotImplemented inherits ProgramError;
    	    	    exception OutOfMemory inherits ProgramError;
    	    	exception LicenseError inherits Failure;
    	    	    exception LicenseNotFound inherits LicenseError;
    	    	    exception TooManyUsers inherits LicenseError;

    pointer PErrorHandler  to ErrorHandler; 
    
    
    -- 
    --  Mutex: a class to synchronize access to shared data 
    --  from threads within one process
    --
    imported Mutex;
    
    -- 
    --  Memory manager  
    --
    Allocate (aSize: Size from Standard)  
    	returns Address from Standard; 
    ---Purpose:  Allocates memory blocks  
    --           aSize - bytes to  allocate 
    
    Free (aStorage: Address from Standard); 
    ---Purpose:  Deallocates memory blocks
    --           aStorage - previously allocated memory block to be freed

    ---C++: alias "template <typename T> static inline void Free (T*& thePtr) { Free ((void*)thePtr); thePtr = 0; }"

    Reallocate(aStorage: Address from Standard;
               aNewSize: Size from Standard)  
    	returns Address from Standard; 
    ---Purpose:  Reallocates memory blocks 
    --           aStorage - previously allocated memory block 
    --           aNewSize - new size in bytes 

    AllocateAligned (theSize  : Size from Standard;
                     theAlign : Size from Standard)
    returns Address from Standard;
    ---Purpose:  Allocates aligned memory blocks.
    -- Should be used with CPU instructions which require specific alignment.
    -- For example: SSE requires 16 bytes, AVX requires 32 bytes.
    -- @param theSize  bytes to allocate
    -- @param theAlign alignment in bytes

    FreeAligned (thePtrAligned : Address from Standard);
    ---Purpose:  Deallocates memory blocks
    -- @param thePtrAligned the memory block previously allocated with AllocateAligned()
    ---C++: alias "template <typename T> static inline void FreeAligned (T*& thePtrAligned) { FreeAligned ((void* )thePtrAligned); thePtrAligned = 0; }"

    Purge returns Integer from Standard; 
    ---Purpose:  Deallocates the storage retained on the free list 
    --           and clears the list. 
    --           Returns non-zero if some memory has been actually freed.

end Standard;
