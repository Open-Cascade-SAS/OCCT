-- File:        AdvancedBrepShapeRepresentation.cdl
-- Created:     Mon Dec  4 12:02:22 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWAdvancedBrepShapeRepresentation from RWStepShape

	---Purpose : Read & Write Module for AdvancedBrepShapeRepresentation

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     AdvancedBrepShapeRepresentation from StepShape,
     EntityIterator from Interface

is

	Create returns RWAdvancedBrepShapeRepresentation;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable AdvancedBrepShapeRepresentation from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : AdvancedBrepShapeRepresentation from StepShape);

	Share(me; ent : AdvancedBrepShapeRepresentation from StepShape; iter : in out EntityIterator);

end RWAdvancedBrepShapeRepresentation;
