-- File:	MeshAlgo_Edge.cdl
-- Created:	Tue May 11 16:38:19 1993
-- Author:	Didier PIFFAULT
--		<dpf@nonox>
---Copyright:	 Matra Datavision 1993

-- signature
deferred class Edge from MeshAlgo 

	---Purpose: Describes the data structure of a Edge.


uses    Integer from Standard,
    	Boolean from Standard,
    	DegreeOfFreedom from MeshDS


is      Initialize     (node1, node2 : Integer from Standard;
    	    	    	canMove      : DegreeOfFreedom from MeshDS);
        ---Purpose: Contructs an Edge beetween to vertices.


    	FirstNode     (me)
        ---Purpose: Give the index of first node of the Edge.
    	    	    returns Integer from Standard;

    	LastNode      (me)
        ---Purpose: Give the index of Last node of the Edge.
    	    	    returns Integer from Standard;

	Movability     (me)
    	    returns DegreeOfFreedom from MeshDS;

	SetMovability     (me      : in out;
    	    	    	   canMove : DegreeOfFreedom from MeshDS);

	SameOrientation(me; Other : Edge from MeshAlgo)
	    returns Boolean from Standard;


---Purpose: For maping the Edges.
--          Same Edge -> Same HashCode
--          Different Edges -> Not IsEqual but can have same HashCode 

    	HashCode      (me;
    	    	       Upper : Integer from Standard)
	---C++: function call
    	        returns Integer from Standard;
		    
    	IsEqual       (me; Other: Edge from MeshAlgo)
	    ---C++: alias operator ==
    	    	    returns Boolean from Standard;

end Edge;
