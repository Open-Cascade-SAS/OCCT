-- Created by: Peter KURNEV
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ShellSplitter from BOPAlgo 
    	inherits Algo from BOPAlgo 
	 
	---Purpose:  
        -- The class provides the splitting of the set of connected faces 
	-- on separate loops    
uses   
    BaseAllocator from BOPCol, 
    Shape from TopoDS,
    ListOfShape from BOPCol, 
    ConnexityBlock from BOPTools, 
    ListOfConnexityBlock from BOPTools 
    
    
--raises

is 
    Create 
    	returns ShellSplitter from BOPAlgo; 
    ---C++: alias "Standard_EXPORT virtual ~BOPAlgo_ShellSplitter();" 
    ---Purpose: empty constructor
     
    Create(theAllocator: BaseAllocator from BOPCol)  
    	returns ShellSplitter from BOPAlgo; 
    ---Purpose:  constructor 
    
    AddStartElement(me:out; 
    	    theS: Shape from TopoDS); 
    ---Purpose: adds a face <theS> to process 	           
    
    StartElements(me)  
    	returns ListOfShape from BOPCol;
    ---C++: return const & 
    ---Purpose: return the faces to process 
    
    Perform(me:out) 
	is redefined;  
    ---Purpose: performs the algorithm 	
	  
    Shells(me) 
	returns ListOfShape from BOPCol; 
    ---C++: return const & 	 
    ---Purpose: returns the loops 
     
    MakeConnexityBlocks(me:out)  
    	is protected;  
     
    MakeShells (me:out)  
    	is protected;   
	
    SplitBlock(myclass; 
    	    theCB:out ConnexityBlock from BOPTools);  
        
fields  
    myStartShapes: ListOfShape from BOPCol is protected; 
    myShells: ListOfShape from BOPCol is protected; 
    myLCB   : ListOfConnexityBlock from BOPTools is protected; 
   
end ShellSplitter;
