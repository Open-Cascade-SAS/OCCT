-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class FillAreaStyle from StepVisual 

inherits TShared from MMgt

uses

	HAsciiString from TCollection, 
	HArray1OfFillStyleSelect from StepVisual, 
	FillStyleSelect from StepVisual
is

	Create returns mutable FillAreaStyle;
	---Purpose: Returns a FillAreaStyle

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aFillStyles : mutable HArray1OfFillStyleSelect from StepVisual) is virtual;

	-- Specific Methods for Field Data Access --

	SetName(me : mutable; aName : mutable HAsciiString);
	Name (me) returns mutable HAsciiString;
	SetFillStyles(me : mutable; aFillStyles : mutable HArray1OfFillStyleSelect);
	FillStyles (me) returns mutable HArray1OfFillStyleSelect;
	FillStylesValue (me; num : Integer) returns FillStyleSelect;
	NbFillStyles (me) returns Integer;

fields

	name : HAsciiString from TCollection;
	fillStyles : HArray1OfFillStyleSelect from StepVisual; -- a SelectType

end FillAreaStyle;
