-- Created on: 1993-04-06
-- Created by: Philippe DAUTRY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class CartesianPoint from PGeom2d inherits Point from PGeom2d

        ---Purpose : Point defined  in  3D space with its 3  cartesian
        --         coordinates X, Y, Z.
        --         
    	---See Also : CartesianPoint from Geom2d.

uses Pnt2d from gp

is


  Create returns mutable CartesianPoint from PGeom2d;
        ---Purpose : Returns a CartesianPoint with default values..
	---Level: Internal 


  Create (aPnt2d : Pnt2d from gp) returns mutable CartesianPoint from PGeom2d;
        ---Purpose : Returns a CartesianPoint built with <aPnt2d>.
	---Level: Internal 


  Pnt (me : mutable; aPnt2d : Pnt2d from gp);
        ---Purpose : Set the field Pnt2d.
	---Level: Internal 


  Pnt (me)  returns Pnt2d;
        ---Purpose : Returns the value of the field Pnt2d.
	---Level: Internal 


fields

    pnt : Pnt2d from gp;

end;
