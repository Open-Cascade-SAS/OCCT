-- File:	RWStepDimTol_RWSymmetryTolerance.cdl
-- Created:	Wed Jun  4 13:34:34 2003 
-- Author:	Galina KULIKOVA
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWSymmetryTolerance from RWStepDimTol

    ---Purpose: Read & Write tool for SymmetryTolerance

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    SymmetryTolerance from StepDimTol

is
    Create returns RWSymmetryTolerance from RWStepDimTol;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : SymmetryTolerance from StepDimTol);
	---Purpose: Reads SymmetryTolerance

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: SymmetryTolerance from StepDimTol);
	---Purpose: Writes SymmetryTolerance

    Share (me; ent : SymmetryTolerance from StepDimTol;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWSymmetryTolerance;
