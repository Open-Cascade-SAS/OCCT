-- Created on: 1994-04-21
-- Created by: s:	Christophe GUYOT & Frederic UNTEREINER
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class TopoSurface  from IGESToBRep inherits CurveAndSurface from IGESToBRep

    ---Purpose : Provides methods to transfer topologic surfaces entities 
    --           from IGES to CASCADE.

uses   

    CurveAndSurface      from IGESToBRep,
    IGESEntity           from IGESData,
    RuledSurface         from IGESGeom,
    SurfaceOfRevolution  from IGESGeom,
    TabulatedCylinder    from IGESGeom,
    OffsetSurface        from IGESGeom,
    Plane                from IGESGeom,
    TrimmedSurface       from IGESGeom,
    BoundedSurface       from IGESGeom,
    PlaneSurface         from IGESSolid,
    SingleParent         from IGESBasic,
    Shape                from TopoDS,
    Face                 from TopoDS,
    Pln                  from gp,
    Trsf                 from gp,
    Trsf2d               from gp


is

    Create returns TopoSurface;
    ---Purpose : Creates  a tool TopoSurface  ready  to  run, with
    --         epsilons  set  to  1.E-04,  TheModeTopo  to  True,  the
    --         optimization of  the continuity to False.

    Create(CS : CurveAndSurface from IGESToBRep) returns TopoSurface;
    ---Purpose : Creates a tool TopoSurface ready to run and sets its
    --         fields as CS's.

    Create(eps        : Real;
    	   epsGeom    : Real;
    	   epsCoeff   : Real;
    	   mode       : Boolean; 
	   modeapprox : Boolean; 
    	   optimized  : Boolean)
        returns TopoSurface;
    ---Purpose : Creates a tool TopoSurface ready to run.

    TransferTopoSurface         (me    : in out;
    	    	    	    	 start : IGESEntity from IGESData)
    	returns Shape from TopoDS;
	
    TransferTopoBasicSurface    (me    : in out;
    	    	    	    	 start : IGESEntity from IGESData)
    	returns Shape from TopoDS;
	
    TransferRuledSurface        (me    : in out;
    	    	    	    	 start : RuledSurface from IGESGeom)
    	returns Shape from TopoDS;
	
    TransferSurfaceOfRevolution (me    : in out;
    	    	    	    	 start : SurfaceOfRevolution from IGESGeom)
    	returns Shape from TopoDS;

    TransferTabulatedCylinder   (me    : in out;
    	    	    	         start : TabulatedCylinder from IGESGeom)
    	returns Shape from TopoDS;

    TransferOffsetSurface       (me    : in out;
    	    	    	         start : OffsetSurface from IGESGeom)
    	returns Shape from TopoDS;

    TransferTrimmedSurface      (me    : in out;
    	    	    	         start : TrimmedSurface from IGESGeom)
    	returns Shape from TopoDS;

    TransferBoundedSurface      (me    : in out;
    	    	    	         start : BoundedSurface from IGESGeom)
    	returns Shape from TopoDS;

    TransferPlane               (me    : in out;
    	    	    	         start : Plane from IGESGeom)
    	returns Shape from TopoDS;

    TransferPlaneSurface        (me    : in out;
    	    	    	         start : PlaneSurface from IGESSolid)
    	returns Shape from TopoDS;

    TransferPerforate           (me    : in out;
                                 start : SingleParent from IGESBasic)
        returns Shape from TopoDS;

    TransferPlaneParts          (me    : in out;
                                 start : Plane from IGESGeom;
                                 gplan : out Pln  from gp;
                                 locat : out Trsf from gp;
                                 first : Boolean)
        returns Shape from TopoDS  is private;

    ParamSurface                (me      : in out;
    	    	    	    	 start   : IGESEntity from IGESData;
				 trans   : out Trsf2d from gp;
				 uFact   : out Real)
    	returns Shape from TopoDS;
    --             ---Purpose : Set the surface parameters:
    --           IsRevol : True for TabulatedCylinder or SurfaceOfRevolution
    --           ParamU ,Paramv, Length used for 2d Curves parametrization.
    
fields

    TheULength : Real from Standard;
    
end TopoSurface;
