-- Created on: 1993-01-27
-- Created by: Philippe DAUTRY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred generic class Iterator from Sweep (TheShape as any)

	---Purpose: This  is a  signature class describing   iteration
	--          services   required      by the Swept   Primitives
	--          algorithms from  a Directing or a Generating Line.
	--          This  tool is  used   to  iterate   on the  direct
	--          sub-shapes  of a  Shape. 
	--          

uses

    Orientation from TopAbs

raises

    NoMoreObject from Standard,
    NoSuchObject from Standard

is

    Init(me : in out; aShape: TheShape)
	---Purpose: Resest the Iterator on sub-shapes of <aShape>.
    is deferred;
    
    More(me) returns Boolean
	---Purpose: Returns True if there is a current sub-shape.
	--          
	-- -C++: inline
    is deferred;
    
    Next(me : in out)
	---Purpose: Moves to the next sub-shape.
    raises
    	NoMoreObject from Standard
    is deferred;
    
    Value(me) returns TheShape
	---Purpose: Returns the current sub-shape.
    raises
    	NoSuchObject from Standard
	-- -C++: return const &
	-- -C++: inline
    is deferred;
    
    Orientation(me) returns Orientation from TopAbs
	---Purpose: Returns the orientation of the current sub-shape.
    raises
    	NoSuchObject from Standard
	---C++: return const &
	---C++: inline
    is deferred;
    
end Iterator;
