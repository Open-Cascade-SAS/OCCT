-- Created on: 1997-02-10
-- Created by: Odile Olivier
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


--  SAV : OCC218 06/03/02 : Add(...) overloaded to take into account arrow & text
--                          aspects.

class XYZAxisPresentation from DsgPrs
    	---Purpose: A framework for displaying the axes of an XYZ trihedron.
uses

    Presentation from Prs3d,
    LineAspect   from Prs3d,
    Pnt          from gp,
    Dir          from gp,
    ArrowAspect from Prs3d,
    TextAspect from Prs3d

is

    Add(myclass;
    	aPresentation: Presentation from Prs3d;
    	anLineAspect : LineAspect from Prs3d;
    	aDir         : Dir from gp;
	aVal         : Real from Standard;
	aText        : CString from Standard;
    	aPfirst      : Pnt    from gp;
    	aPlast       : Pnt    from gp);
	 
    	---Purpose: Draws each axis of a trihedron displayed in the
    	-- presentation aPresentation and with lines shown by
    	-- the values of aLineAspect. Each axis is defined by:
    	-- -   the first and last points aPfirst and aPlast
    	-- -   the direction aDir and
    	-- -   the value aVal which provides a value for length.
    	--  The value for length is provided so that the trihedron
    	-- can vary in length relative to the scale of shape display.
    	-- Each axis will be identified as X, Y, or Z by the text aText.


    Add(myclass;
    	aPresentation : Presentation from Prs3d;
    	aLineAspect   : LineAspect from Prs3d;
    	anArrowAspect : ArrowAspect from Prs3d;
    	aTextAspect   : TextAspect from Prs3d;
    	aDir          : Dir from gp;
	aVal          : Real from Standard;
	aText         : CString from Standard;
    	aPfirst       : Pnt    from gp;
    	aPlast        : Pnt    from gp);
	 
    	---Purpose: draws the presentation X ,Y ,Z axis

end XYZAxisPresentation;
