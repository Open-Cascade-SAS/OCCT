-- Created on: 1994-12-16
-- Created by: Frederic MAUPAS
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class TranslateEdge from StepToTopoDS
    inherits Root from StepToTopoDS
    
    ---Purpose:
    --         

uses

    Edge               from StepShape,
    Tool               from StepToTopoDS,
    TranslateEdgeError from StepToTopoDS,
    Shape              from TopoDS,
    Edge               from TopoDS,
    Vertex             from TopoDS,
    Curve              from Geom2d,
    Surface            from Geom,
    EdgeCurve          from StepShape,
    Curve              from StepGeom,
    Vertex             from StepShape,
    Pcurve             from StepGeom,
    NMTool             from StepToTopoDS

raises NotDone from StdFail

is

    Create returns TranslateEdge;
    
    Create (E      : Edge from StepShape;
            T      : in out Tool from StepToTopoDS;
            NMTool : in out NMTool from StepToTopoDS)
    	returns TranslateEdge;
	    
    Init (me     : in out;
          E      : Edge from StepShape;
          T      : in out Tool from StepToTopoDS;
          NMTool : in out NMTool from StepToTopoDS);

    MakeFromCurve3D (me : in out; C3D : Curve from StepGeom;
    	    	     EC     : EdgeCurve from StepShape;        -- for messages
		     Vend   : Vertex from StepShape;      -- case of null edge
		     preci  : Real; E : in out Edge from TopoDS;
		     V1, V2 : in out Vertex from TopoDS;
		     T      : in out Tool from StepToTopoDS);
    ---Purpose:  Warning! C3D is assumed to be a Curve 3D ...
    --    other cases to checked before calling this

    MakePCurve (me; PCU : Pcurve from StepGeom; ConvSurf : Surface from Geom)
    	returns Curve from Geom2d;
    --  Null if failed

    Value (me) returns Shape from TopoDS
    	raises NotDone
	is static;
	---C++: return const &

    Error (me) returns TranslateEdgeError from StepToTopoDS;
    
fields

    myError  : TranslateEdgeError from StepToTopoDS;
    
    myResult : Shape              from TopoDS;
    
end TranslateEdge;
