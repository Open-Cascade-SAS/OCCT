-- Created on: 1992-09-28
-- Created by: Remi GILET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class MakeArcOfHyperbola from GC inherits Root from GC
    	---Purpose: Implements construction algorithms for an arc
    	-- of hyperbola in 3D space. The result is a Geom_TrimmedCurve curve.
    	-- A MakeArcOfHyperbola object provides a framework for:
    	-- -   defining the construction of the arc of hyperbola,
    	-- -   implementing the construction algorithm, and
    	-- -   consulting the results. In particular, the
    	--   Value function returns the constructed arc of hyperbola.
        
uses Pnt          from gp,
     Hypr         from gp,
     Dir          from gp,
     Ax1          from gp,
     Real         from Standard,
     TrimmedCurve from Geom

raises NotDone from StdFail

is

Create(Hypr           : Hypr    from gp       ;
       Alpha1, Alpha2 : Real    from Standard ;
       Sense          : Boolean from Standard ) returns MakeArcOfHyperbola;
    	---Purpose: Creates an arc of Hyperbola (TrimmedCurve from Geom) from 
    	--          a Hyperbola between two parameters Alpha1 and Alpha2
    	--          (given in radians).

Create(Hypr  : Hypr    from gp       ;
       P     : Pnt     from gp       ;
       Alpha : Real    from Standard ;
       Sense : Boolean from Standard ) returns MakeArcOfHyperbola;
    	---Purpose: Creates an arc of Hyperbola (TrimmedCurve from Geom) from 
    	--          a Hyperbola between point <P> and the parameter
        --          Alpha (given in radians).

Create(Hypr  : Hypr    from gp ;
       P1    : Pnt     from gp ;
       P2    : Pnt     from gp ;
       Sense : Boolean from Standard ) returns MakeArcOfHyperbola;
    	---Purpose: Creates an arc of Hyperbola (TrimmedCurve from Geom) from 
    	--          a Hyperbola between two points P1 and P2.
    	-- The orientation of the arc of hyperbola is:
    	-- -   the sense of Hypr if Sense is true, or
    	-- -   the opposite sense if Sense is false.
    
Value(me) returns TrimmedCurve from Geom
    raises NotDone
    is static;
    	--- Purpose: Returns the constructed arc of hyperbola.
    	---C++: return const&

Operator(me) returns TrimmedCurve from Geom
    is static;
    	---C++: return const&
    	---C++: alias "Standard_EXPORT operator Handle_Geom_TrimmedCurve() const;"

fields

    TheArc : TrimmedCurve from Geom;
    --The solution from Geom.
    
end MakeArcOfHyperbola;
