-- Created on: 1997-04-17
-- Created by: Christophe MARION
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class EdgeInterferenceTool from HLRBRep

	---Purpose: Implements the  methods required  to  instantiates
	--          the EdgeInterferenceList from HLRAlgo.

uses
    Integer      from Standard,
    Boolean      from Standard,
    Real         from Standard,
    Dir          from gp,
    Orientation  from TopAbs,
    Intersection from HLRAlgo,
    Interference from HLRAlgo,
    Data         from HLRBRep

is
    Create(DS : Data from HLRBRep) returns EdgeInterferenceTool from HLRBRep;

    --- methods to iterate on the Vertices of the Edge
    
    LoadEdge(me : in out)
    is static;
	
    InitVertices(me : in out)
	---C++: inline
    is static;
    
    MoreVertices(me) returns Boolean from Standard
	---C++: inline
    is static;
    
    NextVertex(me : in out)
	---C++: inline
    is static;
    
    CurrentVertex(me) returns Intersection from HLRAlgo
	---C++: inline
    	---C++: return const &
    is static;
    
    CurrentOrientation(me) returns Orientation from TopAbs
	---C++: inline
    is static;
    
    CurrentParameter(me) returns Real from Standard
	---C++: inline
    is static;
    
    -- Data on the Edge

    IsPeriodic(me) returns Boolean from Standard
	---C++: inline
    is static;

    EdgeGeometry(me; Param :     Real from Standard;
    	    	     Tgt   : out Dir  from gp;
		     Nrm   : out Dir  from gp;
		     Curv  : out Real from Standard)
	---Purpose: Returns local geometric description of the Edge at
	--          parameter   <Para>.  See  method  Reset  of  class
	--          EdgeFaceTransition from TopCnx for other arguments.
    is static;
    
    -- Data on Interferences
    
    ParameterOfInterference(me; I : Interference from HLRAlgo) 
    returns Real from Standard 
    	---C++: inline
    is static;
    
    SameInterferences(me; I1, I2 : Interference from HLRAlgo) 
    returns Boolean from Standard 
	---Purpose: True if   the  two interferences are on   the same
	--          geometric locus.
    is static;
    
    SameVertexAndInterference(me; I : Interference from HLRAlgo)
    returns Boolean from Standard
	---Purpose: True if the  Interference and the  current  Vertex
	--          are on the same geometric locus.
    is static;
    
    InterferenceBoundaryGeometry(me; I    :     Interference from HLRAlgo;
    	                             Tang : out Dir          from gp;       
   	                             Norm : out Dir          from gp;       
    	                             Curv : out Real         from Standard)
	---Purpose: Returns   the  geometry of  the   boundary  at the
	--          interference  <I>.  See the AddInterference method
	--          of the class  EdgeFaceTransition  from  TopCnx for
	--          the other arguments.
    is static;    	
    
fields
    myDS   : Data         from HLRBRep;
    inter  : Intersection from HLRAlgo [2];
    cur    : Integer      from Standard;
    
end EdgeInterferenceTool;
