-- Created on: 1994-03-17
-- Created by: Bruno DUMORTIER
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class ProjectPointOnSurf from GeomAPI

    	--- Purpose:
    	-- This class implements methods for  computing all the orthogonal
    	--  projections of a point onto a  surface. 

uses
    Surface   from Geom,
    ExtPS     from Extrema,
    ExtAlgo from Extrema,
    Pnt       from gp,
    Length    from Quantity,
    Parameter from Quantity,
--modified by NIZNHY-PKV Thu Apr  4 10:37:24 2002  f
    Surface from GeomAdaptor 
--modified by NIZNHY-PKV Thu Apr  4 10:37:28 2002  t
raises
    OutOfRange from Standard,
    NotDone    from StdFail
    
    
is

    Create
	---Purpose: Creates an empty object. Use the
    	-- Init function for further initialization.          
    returns ProjectPointOnSurf from GeomAPI;
    
    
    Create(P          : Pnt     from gp;
    	   Surface    : Surface from Geom;
    	   Algo : ExtAlgo from Extrema = Extrema_ExtAlgo_Grad)
        ---Purpose: Create the projection  of a point <P> on a surface
        --          <Surface> 
	---Level: Public          
    returns ProjectPointOnSurf from GeomAPI;

    Create(P          : Pnt     from gp;
    	   Surface    : Surface from Geom;
    	   Tolerance  : Real    from Standard;
    	   Algo : ExtAlgo from Extrema = Extrema_ExtAlgo_Grad)
        ---Purpose: Create the projection  of a point <P> on a surface
        --          <Surface> 
	---Level: Public          
    returns ProjectPointOnSurf from GeomAPI;
    

        ---Purpose: Create the projection of a point <P>  on a surface
        --          <Surface>. The solution are computed in the domain
        --          [Umin,Usup] [Vmin,Vsup] of the surface.
	---Level: Public          

    Create(P          : Pnt       from gp;
    	   Surface    : Surface   from Geom;
    	   Umin, Usup, 
    	   Vmin, Vsup : Parameter from Quantity;
           Tolerance  : Real      from Standard;
    	   Algo : ExtAlgo from Extrema = Extrema_ExtAlgo_Grad)
    returns ProjectPointOnSurf from GeomAPI;

    Create(P          : Pnt       from gp;
    	   Surface    : Surface   from Geom;
    	   Umin, Usup, 
    	   Vmin, Vsup : Parameter from Quantity;
    	   Algo : ExtAlgo from Extrema = Extrema_ExtAlgo_Grad)
    returns ProjectPointOnSurf from GeomAPI;


        ---Purpose: Init the projection  of a point <P> on a surface
        --          <Surface> 
	---Level: Public          

    Init(me : in out;
    	 P          : Pnt     from gp;
	 Surface    : Surface from Geom;
    	 Tolerance  : Real    from Standard;
    	 Algo : ExtAlgo from Extrema = Extrema_ExtAlgo_Grad)
    is static;

    Init(me : in out;
    	 P          : Pnt     from gp;
	 Surface    : Surface from Geom;
	 Algo : ExtAlgo from Extrema = Extrema_ExtAlgo_Grad)
    is static;


        ---Purpose: Init the projection of a point <P>  on a surface
        --          <Surface>. The solution are computed in the domain
        --          [Umin,Usup] [Vmin,Vsup] of the surface.
	---Level: Public          

    Init(me : in out;
    	 P          : Pnt       from gp;
	 Surface    : Surface   from Geom;
    	 Umin, Usup, 
    	 Vmin, Vsup : Parameter from Quantity;
    	 Tolerance  : Real    from Standard;
    	 Algo : ExtAlgo from Extrema = Extrema_ExtAlgo_Grad)
	---Level: Public          
    is static;

    Init(me : in out;
    	 P          : Pnt       from gp;
	 Surface    : Surface   from Geom;
    	 Umin, Usup, 
    	 Vmin, Vsup : Parameter from Quantity;
    	 Algo : ExtAlgo from Extrema = Extrema_ExtAlgo_Grad)
    is static;


        ---Purpose: Init the projection for many points on a surface
        --          <Surface>. The solutions will be computed in the domain
        --          [Umin,Usup] [Vmin,Vsup] of the surface.
	---Level: Public          

    Init(me : in out;
	 Surface    : Surface   from Geom;
    	 Umin, Usup, 
    	 Vmin, Vsup : Parameter from Quantity;
	 Tolerance  : Real      from Standard;
	 Algo : ExtAlgo from Extrema = Extrema_ExtAlgo_Grad)
    is static;

    Init(me : in out;
	 Surface    : Surface   from Geom;
    	 Umin, Usup, 
    	 Vmin, Vsup : Parameter from Quantity;
    	 Algo : ExtAlgo from Extrema = Extrema_ExtAlgo_Grad)
    is static;


    Perform (me: in out; P: Pnt from gp)
    	---Purpose: Performs the projection of a point on the current surface.
    	---Level : Public.
    is static;


    IsDone (me) returns Boolean from Standard is static;


    NbPoints(me)
	---Purpose: Returns the number of computed orthogonal projection points.
    	-- Note: if projection fails, NbPoints returns 0.
    returns Integer	
    	---C++: alias "Standard_EXPORT operator Standard_Integer() const;"
    is static;

    
    Point(me; Index : Integer from Standard)
	---Purpose: Returns the orthogonal projection
    	-- on the surface. Index is a number of a computed point.
    	-- Exceptions
    	-- Standard_OutOfRange if Index is not in the range [ 1,NbPoints ], where
    	-- NbPoints is the number of solution points.        
    returns Pnt from gp
    raises OutOfRange from Standard
	
    is static;
    
    
    Parameters(me; Index :     Integer   from Standard;
                   U, V  : out Parameter from Quantity)
        ---Purpose: Returns the parameters (U,V) on the
    	-- surface of the orthogonal projection. Index is a number of a
    	-- computed point.
    	-- Exceptions
    	-- Standard_OutOfRange if Index is not in the range [ 1,NbPoints ], where
    	-- NbPoints is the number of solution points.        
    raises OutOfRange from Standard
	
    is static;
    
    
    Distance(me; Index : Integer from Standard)
    returns Length from Quantity
	---Purpose: Computes the distance between the
    	-- point and its orthogonal projection on the surface. Index is a number
    	-- of a computed point.
    	-- Exceptions
    	-- Standard_OutOfRange if Index is not in the range [ 1,NbPoints ], where
    	-- NbPoints is the number of solution points.     
    raises OutOfRange from Standard
	
    is static;


    NearestPoint(me)
	---Purpose: Returns the nearest orthogonal projection of the point
    	-- on the surface.
    	-- Exceptions
    	-- StdFail_NotDone if projection fails.       
    returns Pnt from gp	
    	---C++: alias "Standard_EXPORT operator gp_Pnt() const;"
    raises NotDone from StdFail
    is static;
    
    
    LowerDistanceParameters(me; U, V : out Parameter from Quantity)
	---Purpose: Returns the parameters (U,V) on the
    	-- surface of the nearest computed orthogonal projection of the point.
    	-- Exceptions
    	-- StdFail_NotDone if projection fails.      
    raises NotDone from StdFail
    is static;


    LowerDistance(me)
	---Purpose: Computes the distance between the
    	-- point and its nearest orthogonal projection on the surface. 
    	-- Exceptions
    	-- StdFail_NotDone if projection fails.        
    returns Length from Quantity
 	---C++: alias "Standard_EXPORT operator Standard_Real() const;"
   raises NotDone from StdFail
    is static;
    
    
    Extrema(me)
	---Purpose: return the algorithmic object from Extrema
	---Level: Advanced
	---C++: return const&
	---C++: inline      
    returns ExtPS from Extrema
    is static;
	    

    Init(me : in out) is static private;
    	---Level: Private

fields

    myIsDone : Boolean from Standard;
    myIndex  : Integer from Standard;    -- index of the nearest solution
    myExtPS  : ExtPS   from Extrema; 
--modified by NIZNHY-PKV Thu Apr  4 10:36:31 2002  f 
    myGeomAdaptor:  Surface from GeomAdaptor; 
--modified by NIZNHY-PKV Thu Apr  4 10:36:33 2002  t
end ProjectPointOnSurf;
