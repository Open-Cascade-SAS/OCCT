-- Created on: 1996-03-08
-- Created by: Robert COUBLANC
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class FaceFilter from StdSelect inherits Filter from SelectMgr

	---Purpose: A framework to define a filter to select a specific type of face.
    	-- The types available include:
    	-- -   any face
    	-- -   a planar face
    	-- -   a cylindrical face
    	-- -   a spherical face
    	-- -   a toroidal face
    	-- -   a revol face.

uses
    TypeOfFace from StdSelect,
    Shape from TopoDS,
    EntityOwner from SelectMgr,
    ShapeEnum from TopAbs
is

    Create (aTypeOfFace: TypeOfFace from StdSelect)
    returns FaceFilter from StdSelect;
    	---Purpose: Constructs a face filter object defined by the type of face aTypeOfFace.    
    SetType(me:mutable;aNewType : TypeOfFace from StdSelect);  
    	--- Purpose: Sets the type of face aNewType. aNewType is to be highlighted in selection.   
    Type(me) returns TypeOfFace from StdSelect;
    	--- Purpose: Returns the type of face to be highlighted in selection.   
    IsOk (me;anobj : EntityOwner from SelectMgr) 
    returns Boolean from Standard is redefined virtual;
  
    ActsOn(me; aStandardMode : ShapeEnum from TopAbs)
    returns Boolean from Standard is redefined virtual;
   
fields

    mytype : TypeOfFace from StdSelect;

end FaceFilter;
