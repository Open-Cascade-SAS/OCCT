-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ContextDependentOverRidingStyledItem from StepVisual 

inherits OverRidingStyledItem from StepVisual 

uses

	HArray1OfStyleContextSelect from StepVisual, 
	StyleContextSelect from StepVisual, 
	HAsciiString from TCollection, 
	HArray1OfPresentationStyleAssignment from StepVisual, 
	RepresentationItem from StepRepr, 
	StyledItem from StepVisual
is

	Create returns mutable ContextDependentOverRidingStyledItem;
	---Purpose: Returns a ContextDependentOverRidingStyledItem


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aStyles : mutable HArray1OfPresentationStyleAssignment from StepVisual;
	      aItem : mutable RepresentationItem from StepRepr;
	      aOverRiddenStyle : mutable StyledItem from StepVisual) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aStyles : mutable HArray1OfPresentationStyleAssignment from StepVisual;
	      aItem : mutable RepresentationItem from StepRepr;
	      aOverRiddenStyle : mutable StyledItem from StepVisual;
	      aStyleContext : mutable HArray1OfStyleContextSelect from StepVisual) is virtual;

	-- Specific Methods for Field Data Access --

	SetStyleContext(me : mutable; aStyleContext : mutable HArray1OfStyleContextSelect);
	StyleContext (me) returns mutable HArray1OfStyleContextSelect;
	StyleContextValue (me; num : Integer) returns StyleContextSelect;
	NbStyleContext (me) returns Integer;

fields

	styleContext : HArray1OfStyleContextSelect from StepVisual; -- a SelectType

end ContextDependentOverRidingStyledItem;
