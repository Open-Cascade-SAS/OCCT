-- File:	RWStepBasic_RWProductDefinitionRelationship.cdl
-- Created:	Mon Jul  3 19:47:51 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class RWProductDefinitionRelationship from RWStepBasic

    ---Purpose: Read & Write tool for ProductDefinitionRelationship

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    ProductDefinitionRelationship from StepBasic

is
    Create returns RWProductDefinitionRelationship from RWStepBasic;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : ProductDefinitionRelationship from StepBasic);
	---Purpose: Reads ProductDefinitionRelationship

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: ProductDefinitionRelationship from StepBasic);
	---Purpose: Writes ProductDefinitionRelationship

    Share (me; ent : ProductDefinitionRelationship from StepBasic;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWProductDefinitionRelationship;
