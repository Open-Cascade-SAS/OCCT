-- Created on: 1993-07-09
-- Created by: Isabelle GRIGNON
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Add2dCurve from BndLib
       	---Purpose: Computes the bounding box for a curve in 2d .
    	-- Functions to add a 2D curve to a bounding box.
    	-- The 2D curve is defined from a Geom2d curve.
        
uses Box2d   from Bnd,
     Curve2d from Adaptor2d


is

    Add(myclass; C   :        Curve2d from Adaptor2d;
    	    	 Tol :        Real    from Standard; 
    	    	 B   : in out Box2d   from Bnd);
    	---Purpose: Adds to the bounding box B the curve C
        --  B is then enlarged by the tolerance value Tol.
    	-- Note: depending on the type of curve, one of the following
    	-- representations of the curve C is used to include it in the bounding box B:
    	-- -   an exact representation if C is built from a line, a circle   or a conic curve,
    	-- -   the poles of the curve if C is built from a Bezier curve or   a BSpline curve,
    	-- -   if not, the points of an approximation of the curve C.
    	-- Warning
    	-- C is an adapted curve, that is, an object which is an interface between:
    	-- -   the services provided by a 2D curve from the package Geom2d
    	-- -   and those required of the curve by the computation algorithm.
    	--  The adapted curve is created in the following way:
    	--    Handle(Geom2d_Curve) mycurve = ...
    	-- ;
    	--    Geom2dAdaptor_Curve C(mycurve);
    	-- The bounding box B is then enlarged by adding it:
    	--    Bnd_Box2d B;
    	-- // ...
    	--    Standard_Real Tol = ... ;
    	--    Add2dCurve::Add ( C, Tol, B );
    	-- Exceptions
    	-- Standard_Failure if the curve is built from:
    	-- -   a Geom_Line, or
    	-- -   a Geom_Parabola, or
    	-- -   a Geom_Hyperbola,
    	-- and P1 and P2 are either two negative infinite real
    	-- numbers, or two positive infinite real numbers.
        
    Add(myclass; C       :        Curve2d from Adaptor2d;
    	    	 U1,U2   :        Real    from Standard;
    	         Tol     :        Real    from Standard; 
    	    	 B       : in out Box2d   from Bnd);
    	---Purpose: Adds to the bounding box Bthe arc of the curve C limited by the two parameter
    	--  values P1 and P2.
        --  B is then enlarged by the tolerance value Tol.
    	-- Note: depending on the type of curve, one of the following
    	-- representations of the curve C is used to include it in the bounding box B:
    	-- -   an exact representation if C is built from a line, a circle   or a conic curve,
    	-- -   the poles of the curve if C is built from a Bezier curve or   a BSpline curve,
    	-- -   if not, the points of an approximation of the curve C.
    	-- Warning
    	-- C is an adapted curve, that is, an object which is an interface between:
    	-- -   the services provided by a 2D curve from the package Geom2d
    	-- -   and those required of the curve by the computation algorithm.
    	--  The adapted curve is created in the following way:
    	--    Handle(Geom2d_Curve) mycurve = ...
    	-- ;
    	--    Geom2dAdaptor_Curve C(mycurve);
    	-- The bounding box B is then enlarged by adding it:
    	--    Bnd_Box2d B;
    	-- // ...
    	--    Standard_Real Tol = ... ;
    	--    Add2dCurve::Add ( C, Tol, B );
    	-- Exceptions
    	-- Standard_Failure if the curve is built from:
    	-- -   a Geom_Line, or
    	-- -   a Geom_Parabola, or
    	-- -   a Geom_Hyperbola,
    	-- and P1 and P2 are either two negative infinite real
    	-- numbers, or two positive infinite real numbers.      
        
        
end Add2dCurve;
