-- Created on: 2003-02-04
-- Created by: data exchange team
-- Copyright (c) 2003-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class ElementOrElementGroup from StepFEA
inherits SelectType from StepData

    ---Purpose: Representation of STEP SELECT type ElementOrElementGroup

uses
    ElementRepresentation from StepFEA,
    ElementGroup from StepFEA

is
    Create returns ElementOrElementGroup from StepFEA;
	---Purpose: Empty constructor

    CaseNum (me; ent: Transient) returns Integer;
	---Purpose: Recognizes a kind of ElementOrElementGroup select type
	--          1 -> ElementRepresentation from StepFEA
	--          2 -> ElementGroup from StepFEA
	--          0 else

    ElementRepresentation (me) returns ElementRepresentation from StepFEA;
	---Purpose: Returns Value as ElementRepresentation (or Null if another type)

    ElementGroup (me) returns ElementGroup from StepFEA;
	---Purpose: Returns Value as ElementGroup (or Null if another type)

end ElementOrElementGroup;
