-- Created on: 1993-01-11
-- Created by: CKY / Contract Toubro-Larsen ( Anand NATRAJAN )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class FlowLineSpec from IGESAppli  inherits IGESEntity

        ---Purpose: defines FlowLineSpec, Type <406> Form <14>
        --          in package IGESAppli
        --          Attaches one or more text strings to entities being
        --          used to represent a flow line

uses

        HAsciiString          from TCollection,
        HArray1OfHAsciiString from Interface

raises OutOfRange

is

        Create returns mutable FlowLineSpec;

        -- Specific Methods pertaining to the class

        Init (me : mutable; allProperties : HArray1OfHAsciiString);
        ---Purpose : This method is used to set the fields of the class
        --           FlowLineSpec
        --       - allProperties : primary flow line specification and modifiers

        NbPropertyValues (me) returns Integer;
        ---Purpose : returns the number of property values

        FlowLineName (me) returns HAsciiString from TCollection;
        ---Purpose : returns primary flow line specification name

        Modifier (me; Index : Integer) returns HAsciiString from TCollection
        raises OutOfRange;
        ---Purpose : returns specified modifier element
        -- raises exception if Index <= 1 or Index > NbPropertyValues

fields

--
-- Class    : IGESAppli_FlowLineSpec
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class FlowLineSpec.
--
-- Reminder : A FlowLineSpec instance is defined by :
--            - primary flow line specification name and modifiers

        theNameAndModifiers : HArray1OfHAsciiString;

end FlowLineSpec;
