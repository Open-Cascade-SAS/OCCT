-- Created on: 1993-01-11
-- Created by: CKY / Contract Toubro-Larsen ( Arun MENON )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PinNumber from IGESAppli  inherits IGESEntity

        ---Purpose: defines PinNumber, Type <406> Form <8>
        --          in package IGESAppli
        --          Used to attach a text string representing a component
        --          pin number to an entity being used to represent an
        --          electrical component's pin

uses

        HAsciiString from TCollection

is

        Create returns mutable PinNumber;

        -- Specific Methods pertaining to the class

        Init (me        : mutable;
              nbPropVal : Integer;
              aValue    : HAsciiString);
        ---Purpose : This method is used to set the fields of the class
        --           PinNumber
        --       - nbPropVal : Number of property values (always = 1)
        --       - aValue    : Pin Number value

        NbPropertyValues (me) returns Integer;
        ---Purpose : returns the number of property values
        -- is always 1

        PinNumberVal (me) returns HAsciiString from TCollection;
        ---Purpose : returns the pin number value

fields

--
-- Class    : IGESAppli_PinNumber
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class PinNumber.
--
-- Reminder : A PinNumber instance is defined by :
--            - Number of property values (always = 1)
--            - Pin Number value

        theNbPropertyValues : Integer;
        thePinNumber        : HAsciiString;

end PinNumber;
