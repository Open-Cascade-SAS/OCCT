-- Created on: 1993-11-26
-- Created by: Modelistation
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ALineToWLine from IntPatch

uses 
    WLine from IntPatch,
    ALine from IntPatch,
    Quadric from IntSurf

is 

    Create(Quad1 : Quadric from IntSurf;
    	   Quad2 : Quadric from IntSurf)
    
    	returns ALineToWLine from IntPatch;
	
    Create(Quad1       : Quadric from IntSurf;
           Quad2       : Quadric from IntSurf;
           Deflection  : Real from Standard;
    	   PasMaxUV    : Real from Standard;
           NbMaxPoints : Integer from Standard) 
    
    	returns ALineToWLine from IntPatch;
	
	
    SetTolParam(me:out; 
    	    aT:Real from Standard); 
	 
    TolParam(me) 
    	returns Real from Standard; 
	 
    SetTolOpenDomain(me:out; 
    	    aT:Real from Standard); 
	 
    TolOpenDomain(me) 
    	returns Real from Standard; 
	 
    SetTolTransition(me:out; 
    	    aT:Real from Standard); 
	 
    TolTransition(me) 
    	returns Real from Standard;  

    SetTol3D(me:out; 
    	    aT:Real from Standard); 
	 
    Tol3D(me) 
    	returns Real from Standard;  
     
    SetConstantParameter(me);
    
    SetUniformAbscissa(me);
    
    SetUniformDeflection(me);
    
    MakeWLine(me; aline: ALine from IntPatch)
    
    	returns WLine from IntPatch;
	
    MakeWLine(me; aline: ALine from IntPatch; paraminf,paramsup: Real from Standard)
    	returns WLine from IntPatch; 
    
fields
    quad1         : Quadric from IntSurf;
    quad2         : Quadric from IntSurf;
    deflectionmax : Real    from Standard;
    nbpointsmax   : Integer from Standard;
    type          : Integer from Standard; -- 0: Constant Parameter
                                           -- 1: Uniform Abscissa
                                           -- 2: Uniform Deflection
    myTolParam      : Real from Standard; 
    myTolOpenDomain : Real from Standard; 
    myTolTransition : Real from Standard; 
    myTol3D         : Real from Standard;        

end;
