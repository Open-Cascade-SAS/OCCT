-- Created on: 1992-11-18
-- Created by: Christian CAILLET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class SelectType  from IFSelect   inherits SelectAnyType

    ---Purpose : A SelectType keeps or rejects Entities of which the Type
    --           is Kind of a given Cdl Type

uses Type, AsciiString from TCollection, Transient

is

    Create returns mutable SelectType;
    ---Purpose : Creates a SelectType. Default is no filter

    Create (atype : Type) returns mutable SelectType;
    ---Purpose : Creates a SelectType for a given Type

    SetType (me : mutable; atype : Type);
    ---Purpose : Sets a TYpe for filter

    TypeForMatch (me) returns Type;
    ---Purpose : Returns the Type to be matched for select : this is the type
    --           given at instantiation time

    ExtractLabel (me) returns AsciiString from TCollection;
    ---Purpose : Returns a text defining the criterium.
    --           (should by gotten from Type of Entity used for instantiation)

fields

    thetype : Type;

end SelectType;
