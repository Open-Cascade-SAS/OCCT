-- File:	IGESDimen_ToolAngularDimension.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolAngularDimension  from IGESDimen

    ---Purpose : Tool to work on a AngularDimension. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses AngularDimension from IGESDimen,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolAngularDimension;
    ---Purpose : Returns a ToolAngularDimension, ready to work


    ReadOwnParams (me; ent : mutable AngularDimension;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : AngularDimension;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : AngularDimension;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a AngularDimension <ent>, from
    --           its specific (own) parameters

    DirChecker (me; ent : AngularDimension) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : AngularDimension;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : AngularDimension; entto : mutable AngularDimension;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : AngularDimension;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolAngularDimension;
