-- Created by: Sergey RUIN
-- Copyright (c) 2001-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class CompoundDelta from TDocStd inherits Delta from TDF

	---Purpose: A delta set is available at <aSourceTime>. If
	--          applied, it restores the TDF_Data in the state it
	--          was at <aTargetTime>.

uses

    OStream from Standard

is


    Create;
	---Purpose: Creates a compound delta.

--    SetValidTime(me : mutable;  aBeginTime, anEndTime : Integer from Standard) is private;
    ---Purpose: Validates <me> at <aBeginTime>. If applied, it
    --          restores the TDF_Data in the state it was at
    --          <anEndTime>. Reserved to TDF_Data.
    
--    AppendAttributeDelta(me : mutable; anAttributeDelta : AttributeDelta from TDF) is private;
    
friends

    class Document from TDocStd

end Delta;

