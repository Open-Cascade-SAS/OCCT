-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class AutoDesignDateAndTimeItem from StepAP214 inherits SelectType from StepData

	-- <AutoDesignDateAndTimeItem> is an EXPRESS Select Type construct translation.
	-- it gathers : ApprovalPersonOrganization, AutoDesignDateAndPersonAssignment

uses

	ApprovalPersonOrganization from StepBasic,
	AutoDesignDateAndPersonAssignment from StepAP214,
	ProductDefinitionEffectivity from StepBasic
is

	Create returns AutoDesignDateAndTimeItem;
	---Purpose : Returns a AutoDesignDateAndTimeItem SelectType

	CaseNum (me; ent : Transient) returns Integer;
	---Purpose: Recognizes a AutoDesignDateAndTimeItem Kind Entity that is :
	--        1 -> ApprovalPersonOrganization
	--        2 -> AutoDesignDateAndPersonAssignment
	--        0 else

	ApprovalPersonOrganization (me) returns any ApprovalPersonOrganization;
	---Purpose : returns Value as a ApprovalPersonOrganization (Null if another type)

	AutoDesignDateAndPersonAssignment (me) returns any AutoDesignDateAndPersonAssignment;
	---Purpose : returns Value as a AutoDesignDateAndPersonAssignment (Null if another type)

    	ProductDefinitionEffectivity (me) returns ProductDefinitionEffectivity;

end AutoDesignDateAndTimeItem;
