-- File:        ApprovalRelationship.cdl
-- Created:     Mon Dec  4 12:02:23 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWApprovalRelationship from RWStepBasic

	---Purpose : Read & Write Module for ApprovalRelationship

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     ApprovalRelationship from StepBasic,
     EntityIterator from Interface

is

	Create returns RWApprovalRelationship;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable ApprovalRelationship from StepBasic);

	WriteStep (me; SW : in out StepWriter; ent : ApprovalRelationship from StepBasic);

	Share(me; ent : ApprovalRelationship from StepBasic; iter : in out EntityIterator);

end RWApprovalRelationship;
