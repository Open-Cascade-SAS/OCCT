-- Created on: 1999-01-05
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Explorer from TopOpeBRepDS

uses

    Shape from TopoDS,
    Edge from TopoDS,
    Face from TopoDS,
    Vertex from TopoDS,
    ShapeEnum from TopAbs,
    HDataStructure from TopOpeBRepDS

raises

    NoMoreObject from Standard,
    NoSuchObject from Standard

is

    Create returns Explorer;

    Create(HDS:HDataStructure;T:ShapeEnum = TopAbs_SHAPE;findkeep : Boolean = Standard_True) returns Explorer;
    
    Init(me:in out;HDS:HDataStructure;T:ShapeEnum = TopAbs_SHAPE;findkeep : Boolean = Standard_True);

    Type(me) returns ShapeEnum from TopAbs;

    More(me) returns Boolean;

    Next(me : in out) raises NoMoreObject; -- when More returned False

    Current(me) returns Shape raises NoSuchObject from Standard; -- when More returns False;
    ---C++: return const &

    Index(me) returns Integer raises NoSuchObject from Standard; -- when More returns False;

    Face(me) returns Face raises NoSuchObject from Standard; -- when More returns False;
    ---C++: return const &

    Edge(me) returns Edge raises NoSuchObject from Standard; -- when More returns False;
    ---C++: return const &

    Vertex(me) returns Vertex raises NoSuchObject from Standard; -- when More returns False;
    ---C++: return const &        


    Find(me:in out) is private;
    
fields

    myHDS : HDataStructure from TopOpeBRepDS;
    myT : ShapeEnum from TopAbs;
    myI,myN : Integer;
    myB : Boolean;
    myFK : Boolean;

end Explorer from TopOpeBRepDS;
