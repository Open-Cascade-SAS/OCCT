-- Created on: 1992-11-18
-- Created by: Christian CAILLET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SelectType  from IFSelect   inherits SelectAnyType

    ---Purpose : A SelectType keeps or rejects Entities of which the Type
    --           is Kind of a given Cdl Type

uses Type, AsciiString from TCollection, Transient

is

    Create returns SelectType;
    ---Purpose : Creates a SelectType. Default is no filter

    Create (atype : Type) returns SelectType;
    ---Purpose : Creates a SelectType for a given Type

    SetType (me : mutable; atype : Type);
    ---Purpose : Sets a TYpe for filter

    TypeForMatch (me) returns Type;
    ---Purpose : Returns the Type to be matched for select : this is the type
    --           given at instantiation time

    ExtractLabel (me) returns AsciiString from TCollection;
    ---Purpose : Returns a text defining the criterium.
    --           (should by gotten from Type of Entity used for instantiation)

fields

    thetype : Type;

end SelectType;
