-- File:	StepRepr_CompoundRepresentationItem.cdl
-- Created:	Tue Apr 24 17:51:25 2001
-- Author:	Christian CAILLET
--		<cky@photox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 2001

class CompoundRepresentationItem  from StepRepr
  inherits RepresentationItem  from StepRepr

    ---Purpose : Added for Dimensional Tolerances

uses
    HAsciiString from TCollection,
    HArray1OfRepresentationItem from StepRepr

is

    Create returns CompoundRepresentationItem;

    Init (me : mutable;
             aName : mutable HAsciiString from TCollection;
	     item_element : HArray1OfRepresentationItem from StepRepr);

    ItemElement (me) returns HArray1OfRepresentationItem from StepRepr;
    NbItemElement (me) returns Integer;
    SetItemElement (me : mutable; item_element : HArray1OfRepresentationItem from StepRepr);
    ItemElementValue (me; num : Integer) returns RepresentationItem;
    SetItemElementValue (me : mutable; num : Integer;
    	anelement : RepresentationItem);

fields

    theItemElement : HArray1OfRepresentationItem from StepRepr;

end CompoundRepresentationItem;
