-- File:        AutoDesignPresentedItem.cdl
-- Created:     Mon Dec  4 12:02:23 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWAutoDesignPresentedItem from RWStepAP214

	---Purpose : Read & Write Module for AutoDesignPresentedItem

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     AutoDesignPresentedItem from StepAP214,
     EntityIterator from Interface

is

	Create returns RWAutoDesignPresentedItem;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable AutoDesignPresentedItem from StepAP214);

	WriteStep (me; SW : in out StepWriter; ent : AutoDesignPresentedItem from StepAP214);

	Share(me; ent : AutoDesignPresentedItem from StepAP214; iter : in out EntityIterator);

end RWAutoDesignPresentedItem;
