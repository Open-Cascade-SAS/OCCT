-- Created on: 1999-04-01
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Marker from TopOpeBRepDS inherits TShared from MMgt    	
uses
    HArray1OfBoolean from TColStd,
    AsciiString from TCollection
is
    Create returns mutable Marker;
    Reset(me:mutable);
    Set(me:mutable;i:Integer;b:Boolean);
    Set(me:mutable;b:Boolean;n:Integer;a:Address);
    GetI(me;i:Integer) returns Boolean;
    Allocate(me:mutable;n:Integer);    
fields
    myhe : HArray1OfBoolean from TColStd;
    myne : Integer;   
end Marker from TopOpeBRepDS;
