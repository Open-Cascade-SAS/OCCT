-- Created on: 1996-11-14
-- Created by: Philippe MANGIN
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class PrefAndRec from AdvApprox inherits Cutting from AdvApprox

    ---Purpose : 
    -- inherits class Cutting; contains a list of preferential points (pi)i
    -- and a list of Recommended points used in cutting management.
    

uses Array1OfReal from TColStd

raises DomainError from Standard
    
is
    Create(RecomendedCut : Array1OfReal;
           PrefferedCut  : Array1OfReal;
           Weight        : Real = 5 ) 
    returns PrefAndRec 
    raises DomainError;  -- if  Weight <= 1
    
    Value(me; a,b : Real;
              cuttingvalue : out Real)
    returns Boolean 
    ---Purpose: 
    --     cuting value is
    --    - the recommended point nerest of (a+b)/2 
    --      if pi is in ]a,b[ or else
    --   -  the preferential point nearest of (a+b) / 2
    --     if pi is in ](r*a+b)/(r+1) , (a+r*b)/(r+1)[ where r = Weight
    --   -  or (a+b)/2 else.
    is redefined;


fields
    myRecCutting : Array1OfReal from TColStd;
    myPrefCutting: Array1OfReal from TColStd;
    myWeight     : Real;
end PrefAndRec;
