-- Created on: 2002-04-10
-- Created by: QA Admin
-- Copyright (c) 2002-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class  MyText  from  QABugs  inherits  InteractiveObject  from  AIS 
uses 
    ExtendedString from TCollection, 
    Pnt from gp, 
    PresentationManager3d from PrsMgr, 
    Presentation from Prs3d,
    NameOfColor  from  Quantity,
    Selection from SelectMgr
is 
    Create(aText  :ExtendedString  from  TCollection;aPosition  : Pnt  from  gp)
    returns mutable MyText from QABugs;
    Create(aText  :ExtendedString  from  TCollection;aPosition  : Pnt  from  gp;aFont :  CString from Standard; aColor : NameOfColor  from  Quantity; aHeight :Real  from  Standard)
    returns mutable MyText from QABugs;

    NbPossibleSelection(me)
    returns Integer from Standard
    is redefined virtual protected;
    
    Compute(me:mutable;
            aPresentationManager: PresentationManager3d from PrsMgr;
            aPresentation: mutable Presentation from Prs3d;
            aMode: Integer from Standard = 0)
    is redefined virtual protected;

    ComputeSelection(me:mutable; aSelection :mutable Selection from SelectMgr;
                                 aMode      : Integer) is redefined virtual protected;

fields
        myPosition                   : Pnt from gp;
        myText                       : ExtendedString from TCollection;
        myNameOfColor                : NameOfColor from Quantity;
        myNameOfFont                 : CString from Standard;
        myHeight                     : Real from Standard;
end MyText;
    
