-- Created on: 1994-04-05
-- Created by: Yves FRICAUD
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



private class FunctionInter from Bisector  
inherits FunctionWithDerivative from math 

        ---Purpose:                           2                      2 
	--          F(u) =  (PC(u) - PBis1(u))   + (PC(u) - PBis2(u))

uses 
    Curve   from Geom2d,
    Curve   from Bisector
	--          

is

    Create  returns FunctionInter from Bisector;
    
    Create (C     : Curve   from Geom2d ;
            Bis1  : Curve   from Bisector;
	    Bis2  : Curve   from Bisector)  
    returns FunctionInter from Bisector;
    
    Perform (me    : in out;
    	     C     : Curve   from Geom2d ;
             Bis1  : Curve   from Bisector;
	     Bis2  : Curve   from Bisector)
    is static;	     	
	     
    Value(me : in out; X : Real; F : out Real) 
    	---Purpose: Computes the values of the Functions for the variable <X>.
    returns Boolean
    is static;
    
    Derivative(me : in out; X : Real; D : out Real) 
    returns Boolean;

    Values(me : in out ; X  : Real; F  : out Real; D  : out Real)    
    	---Purpose: Returns the values of the functions and the derivatives
    	--          for the variable <X>.
    returns Boolean
    is static;
    
fields
    
    curve     : Curve from Geom2d;
    bisector1 : Curve from Bisector;
    bisector2 : Curve from Bisector;
    
end FunctionInter;
