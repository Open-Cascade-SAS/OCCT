-- Created on: 1998-07-24
-- Created by: Christian CAILLET
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MaterialDesignation  from StepRepr

inherits TShared  from MMgt

uses

	HAsciiString from TCollection, 
	CharacterizedDefinition from StepRepr

is

    Create returns mutable MaterialDesignation;

    Init (me : mutable;
    	  aName : mutable HAsciiString from TCollection;
	  aOfDefinition : CharacterizedDefinition);


	-- Specific Methods for Field Data Access --

	SetName(me : mutable; aName : mutable HAsciiString);
	Name (me) returns mutable HAsciiString;
    	SetOfDefinition (me : mutable; aOfDefinition : CharacterizedDefinition);
	OfDefinition (me) returns CharacterizedDefinition;

fields

    	name : HAsciiString from TCollection;
    	ofDefinition : CharacterizedDefinition;

end MaterialDesignation;
