-- Created on: 2000-09-07
-- Created by: TURIN  Anatoliy <ati@nnov.matra-dtv.fr>
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DocumentStorageDriver from StdDrivers inherits DocumentStorageDriver from MDocStd

	---Purpose: storage driver of a  Part document


uses Document from CDM, 
     MessageDriver from CDM,
     Document     from PCDM,
     SequenceOfDocument from PCDM,
     ExtendedString from  TCollection,
     ASDriverTable from MDF


is

    Create
    returns DocumentStorageDriver from StdDrivers;
    
    Make(me : mutable; aDocument :     Document from CDM;
                       Documents : out SequenceOfDocument from PCDM)
    is redefined; 
    
    AttributeDrivers(me : mutable;  theMessageDriver : MessageDriver from CDM)
    returns ASDriverTable from MDF
    is redefined;
    
end DocumentStorageDriver;
