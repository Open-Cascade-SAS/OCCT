-- Created on: 2001-01-04
-- Copyright (c) 2001-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ArrayOfPoints from Graphic3d inherits ArrayOfPrimitives from Graphic3d

is

  -- constructor
  Create (maxVertexs: Integer from Standard;
          hasVColors: Boolean from Standard = Standard_False)
  returns ArrayOfPoints from Graphic3d;
  ---Purpose: Creates an array of points,
  -- a single pixel point is drawn at each vertex.
  -- The array must be filled using the AddVertex(Point) method. 
  -- When <hasVColors> is TRUE , you must use only AddVertex(Point,Color) method.

end;
