-- Created on: 1994-03-22
-- Created by: Frederic UNTEREINER
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package IGESToBRep

    ---Purpose : Provides tools in order to transfer IGES entities
    --         to CAS.CADE.

uses

    Interface,
    Transfer,
    MoniTool,
    Message,
    IGESData,
    IGESBasic,
    IGESGeom,
    IGESSolid,
    gp,
    Geom,
    Geom2d,
    TColGeom,
    TColGeom2d,
    TColStd,
    TopoDS,
    TopTools,
    ShapeExtend,
    ShapeAnalysis
    
is

    class CurveAndSurface;
    	class BasicSurface;
    	class BasicCurve;
    	class TopoSurface;
    	class TopoCurve;
    	class BRepEntity;

    class IGESBoundary;
    class Reader;
    class Actor;
    class AlgoContainer;
    class ToolContainer;
 
    Init;                                                                                                                
        ---Purpose: Creates and initializes default AlgoContainer.     
 
    SetAlgoContainer (aContainer: AlgoContainer from IGESToBRep);                                                          
        ---Purpose: Sets default AlgoContainer                                                                           
                                                                                                                         
    AlgoContainer returns AlgoContainer from IGESToBRep;                                                                   
        ---Purpose: Returns default AlgoContainer    
	
    IsCurveAndSurface(start : IGESEntity from IGESData)
    	returns Boolean;
        ---Purpose: Return True if the IGESEntity can be transfered by
    	--          TransferCurveAndSurface.
    	--          ex: All IGESEntity from IGESGeom


    IsBasicCurve  (start : IGESEntity from IGESData)
    	returns Boolean;
    	---Purpose: Return True if the IGESEntity can be transfered by
    	--          TransferBasicCurve.
    	--          ex: CircularArc, ConicArc, Line, CopiousData,
    	--              BSplineCurve, SplineCurve... from IGESGeom :
    	--              104,110,112,126


    IsBasicSurface(start : IGESEntity from IGESData)
    	returns Boolean;
      	---Purpose: Return True if the IGESEntity can be transfered by
    	--          TransferBasicSurface.
    	--          ex: BSplineSurface, SplineSurface... from IGESGeom :
    	--              114,128
     

    IsTopoCurve(start : IGESEntity from IGESData)
    	returns Boolean;
      	---Purpose: Return True if the IGESEntity can be transfered by
    	--          TransferTopoCurve.         
    	--          ex: all Curves from IGESGeom :
    	--              all basic curves,102,130,142,144

     
    IsTopoSurface(start : IGESEntity from IGESData)
    	returns Boolean;
     	---Purpose: Return True if the IGESEntity can be transfered by
    	--          TransferTopoSurface.
    	--          ex: All Surfaces from IGESGeom : 
    	--              all basic surfaces,108,118,120,122,141,143
     

    IsBRepEntity  (start : IGESEntity from IGESData)
    	returns Boolean;
    	---Purpose: Return True if the IGESEntity can be transfered by
    	--          TransferBRepEntity.
    	--          ex: VertexList, EdgeList, Loop, Face, Shell, 
    	--              Manifold Solid BRep Object from IGESSolid :
    	--              502, 504, 508, 510, 514, 186.

    WriteShape(shape  : Shape from TopoDS;
    	       number : Integer from Standard);
    	---Purpose: Creates  a file  Shape_'number' with the shape being
    	--          able to be restored by Draw.

    IGESCurveToSequenceOfIGESCurve (curve   : IGESEntity from IGESData;
    	    	    	    	    sequence: out HSequenceOfTransient from TColStd)
    returns Integer;
    
    TransferPCurve (fromedge: Edge from TopoDS;
    	    	    toedge  : Edge from TopoDS;
    	    	    face    : Face from TopoDS)
    returns Boolean;
    
end IGESToBRep;


