-- Created on: 1994-05-26
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Transition from TopOpeBRepDS 

uses

    State from TopAbs,
    Orientation from TopAbs,
    ShapeEnum from TopAbs,
    OStream from Standard

is

    Create returns Transition from TopOpeBRepDS;

    Create(StateBefore,StateAfter : State from TopAbs;
    	   ShapeBefore : ShapeEnum from TopAbs = TopAbs_FACE;
    	   ShapeAfter  : ShapeEnum from TopAbs = TopAbs_FACE) 
    returns Transition from TopOpeBRepDS;

    Create(O : Orientation from TopAbs)
    returns Transition from TopOpeBRepDS;

    Set(me : in out; 
    	StateBefore, StateAfter : State from TopAbs;
	ShapeBefore : ShapeEnum from TopAbs = TopAbs_FACE;
    	ShapeAfter  : ShapeEnum from TopAbs = TopAbs_FACE);

    StateBefore(me : in out; S : State from TopAbs);
    StateAfter(me : in out; S : State from TopAbs);
    ShapeBefore(me : in out; SE : ShapeEnum from TopAbs);
    ShapeAfter(me : in out; SE : ShapeEnum from TopAbs);
    Before(me : in out; S : State from TopAbs;ShapeBefore : ShapeEnum from TopAbs = TopAbs_FACE);
    After(me : in out; S : State from TopAbs;ShapeAfter : ShapeEnum from TopAbs = TopAbs_FACE);

    Index(me : in out; I : Integer);
    IndexBefore(me : in out; I : Integer);
    IndexAfter(me : in out; I : Integer);

    Before(me) returns State from TopAbs;
    ONBefore(me) returns ShapeEnum from TopAbs;
    After(me) returns State from TopAbs;
    ONAfter(me) returns ShapeEnum from TopAbs;
    ShapeBefore(me) returns ShapeEnum from TopAbs;
    ShapeAfter(me) returns ShapeEnum from TopAbs;
    Index(me) returns Integer; -- index of ShapeBefore (may be null)
    IndexBefore(me) returns Integer; -- index of ShapeBefore (may be null)
    IndexAfter(me) returns Integer;  -- index of ShapeAfter (may be null)

    Set(me : in out; O : Orientation from TopAbs);
    ---Purpose: set the transition corresponding to orientation <O>
    --
    --       O       Before  After
    --       
    --   FORWARD       OUT    IN 
    --   REVERSED      IN     OUT
    --   INTERNAL      IN     IN
    --   EXTERNAL      OUT    OUT
    -- 

    Orientation(me; S : State from TopAbs;
    	    	    T : ShapeEnum from TopAbs = TopAbs_FACE) 

    ---Purpose: returns the orientation corresponding to state <S> 
    -- 
    -- Before and After not equal TopAbs_ON :
    -- --------------------------------------                   
    -- Before  After   Computed orientation
    -- 
    --  S      not S   REVERSED (we leave state S)
    --  not S  S       FORWARD  (we enter state S)
    --  S      S       INTERNAL (we stay in state S)
    --  not S  not S   EXTERNAL (we stay outside state S)
    returns Orientation from TopAbs;

    OrientationON(me; S : State from TopAbs;
    	    	      T : ShapeEnum from TopAbs) 

    ---Purpose: returns the orientation corresponding to state <S> 
    --          (if one at least of the internal states is ON)
    returns Orientation from TopAbs
    is static private;

    Complement(me) returns Transition from TopOpeBRepDS;

    IsUnknown(me) returns Boolean from Standard;
    ---Purpose: returns True if both states are UNKNOWN
    
    DumpA(me; OS : in out OStream from Standard) returns OStream; 
    ---C++: return &

    DumpB(me; OS : in out OStream from Standard) returns OStream;
    ---C++: return &

    Dump(me; OS : in out OStream from Standard) returns OStream;    
    ---C++: return &
        
fields

    myStateBefore, myStateAfter : State from TopAbs;
    myShapeBefore, myShapeAfter : ShapeEnum from TopAbs;
    myIndexBefore, myIndexAfter : Integer from Standard;
    
end Transition from TopOpeBRepDS;
