-- Created by: Peter KURNEV
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Tools from BOPAlgo 

---Purpose: 

uses  
    BaseAllocator from BOPCol, 
    IndexedDataMapOfIntegerListOfInteger from BOPCol,  
    DataMapOfIntegerListOfInteger from BOPCol, 
    PDS from BOPDS, 
    PaveBlock from BOPDS,  
    IndexedDataMapOfPaveBlockListOfInteger from BOPDS, 
    IndexedDataMapOfPaveBlockListOfPaveBlock from BOPDS, 
    DataMapOfIntegerListOfPaveBlock from BOPDS
--raises

is
    --- 
    --- static methods 
    --- 
    MakeBlocksCnx(myclass; 
        theMILI     :IndexedDataMapOfIntegerListOfInteger from BOPCol; 
        theMBlocks  :out DataMapOfIntegerListOfInteger from BOPCol; 
        theAllocator:out BaseAllocator from BOPCol);  

    MakeBlocks(myclass; 
        theMILI     :IndexedDataMapOfPaveBlockListOfPaveBlock from BOPDS; 
        theMBlocks  :out DataMapOfIntegerListOfPaveBlock from BOPDS; 
        theAllocator:out BaseAllocator from BOPCol); 
 
    PerformCommonBlocks(myclass; 
        theMBlocks  :out IndexedDataMapOfPaveBlockListOfPaveBlock from BOPDS; 
        theAllocator:out BaseAllocator from BOPCol; 
        pDS: out PDS from BOPDS);
    
    FillMap(myclass; 
        tneN1:Integer from Standard; 
        tneN2:Integer from Standard; 
        theMILI : out IndexedDataMapOfIntegerListOfInteger from BOPCol; 
        theAllocator: out BaseAllocator from BOPCol); 
    
     
    FillMap(myclass; 
        tnePB1:PaveBlock from BOPDS; 
        tnePB2:PaveBlock from BOPDS; 
        theMILI : out IndexedDataMapOfPaveBlockListOfPaveBlock from BOPDS; 
        theAllocator: out BaseAllocator from BOPCol);
 
    FillMap(myclass; 
        tnePB1:PaveBlock from BOPDS; 
        tneF:Integer from Standard;  
        theMILI : out IndexedDataMapOfPaveBlockListOfInteger from BOPDS; 
        theAllocator: out BaseAllocator from BOPCol); 
 
    PerformCommonBlocks(myclass; 
        theMBlocks  :IndexedDataMapOfPaveBlockListOfInteger from BOPDS; 
        theAllocator:out BaseAllocator from BOPCol; 
        pDS: out PDS from BOPDS);
--fields

end Tools;
