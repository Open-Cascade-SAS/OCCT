-- Created on: 2003-05-06
-- Created by: Michael KLOKOV
-- Copyright (c) 2003-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Tools from QANewModTopOpe
uses
    Edge from TopoDS,
    Shape from TopoDS,
    State from TopAbs,
    PPaveFiller from BOPAlgo, 
    PBOP from BOPAlgo,
    ListOfShape from TopTools,
    IndexedDataMapOfShapeListOfShape from TopTools

is

    NbPoints(myclass; theDSFiller: PPaveFiller from BOPAlgo)
    	returns Integer from Standard;

    NewVertex(myclass; theDSFiller: PPaveFiller from BOPAlgo;
    	    	       theIndex   : Integer from Standard)
    	returns Shape from TopoDS;

    HasSameDomain(myclass; theBuilder: PBOP from BOPAlgo;
    	    	    	   theFace    : Shape from TopoDS)
    	returns Boolean from Standard;
    
    SameDomain(myclass; theBuilder: PBOP from BOPAlgo;
    	    	    	theFace    : Shape from TopoDS;
    	    	    	theResultList: out ListOfShape from TopTools);

    IsSplit(myclass; theDSFiller: PPaveFiller from BOPAlgo;
    	    	     theEdge    : Shape from TopoDS;
    	    	     theState   : State from TopAbs)
    	returns Boolean from Standard;
	---Warning: This method could be called only after boolean operation,
	---         arguments of which was solids or compounds of solids.
	---

    Splits(myclass; theDSFiller: PPaveFiller from BOPAlgo;
    	    	    theEdge    : Shape from TopoDS;
    	    	    theState   : State from TopAbs;
    	    	    theResultList: out ListOfShape from TopTools);
	---Warning: This method could be called only after boolean operation,
	---         arguments of which was solids or compounds of solids.
	---

    SplitE(myclass; theEdge  : Edge from TopoDS;
    	    	    theSplits: out ListOfShape from TopTools)
    	returns Boolean from Standard;

    EdgeCurveAncestors(myclass; theDSFiller: PPaveFiller from BOPAlgo;
    	    	    	    	theEdge    : Shape from TopoDS;
				theFace1   : out Shape from TopoDS;
				theFace2   : out Shape from TopoDS)
    	returns Boolean from Standard;
    
    EdgeSectionAncestors(myclass; theDSFiller: PPaveFiller from BOPAlgo;
    	    	    	    	  theEdge    : Shape from TopoDS;
    	    	    	    	  LF1,LF2    : out ListOfShape from TopTools;
				  LE1,LE2 : out ListOfShape from TopTools)
    	returns Boolean from Standard;

    BoolOpe(myclass; theFace1: Shape from TopoDS;
    	    	     theFace2: Shape from TopoDS;
		     IsCommonFound: out Boolean from Standard;
    	    	     theHistoryMap: out IndexedDataMapOfShapeListOfShape from TopTools)
    	returns Boolean from Standard;

end Tools from QANewModTopOpe;
