-- Created on: 1998-06-03
-- Created by: data exchange team
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package ShapeAnalysis 

    ---Purpose: This package is intended to analyze geometrical objects
-- and topological shapes. Analysis domain includes both
-- exploring geometrical and topological properties of
-- shapes and checking their conformance to Open CASCADE requirements.
-- The directions of analysis provided by tools of this package are:
-- computing quantities of subshapes,  
-- computing parameters of points on curve and surface,  
-- computing surface singularities,  
-- checking edge and wire consistency,  
-- checking edges order in the wire,  
-- checking face bounds orientation,  
-- checking small faces,  
-- analyzing shape tolerances,  
-- analyzing of free bounds of the shape.  

uses
    gp,
    TColStd,
    TCollection,
    TColgp,
    Bnd,
    Geom, 
    Geom2d,
    GeomAdaptor,
    Extrema,
    IntRes2d,
    TopAbs,
    TopLoc,
    TopoDS,
    TopTools,
    ShapeExtend,
    Adaptor3d
    
is
 
    class Geom;

    class Curve;

    class Surface;

    class Edge;

    class Wire;

    class WireOrder;

    class WireVertex;

    class CheckSmallFace;                                                                                 

    class Shell;		    

    class ShapeTolerance;

    --class OverlapEdges;  now it is in package OverlapShape of Products
    --- Container for keeping information about
	--          overlapping edges

    --class CheckCoincidenceTool;  now it is in package OverlapShape of Products
    ---Tool for checking coincidence of faces and edges

     -- Class intended for analyzing shape contents
    
    class ShapeContents;

    -- Classes intended for free bounds analysis

    class FreeBounds;

    class FreeBoundData;

    class FreeBoundsProperties;

    class TransferParameters;

	class TransferParametersProj;

    imported SequenceOfFreeBounds;

    imported transient class HSequenceOfFreeBounds;

    imported DataMapOfShapeListOfReal;

    imported DataMapIteratorOfDataMapOfShapeListOfReal;

    --class SequenceOfOverlapEdges instantiates 
    	--Sequence from TCollection (OverlapEdges from ShapeAnalysis); 
	    -- now it is in package OverlapShape of Products
	
    --class IndexedDataMapOfShapeSequenceOfOverlapEdges instantiates
    	--IndexedDataMap from TCollection(Shape          from TopoDS,
	    	    	    	    	--SequenceOfOverlapEdges from ShapeAnalysis,
                                        --ShapeMapHasher from TopTools);
	    -- now it is in package OverlapShape of Products
					

    OuterWire (face: Face from TopoDS) returns Wire from TopoDS;
        ---Purpose: Returns the outer wire on the face <Face>.
	--          This is replacement of the method BRepTools::OuterWire
	--          until it works badly.
	--          Returns the first wire oriented as outer according to
	--          FClass2d_Classifier. If none, last wire is returned.

    TotCross2D(sewd: WireData from ShapeExtend; aFace: Face from TopoDS)
    returns Real;
    	---Purpose: Returns a total area of 2d wire
	
    ContourArea(theWire : Wire from TopoDS) returns Real;
       --sewd: WireData from ShapeExtend) returns Real;
    	---Purpose: Returns a total area of 3d wire
	
    IsOuterBound (face: Face from TopoDS) returns Boolean;
    	---Purpose: Returns True if <F> has outer bound.
	---Remarks: This method checks only presence of outer bound, it does not
	--          check mutual orientation of the bounds on a face

    AdjustByPeriod(Val: Real; ToVal: Real; Period: Real)
    returns Real;
    	---Purpose: Returns a shift required to move point
        --          <Val> to the range [ToVal-Period/2,ToVal+Period/2].
        --          This shift will be the divisible by Period.
	--          Intended for adjusting parameters on periodic surfaces.
	
    AdjustToPeriod(Val: Real; ValMin: Real; ValMax: Real)
    returns Real;
    	---Purpose: Returns a shift required to move point
        --          <Val> to the range [ValMin,ValMax].
        --          This shift will be the divisible by Period
        --          with Period = ValMax - ValMin.
	--          Intended for adjusting parameters on periodic surfaces.

    FindBounds (shape: Shape  from TopoDS;
		V1   : in out Vertex from TopoDS;
		V2   : in out Vertex from TopoDS);
    	---Purpose: Finds the start and end vertices of the shape
	--          Shape can be of the following type:
	--          vertex: V1 and V2 are the same and equal to <shape>,
	--          edge  : V1 is start and V2 is end vertex (see ShapeAnalysis_Edge
    	--                  methods FirstVertex and LastVertex),
	--          wire  : V1 is start vertex of the first edge, V2 is end vertex
	--                  of the last edge (also see ShapeAnalysis_Edge).
	--                  If wire contains no edges V1 and V2 are nullified
	--          If none of the above V1 and V2 are nullified
	---Remark:  V1 and V2 can be of any orientation
	
    GetFaceUVBounds(F: Face from TopoDS; Umin, Umax, Vmin, Vmax: out Real);
    	---Purpose: Computes exact UV bounds of all wires on the face        
	
end ShapeAnalysis;
