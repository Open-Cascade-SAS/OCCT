-- Created on: 1995-10-24
-- Created by: Mister rmi
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



package PPoly 

	---Purpose: This  package  provides  persistent classes  to
	--          handle :
	--          
	--          * 3D triangular polyhedrons.
	--          
	--          * 3D polygons.
	--          
	--          * 2D polygon.

uses    PCollection,
        PColStd,
   	PColgp

is

    class Triangle;
	---Purpose: A triangle is  a triplet  of integers (indices  of
	--          the nodes).
    
    class Triangulation;
	---Purpose: A   Triangulation  is  a   3D  polyhedron made  of
	--          triangles.  It   is  made  of  a nodes  which  are
	--          indexed. Nodes  have a 3d  value  and a  2d value.
	--          Triangles are triplet of node indices.
	--          
	--          This is a Transient class.


    class Polygon3D;
    	---Purpose: A Polygon3D is  made of  indexed nodes.
    	--          Nodes have a 3d value.

    class Polygon2D;
    	---Purpose: A Polygon2D is made of  indexed nodes.
    	--          Nodes have a 2d value.
	  
    class PolygonOnTriangulation;
    	---Purpose: A polygonOnTriangulation is made of node indices
    	--          referencing a triangulation.

    class HArray1OfTriangle
    instantiates HArray1 from PCollection(Triangle from PPoly);

end PPoly;
