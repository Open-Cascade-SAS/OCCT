-- Created on: 1993-06-24
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class GeomTool from TopOpeBRep 

    ---Purpose: Provide services needed by the DSFiller

uses

    Curve from Geom,
    Curve from Geom2d,
    Face from TopoDS,
    Shape from TopoDS,
    Curve from TopOpeBRepDS,
    LineInter from TopOpeBRep 
    
is

    Create returns GeomTool from TopOpeBRep;
    
    MakeCurves(myclass;
     	       min,max:Real;L:LineInter from TopOpeBRep;
    	       S1,S2:Shape from TopoDS;
     	       C:out Curve from TopOpeBRepDS;
    	       PC1,PC2:out Curve from Geom2d);
    ---Purpose: Make the  DS curve <C> and the pcurves <PC1,PC2> from
    -- intersection line <L> lying on shapes <S1,S2>. <min,max> = <L> bounds

    MakeCurve(myclass;
     	      min,max:Real;L:LineInter from TopOpeBRep;
     	      C : out Curve from Geom);

    MakePrivateCurves
    (myclass;  
     min,max:Real;L:LineInter from TopOpeBRep;S1,S2:Shape from TopoDS;
     C:out Curve from Geom;
     PC1,PC2:out Curve from Geom2d;
     New:out Boolean;
     tolreached2d1,tolreached2d2:out Real);

    MakeBSpline1fromWALKING3d  
    (myclass; L:LineInter from TopOpeBRep) returns Curve from Geom;
 
    MakeBSpline1fromWALKING2d 
    (myclass;L:LineInter from TopOpeBRep;SI:Integer) returns Curve from Geom2d;
 
end GeomTool from TopOpeBRep;
