-- Created on: 1993-01-09
-- Created by: CKY / Contract Toubro-Larsen ( SIVA )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class ToroidalSurface from IGESSolid  inherits IGESEntity

        ---Purpose: defines ToroidalSurface, Type <198> Form Number <0,1>
        --          in package IGESSolid
        --          This entity is defined by the center point, the axis
        --          direction and the major and minor radii. In case of
        --          parametrised surface a reference direction is provided.

uses

        Point           from IGESGeom,
        Direction       from IGESGeom,
        Pnt             from gp

is

        Create returns mutable ToroidalSurface;

        -- Specific Methods pertaining to the class

        Init (me        : mutable;
              aCenter   : Point;
              anAxis    : Direction;
              majRadius : Real;
              minRadius : Real;
              Refdir    : Direction);
        ---Purpose : This method is used to set the fields of the class
        --           ToroidalSurface
        --       - aCenter   : the center point coordinates
        --       - anAxis    : the direction of the axis
        --       - majRadius : the major radius
        --       - minRadius : the minor radius
        --       - Refdir    : the reference direction (parametrised)
        --                     default Null for unparametrised surface

        Center(me) returns Point;
        ---Purpose : returns the center point coordinates of the surface

        TransformedCenter(me) returns Pnt;
        ---Purpose : returns the center point coordinates of the surface
        -- after applying TransformationMatrix

        Axis(me) returns Direction;
        ---Purpose : returns the direction of the axis

        MajorRadius(me) returns Real;
        ---Purpose : returns the major radius of the surface

        MinorRadius(me) returns Real;
        ---Purpose : returns the minor radius of the surface

        ReferenceDir(me) returns Direction;
        ---Purpose : returns the reference direction (parametrised surface)
        -- Null is returned if the surface is not parametrised

        IsParametrised(me) returns Boolean;
        ---Purpose : Returns True if the surface is parametrised, else False

fields

--
-- Class    : IGESSolid_ToroidalSurface
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class ToroidalSurface.
--
-- Reminder : A ToroidalSurface instance is defined by :
--            This entity is defined by the center point, the axis
--            direction and the major and minor radii. In case of
--            parametrised surface a reference direction is provided.
--

        theCenter      : Point;
            -- the center point coordinates of the surface

        theAxis        : Direction;
            -- the direction of the axis

        theMajorRadius : Real;
            -- the major radius of the surface

        theMinorRadius : Real;
            -- the minor radius of the surface

        theRefDir      : Direction;
            -- the reference direction of the surface (parametrised)

end ToroidalSurface;
