-- Created on: 1992-07-21
-- Created by: Laurent PAINNOT
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

generic class CurveLocator from Extrema 
    (Curve1 as any;
     Tool1  as any;   -- as ToolCurve(Curve1)
     Curve2 as any;
     Tool2  as any;   -- as ToolCurve(Curve2)
     POnC   as any;
     Pnt    as any)
					
     
is

    Locate (myclass; P: Pnt; C: Curve1; NbU: Integer; Papp: out POnC);
    ---Purpose: Among a set of points {C(ui),i=1,NbU}, locate the point
    --          P=C(uj) such that:
    --           distance(P,C) = Min{distance(P,C(ui))}


    Locate (myclass; P: Pnt; C: Curve1; NbU: Integer; Umin, Usup: Real;Papp: out POnC);
    ---Purpose: Among a set of points {C(ui),i=1,NbU}, locate the point
    --          P=C(uj) such that:
    --           distance(P,C) = Min{distance(P,C(ui))}
    --           The research is done between umin and usup.


   Locate (myclass; C1: Curve1; C2: Curve2; NbU, NbV: Integer; Papp1, Papp2: out POnC);
    ---Purpose: Among two sets of points {C1(ui),i=1,NbU} and
    --          {C2(vj),j=1,NbV}, locate the two points P1=C1(uk) and 
    --          P2=C2(vl) such that:
    --           distance(P1,P2) = Min {distance(C1(ui),C2(vj))}.


end CurveLocator;
