-- Created on: 2000-08-16
-- Created by: data exchange team
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Color from PXCAFDoc  inherits Attribute from PDF

	---Purpose: 

uses
    Color from Quantity

is
    Create returns mutable Color from PXCAFDoc;
    
    Create (Loc: Color from Quantity) returns mutable Color from PXCAFDoc;
    
    Set (me: mutable; Loc: Color from Quantity);
    
    Get (me) returns Color from Quantity;
    
fields
    myColor : Color from Quantity;
    
end Color;
