-- Created on: 1993-09-29
-- Created by: Denis PASCAL
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class RGNode from GraphTools

uses SC                from GraphTools,
     SequenceOfInteger from TColStd

is

    Create returns RGNode;
    
    Reset (me : in out);
    
    SetVisited (me : in out; v : Integer from Standard);
    
    GetVisited (me) 
    returns Integer from Standard;
    
    AddAdj (me : in out; adj : Integer from Standard);
    
    NbAdj (me) 
    returns Integer from Standard;
    
    GetAdj (me; index : Integer from Standard)
    returns Integer from Standard;

    SetSC (me : in out; SC : SC from GraphTools);

    GetSC (me) 
    returns SC from GraphTools;

fields

    visited : Integer from Standard;
    myAdj   : SequenceOfInteger from TColStd;
    mySC    : SC from GraphTools;

end RGNode;      	

