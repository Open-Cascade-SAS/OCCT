-- Created on: 2003-01-22
-- Created by: data exchange team
-- Copyright (c) 2003-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class FeaCurveSectionGeometricRelationship from StepFEA
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity FeaCurveSectionGeometricRelationship

uses
    CurveElementSectionDefinition from StepElement,
    AnalysisItemWithinRepresentation from StepElement

is
    Create returns FeaCurveSectionGeometricRelationship from StepFEA;
	---Purpose: Empty constructor

    Init (me: mutable; aSectionRef: CurveElementSectionDefinition from StepElement;
                       aItem: AnalysisItemWithinRepresentation from StepElement);
	---Purpose: Initialize all fields (own and inherited)

    SectionRef (me) returns CurveElementSectionDefinition from StepElement;
	---Purpose: Returns field SectionRef
    SetSectionRef (me: mutable; SectionRef: CurveElementSectionDefinition from StepElement);
	---Purpose: Set field SectionRef

    Item (me) returns AnalysisItemWithinRepresentation from StepElement;
	---Purpose: Returns field Item
    SetItem (me: mutable; Item: AnalysisItemWithinRepresentation from StepElement);
	---Purpose: Set field Item

fields
    theSectionRef: CurveElementSectionDefinition from StepElement;
    theItem: AnalysisItemWithinRepresentation from StepElement;

end FeaCurveSectionGeometricRelationship;
