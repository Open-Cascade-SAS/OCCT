-- Created on: 1999-09-20
-- Created by: Peter KURNEV
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class ShapeWithState from TopOpeBRepDS 

	---Purpose: 

uses
    Shape from TopoDS, 
    ListOfShape  from  TopTools,
    State from TopAbs 


is
    Create returns  ShapeWithState from TopOpeBRepDS ;
     
    Part  (me;  aState: State from TopAbs)  returns ListOfShape  from  TopTools ;  
    ---C++:  return  const& 
     
    AddPart (me:out;  aShape:Shape  from  TopoDS;  aState: State from TopAbs);  

    AddParts (me:out; aListOfShape:ListOfShape  from  TopTools;  aState: State from TopAbs);  
     
    SetState  (me:out;  aState: State from TopAbs);  
    
    State  (me)  returns  State from TopAbs; 
     
    SetIsSplitted  (me:out;  anIsSplitted:Boolean  from  Standard); 
     
    IsSplitted  (me)  returns  Boolean  from  Standard; 
    
fields
  
    myPartIn   :  ListOfShape  from  TopTools; 
    myPartOut  :  ListOfShape  from  TopTools; 
    myPartOn   :  ListOfShape  from  TopTools; 
    myState:  State from TopAbs ; 
    myIsSplitted:  Boolean  from  Standard; 
     
end ShapeWithState;
