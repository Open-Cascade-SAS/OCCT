-- Created on: 1993-07-13
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Curve2d from BRepAdaptor inherits Curve from Geom2dAdaptor

	---Purpose: The Curve2d from BRepAdaptor allows to use an Edge
	--          on   a Face like   a  2d   curve. (curve  in   the
	--          parametric space).
	--          
	--          It  has  the methods    of the class Curve2d  from
	--          Adpator. 
	--          
	--          It  is created or  initialized with a  Face and an
	--          Edge.  The methods are  inherited from  Curve from
	--          Geom2dAdaptor. 

uses
    Face from TopoDS,
    Edge from TopoDS

raises
    NullObject from Standard

is

    Create returns Curve2d from BRepAdaptor;
	---Purpose: Creates an uninitialized curve2d.

    Create(E : Edge from TopoDS; F : Face from TopoDS)
    returns Curve2d from BRepAdaptor
	---Purpose: Creates with the pcurve of <E> on <F>.
    raises
    	NullObject from Standard; -- if <E> has no pcurve on <F>
	
    Initialize(me : in out; E : Edge from TopoDS; F : Face from TopoDS)
	---Purpose: Initialize with the pcurve of <E> on <F>.
    raises
    	NullObject from Standard -- if <E> has no pcurve on <F>
    is static;
    
    Edge(me) returns Edge from TopoDS
	---Purpose: Returns the Edge.
	--          
	---C++: return const &
    is static;

    Face(me) returns Face from TopoDS
	---Purpose: Returns the Face.
	--          
	---C++: return const &
    is static;

fields

    myEdge : Edge from TopoDS;
    myFace : Face from TopoDS;
	
end Curve2d;
