-- Created on: 2008-03-27
-- Created by: Sergey ZARITCHNY
-- Copyright (c) 2008-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ExtStringArray_1 from PDataStd inherits Attribute from PDF

	---Purpose: Persistence

uses  HExtendedString          from PCollection,
      HArray1OfExtendedString  from PColStd
     
     
is

    Create returns mutable ExtStringArray_1 from PDataStd;

    Init(me : mutable; lower, upper : Integer from Standard);

    SetValue(me: mutable; Index : Integer from Standard; Value : HExtendedString from PCollection);
    
    Value(me;  Index : Integer from Standard) returns HExtendedString from PCollection;
   
    Lower (me) returns Integer from Standard;      

    Upper (me) returns Integer from Standard;   
     
    SetDelta(me : mutable; delta : Boolean from Standard); 
     
    GetDelta(me) returns Boolean from Standard;
     
fields
    myValue     :  HArray1OfExtendedString from PColStd;
    myDelta  : Boolean from Standard;

end ExtStringArray_1;



