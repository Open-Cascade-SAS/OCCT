-- Created on: 1995-02-16
-- Created by: Dieter THIEMANN
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class FacetedTool from TopoDSToStep

    ---Purpose: This Tool Class provides Information about Faceted Shapes
    --          to be mapped to STEP.

uses

    Shape  from TopoDS,
    FacetedError from TopoDSToStep

is    
    
--  -----------------------------------------------------------
--  just class methods
--  -----------------------------------------------------------


    CheckTopoDSShape(myclass; SH : Shape from TopoDS)
		     returns FacetedError from TopoDSToStep;


end FacetedTool from TopoDSToStep;

