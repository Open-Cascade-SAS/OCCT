-- Created on: 1997-02-10
-- Created by: Odile Olivier
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class XYZPlanePresentation from DsgPrs
    	---Purpose: A framework for displaying the planes of an XYZ trihedron.
uses

    Presentation from Prs3d,
    Drawer       from Prs3d,
    Pnt          from gp

is

    Add(myclass;
    	aPresentation: Presentation from Prs3d;
    	aDrawer      : Drawer from Prs3d;
    	aPt1         : Pnt    from gp;
    	aPt2         : Pnt    from gp;
    	aPt3         : Pnt    from gp);
	 
    	---Purpose: Draws each plane of a trihedron displayed in the
    	-- presentation aPresentation and with attributes
    	-- defined by the attribute manager aDrawer. Each
    	-- triangular plane is defined by the points aPt1 aPt2 and aPt3.

end XYZPlanePresentation;
