-- Created on: 1997-03-05
-- Created by: Joelle CHAUVET
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PlateG0Criterion from GeomPlate inherits Criterion from AdvApp2Var


uses
    SequenceOfXY,SequenceOfXYZ from TColgp,
    Patch,Context from AdvApp2Var,
    CriterionType,CriterionRepartition from AdvApp2Var


is

    Create( Data : SequenceOfXY;
    	    G0Data : SequenceOfXYZ;
            Maximum : Real;
    	    Type : CriterionType  = AdvApp2Var_Absolute;
    	    Repart : CriterionRepartition  = AdvApp2Var_Regular)  returns PlateG0Criterion;
	    
    Value(me; P : in out Patch; C : Context )
    is redefined;
    
    IsSatisfied(me; P : Patch ) returns Boolean
    is redefined;
    

    
fields
    myData : SequenceOfXY;
    myXYZ : SequenceOfXYZ;
    
end PlateG0Criterion;

