-- Created on: 1992-06-22
-- Created by: Gilles DEBARBOUILLE
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class UnitsDictionary from Units 

inherits

        TShared from MMgt 
	---Purpose: This class creates  a dictionary of all  the units
	--          you want to know.

uses

    HAsciiString       from TCollection,
    AsciiString        from TCollection,
    Quantity           from Units,
    QuantitiesSequence from Units,
    Dimensions         from Units


is

    Create returns mutable UnitsDictionary from Units;
    
    ---Level: Internal 
    
    ---Purpose: Returns an empty instance of UnitsDictionary.
    
    Creates(me : mutable ; afilename : CString)
    
    ---Level: Internal 
    
    ---Purpose: Returns a  UnitsDictionary object  which  contains the
    --          sequence  of all   the  units  you want to   consider,
    --          physical quantity by physical quantity.
    
    is static;
    
    Sequence(me) returns any QuantitiesSequence from Units
    
    ---Level: Internal 
    
    ---C++: inline
    
    ---Purpose: Returns   the  head   of   the  sequence  of  physical
    --          quantities.
    
    is static;
    
    UpToDate(me) returns Boolean
    
    ---Level: Internal 
    
    ---Purpose: Returns true if there has been no  modification of the
    --          file Units.dat  since the   creation of the dictionary
    --          object, false otherwise.
    
    is static;
    
    ActiveUnit(me ; aquantity : CString) returns AsciiString from TCollection
    
    ---Level: Internal 
    
    ---Purpose: Returns for <aquantity> the active unit.

    is static;
    
    Dump(me ; alevel : Integer)
    
    ---Level: Internal 
    
    ---C++: inline
    
    ---Purpose: Dumps only  the sequence   of  quantities without  the
    --          units  if  <alevel> is  equal  to zero,  and  for each
    --          quantity all the units stored if <alevel>  is equal to
    --          one.
    
    is static;

    Dump(me ; adimensions : Dimensions)
    
    ---Level: Internal 
    
    ---C++: inline
    
    ---Purpose: Dumps  for a     designated  physical       dimensions
    --          <adimensions> all the previously stored units.
    
    is static;

fields

    thefilename           : HAsciiString from TCollection;
    thetime               : Integer;
    thequantitiessequence : QuantitiesSequence from Units;

end UnitsDictionary;











