-- Created on: 2001-04-24
-- Created by: Christian CAILLET
-- Copyright (c) 2001-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MeasureRepresentationItemAndQualifiedRepresentationItem  from StepShape
    inherits RepresentationItem  from StepRepr

    ---Purpose : Added for Dimensional Tolerances
    --           Complex Type between MeasureRepresentationItem and
    --             QualifiedRepresentationItem

uses
    HArray1OfValueQualifier from StepShape,
    ValueQualifier from StepShape,
    HAsciiString from TCollection,
    Unit               from StepBasic,
    MeasureWithUnit    from StepBasic,
    MeasureValueMember from StepBasic
 
is

    Create returns MeasureRepresentationItemAndQualifiedRepresentationItem;

    Init (me : mutable;
          aName : HAsciiString from TCollection;
          aValueComponent : MeasureValueMember from StepBasic;
          aUnitComponent : Unit from StepBasic;
    	  qualifiers : HArray1OfValueQualifier from StepShape);

    	--  About MeasureReprItem

    SetMeasure (me: mutable; Measure: MeasureWithUnit from StepBasic);
    Measure (me) returns MeasureWithUnit from StepBasic;

    	--  About QualifiedReprItem

    Qualifiers (me) returns HArray1OfValueQualifier from StepShape;
    NbQualifiers (me) returns Integer;
    SetQualifiers (me : mutable; qualifiers : HArray1OfValueQualifier from StepShape);
    QualifiersValue (me; num : Integer) returns ValueQualifier from StepShape;
    SetQualifiersValue (me : mutable; num : Integer; aqualifier : ValueQualifier from StepShape);

fields

    myMeasure: MeasureWithUnit from StepBasic;
    theQualifiers : HArray1OfValueQualifier from StepShape;

end MeasureRepresentationItemAndQualifiedRepresentationItem;
