-- Created on: 1995-12-07
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.





class GeneralModule from RWStepAP214  inherits GeneralModule from StepData
	---Purpose : Defines General Services for StepAP214 Entities
	--           (Share,Check,Copy; Trace already inherited)
	--           Depends (for case numbers) of Protocol from StepAP214

uses Transient,  HAsciiString from TCollection,
     EntityIterator from Interface,
     ShareTool      from Interface,
     Check          from Interface,
     CopyTool       from Interface,
     InterfaceModel from Interface

is

    Create returns mutable GeneralModule from RWStepAP214;
    ---Purpose : Creates a GeneralModule

    FillSharedCase (me; CN : Integer; ent : Transient;
                        iter : in out EntityIterator);
    ---Purpose : Specific filling of the list of Entities shared by an Entity
    --           <ent>, according to a Case Number <CN> (provided by StepAP214
    --           Protocol).

    CheckCase (me; CN : Integer; ent : Transient; shares : ShareTool; ach : in out Check);
    ---Purpose : Specific Checking of an Entity <ent>

    CopyCase (me; CN : Integer; entfrom : Transient; entto : mutable Transient; TC : in out CopyTool);
    ---Purpose : Specific Copy ("Deep") from <entfrom> to <entto> (same type)
    --           by using a CopyTool which provides its working Map.
    --           Use method Transferred from CopyTool to work


    NewVoid (me; CN : Integer; ent : out mutable Transient) returns Boolean;

    CategoryNumber (me; CN : Integer; ent : Transient; shares : ShareTool)
    returns Integer  is redefined;

    Name (me; CN : Integer; ent : Transient; shares : ShareTool from Interface)
    returns HAsciiString from TCollection  is redefined;
    ---Purpose : Returns the name of a STEP Entity according to its type

end GeneralModule;
