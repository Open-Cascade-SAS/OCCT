-- Created on: 1997-03-28
-- Created by: Philippe MANGIN
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



private class SearchSing from ChFi3d inherits FunctionWithDerivative from math

	---Purpose: F(t) = (C1(t) - C2(t)).(C1'(t) - C2'(t));

uses Curve from Geom

is
    Create(C1, C2 : Curve from Geom)
    returns SearchSing from ChFi3d;

    Value(me: in out; X: Real; F: out Real)
    	---Purpose: computes the value of the function <F> for the 
    	--          variable <X>. 
    	--          returns True if the computation was done successfully,
    	--          False otherwise.
    returns Boolean;
    
    Derivative(me: in out; X: Real; D: out Real)
         ---Purpose: computes the derivative <D> of the function 
         --          for the variable <X>.
    	--           Returns True if the calculation were successfully done, 
    	--           False otherwise.

    returns Boolean;    

    Values(me: in out; X: Real; F, D: out Real)
    	---Purpose: computes the value <F> and the derivative <D> of the 
    	--          function for the variable <X>.
    	--          Returns True if the calculation were successfully done,
    	--          False otherwise.

    returns Boolean;

fields
myC1 : Curve from Geom;
myC2 : Curve from Geom;
end SearchSing;
