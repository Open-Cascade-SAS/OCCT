-- Created on: 2012-02-10
-- Created by: Serey ZERCHANINOV
-- Copyright (c) 2012-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class Polygon2d from Intf

	---Purpose: 

uses Pnt2d from gp,
     Box2d from Bnd

raises OutOfRange from Standard

is

    Bounding (me)
        returns Box2d from Bnd;
    ---C++: return const &
    ---C++: inline
    ---Purpose: Returns the bounding box of the polygon.

    Closed (me)
        returns Boolean from Standard is virtual;
    ---Purpose: Returns True if the polyline is closed.

    DeflectionOverEstimation (me) returns Real from Standard is deferred;
    ---Purpose: Returns the tolerance of the polygon.

    NbSegments (me) returns Integer from Standard is deferred;
    ---Purpose: Returns the number of Segments in the polyline.

    Segment (me; theIndex : in Integer from Standard;
                 theBegin, theEnd : in out Pnt2d from gp)
        raises OutOfRange from Standard is deferred;
    ---Purpose: Returns the points of the segment <Index> in the Polygon.

fields

    myBox   : Box2d from Bnd is protected;

end Polygon2d;
