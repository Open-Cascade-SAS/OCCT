-- Created on: 1998-06-30
-- Created by: Christian CAILLET
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class AssemblyComponentUsageSubstitute  from StepRepr    inherits TShared from MMgt

uses
     HAsciiString from TCollection,
     AssemblyComponentUsage from StepRepr

is

    Create returns mutable AssemblyComponentUsageSubstitute;

    Init (me : mutable;
    	  aName : HAsciiString;
	  aDef  : HAsciiString;
	  aBase : AssemblyComponentUsage;
	  aSubs : AssemblyComponentUsage);

    Name (me) returns HAsciiString;
    SetName (me : mutable; aName : HAsciiString);

    Definition (me) returns HAsciiString;
    SetDefinition (me : mutable; aDef : HAsciiString);

    Base (me) returns AssemblyComponentUsage;
    SetBase (me : mutable; aBase : AssemblyComponentUsage);

    Substitute (me) returns AssemblyComponentUsage;
    SetSubstitute (me : mutable; aSubstitute : AssemblyComponentUsage);

fields

    theName : HAsciiString;
    theDef  : HAsciiString;
    theBase : AssemblyComponentUsage;
    theSubs : AssemblyComponentUsage;

end AssemblyComponentUsageSubstitute;
