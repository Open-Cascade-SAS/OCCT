-- Created on: 1998-02-02
-- Created by: Philippe MANGIN
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

private  class LocFunction from GeomFill 

	---Purpose: 

uses 
 LocationLaw from GeomFill,
 Array1OfVec   from TColgp, 
 Mat  from  gp

is 
    Create( Law  :  LocationLaw  from  GeomFill) 
    returns  LocFunction  from  GeomFill; 
     
    
   D0(me : in  out; 
      Param: Real;
      First, Last : Real)
      ---Purpose: compute the section for v = param           
   returns Boolean; 
	
   D1(me : in  out;
      Param: Real;
      First, Last : Real)
      ---Purpose: compute the first  derivative in v direction  of the
      --           section for v =  param 
   returns Boolean;
   
    D2(me : in  out;
      Param: Real;
      First, Last : Real)      
      ---Purpose: compute the second derivative  in v direction of the
      --          section  for v = param  
   returns Boolean; 
    
   DN(me  :  in  out;
      Param       : Real;
      First, Last : Real; 
      Order       :  Integer; 
      Result      :  in  out  Real; 
      Ier         :  out  Integer); 

fields 
  myLaw  :  LocationLaw  from  GeomFill;
  V,  DV,  D2V  :  Array1OfVec  from  TColgp; 
  M,  DM,  D2M  :  Mat  from  gp;
end LocFunction;
