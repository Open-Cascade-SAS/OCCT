-- Created on: 1998-04-08
-- Created by: Andre LIEUTIER
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package NLPlate

uses
     Plate, Geom, TCollection, TColStd,
     math, gp, TColgp,  GeomAbs
is

    class NLPlate;
-- Constraints Class
    deferred  class HGPPConstraint; 
    class  HPG0Constraint; 
    class  HPG0G1Constraint;
    class  HPG0G2Constraint;
    class  HPG0G3Constraint;
    class  HPG1Constraint;
    class  HPG2Constraint;
    class  HPG3Constraint;
--  

-- utilities and internal Classes
    imported StackOfPlate;
    imported ListIteratorOfStackOfPlate;   
    imported SequenceOfHGPPConstraint;   
end NLPlate;
