-- Created on: 1997-01-03
-- Created by: Christian CAILLET
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class PDescr  from StepData    inherits TShared

    ---Purpose : This class is intended to describe the authorized form for a
    --           parameter, as a type or a value for a field
    --           
    --           A PDescr firstly describes a type, which can be SELECT, i.e.
    --           have several members

uses CString, Type from Standard, AsciiString from TCollection,
     Check from Interface,
     EnumTool from StepData, Field from StepData, EDescr from StepData

is

    Create returns PDescr;

    SetName (me : mutable; name : CString);
    Name    (me) returns CString;

    	--  basic settings

    Kind (me) returns Integer  is private;

    SetSelect (me : mutable);
    ---Purpose : Declares this PDescr to be a Select, hence to have members
    --           <me> itself can be the first member

    AddMember (me : mutable; member : PDescr);
    ---Purpose : Adds a member to a SELECT description

    SetMemberName (me : mutable; memname : CString);
    ---Purpose : Sets a name for SELECT member. To be used if a member is for
    --           an immediate type

    SetInteger (me : mutable);
    ---Purpose : Sets <me> for an Integer value

    SetReal    (me : mutable);
    ---Purpose : Sets <me> for a Real value

    SetString  (me : mutable);
    ---Purpose : Sets <me> for a String value

    SetBoolean (me : mutable);
    ---Purpose : Sets <me> for a Boolean value (false,true)

    SetLogical (me : mutable);
    ---Purpose : Sets <me> for a Logical value (false,true,unknown)

    SetEnum    (me : mutable);
    ---Purpose : Sets <me> for an Enum value
    --           Then, call AddEnumDef ordered from the first one (value 0)

    AddEnumDef (me : mutable; enumdef : CString);
    ---Purpose : Adds an enum value as a string

    SetType    (me : mutable; atype : Type from Standard);
    ---Purpose : Sets <me> for an Entity which must match a Type (early-bound)

    SetDescr   (me : mutable; dscnam : CString);
    ---Purpose : Sets <me> for a Described Entity, whose Description must match
    --           the type name  <dscnam>

    AddArity   (me : mutable; arity : Integer = 1);
    ---Purpose : Adds an arity count to <me>, by default 1
    --           1 : a simple field passes to a LIST/ARRAY etc
    --               or a LIST to a LIST OF LIST
    --           2 : a simple field passes to a LIST OF LIST

    SetArity   (me : mutable; arity : Integer = 1);
    ---Purpose : Directly sets the arity count
    --           0 : simple field
    --           1 : LIST or ARRAY etc
    --           2 : LIST OF LIST

    	-- complements

    SetFrom (me : mutable; other : PDescr);
    ---Purpose : Sets <me> as <other> but duplicated
    --           Hence, some definition may be changed

    SetOptional (me : mutable; opt : Boolean = Standard_True);
    ---Purpose : Sets/Unsets <me> to accept undefined values

    SetDerived  (me : mutable; der : Boolean = Standard_True);
    ---Purpose : Sets/Unsets <me> to be for a derived field

    SetField    (me : mutable; name : CString; rank : Integer);
    ---Purpose : Sets <me> to describe a field of an entity
    --           With a name and a rank

    	-- querying

    IsSelect  (me) returns Boolean;
    ---Purpose : Tells if <me> is for a SELECT

    Member    (me; name : CString) returns PDescr;
    ---Purpose : For a SELECT, returns the member whose name matches <name>
    --           To this member, the following question can then be asked
    --           Null Handle if <name> not matched or <me> not a SELECT
    --           
    --           Remark : not to be asked for an entity type
    --           Hence, following IsInteger .. Enum* only apply on <me> and
    --           require Member
    --           While IsType applies on <me> and all Select Members

    IsInteger (me) returns Boolean;
    ---Purpose : Tells if <me> is for an Integer

    IsReal    (me) returns Boolean;
    ---Purpose : Tells if <me> is for a Real value

    IsString  (me) returns Boolean;
    ---Purpose : Tells if <me> is for a String value

    IsBoolean (me) returns Boolean;
    ---Purpose : Tells if <me> is for a Boolean value (false,true)

    IsLogical (me) returns Boolean;
    ---Purpose : Tells if <me> is for a Logical value (false,true,unknown)

    IsEnum    (me) returns Boolean;
    ---Purpose : Tells if <me> is for an Enum value
    --           Then, call AddEnumDef ordered from the first one (value 0)
    --           Managed by an EnumTool

    EnumMax   (me) returns Integer;
    ---Purpose : Returns the maximum integer for a suitable value (count - 1)

    EnumValue (me; name : CString) returns Integer;
    ---Purpose : Returns the numeric value found for an enum text
    --           The text must be in capitals and limited by dots
    --           A non-suitable text gives a negative value to be returned
 
    EnumText  (me; val  : Integer) returns CString;
    ---Purpose : Returns the text which corresponds to a numeric value,
    --           between 0 and EnumMax. It is limited by dots

    IsEntity  (me) returns Boolean;
    ---Purpose : Tells if <me> is for an Entity, either Described or CDL Type

    IsType    (me; atype : Type from Standard) returns Boolean;
    ---Purpose : Tells if <me> is for an entity of a given CDL type (early-bnd)
    --           (works for <me> + nexts if <me> is a Select)

    Type      (me) returns Type from Standard;
    ---Purpose : Returns the type to match (IsKind), for a CDL Entity
    --           (else, null handle)

    IsDescr   (me; descr : EDescr from StepData) returns Boolean;
    ---Purpose : Tells if <me> is for a Described entity of a given EDescr
    --           (does this EDescr match description name ?). For late-bnd
    --           (works for <me> + nexts if <me> is a Select)

    DescrName (me) returns CString;
    ---Purpose : Returns the description (type name) to match, for a Described
    --           (else, empty string)

    Arity (me) returns Integer;
    ---Purpose : Returns the arity of <me>

    Simple (me) returns PDescr;
    ---Purpose : For a LIST or LIST OF LIST, Returns the PDescr for the simpler
    --           PDescr. Else, returns <me>
    --           This allows to have different attributes for Optional for
    --           instance, on a field, and on the parameter of a LIST :
    --           [OPTIONAL] LIST OF [OPTIONAL] ...

    IsOptional (me) returns Boolean;
    ---Purpose : Tells if <me> is Optional

    IsDerived  (me) returns Boolean;
    ---Purpose : Tells if <me> is Derived

    IsField    (me) returns Boolean;
    ---Purpose : Tells if <me> is a Field. Else it is a Type

    FieldName  (me) returns CString;
    FieldRank  (me) returns Integer;

    Check (me; afild : Field; ach : in out Check)  is virtual;
    ---Purpose : Semantic Check of a Field : does it complies with the given
    --           description ?

fields

    thename : AsciiString from TCollection;
    thesel  : Integer;  -- 0 no  1 entity  2 immediate  3 heterog. 4 unknown
    thesnam : AsciiString from TCollection;
    thenext : PDescr;   -- list of members
    thekind : Integer;  -- as Field
    theenum : EnumTool from StepData;
    thetype : Type from Standard;
    thednam : AsciiString from TCollection;
    thearit : Integer;
    thefrom : PDescr;   -- for SetFrom
    theopt  : Boolean;
    theder  : Boolean;
    thefnam : AsciiString from TCollection;
    thefnum : Integer;

end PDescr;
