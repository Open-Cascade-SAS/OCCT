-- Created on: 2002-12-10
-- Created by: data exchange team
-- Copyright (c) 2002-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V2.0

class SurfaceElementPurpose from StepElement
inherits SelectType from StepData

    ---Purpose: Representation of STEP SELECT type SurfaceElementPurpose

uses
    SelectMember from StepData,
    EnumeratedSurfaceElementPurpose from StepElement,
    HAsciiString from TCollection

is
    Create returns SurfaceElementPurpose from StepElement;
	---Purpose: Empty constructor

    CaseNum (me; ent: Transient) returns Integer;
	---Purpose: Recognizes a kind of SurfaceElementPurpose select type
	--          return 0 

    CaseMem (me; ent: SelectMember from StepData) returns Integer is redefined;
	---Purpose: Recognizes a items of select member SurfaceElementPurposeMember
	--          1 -> EnumeratedSurfaceElementPurpose
	--          2 -> ApplicationDefinedElementPurpose
	--          0 else


     NewMember(me) returns SelectMember from StepData is redefined;
	---Purpose: Returns a new select member the type SurfaceElementPurposeMember

    SetEnumeratedSurfaceElementPurpose(me: in out; aVal :EnumeratedSurfaceElementPurpose from StepElement);
	---Purpose: Set Value for EnumeratedSurfaceElementPurpose

    EnumeratedSurfaceElementPurpose (me) returns EnumeratedSurfaceElementPurpose from StepElement;
	---Purpose: Returns Value as EnumeratedSurfaceElementPurpose (or Null if another type)

    SetApplicationDefinedElementPurpose(me: in out; aVal :HAsciiString from TCollection);
	---Purpose: Set Value for ApplicationDefinedElementPurpose

    ApplicationDefinedElementPurpose (me) returns HAsciiString from TCollection;
	---Purpose: Returns Value as ApplicationDefinedElementPurpose (or Null if another type)

end SurfaceElementPurpose;
