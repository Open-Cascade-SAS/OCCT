-- File:        BoxDomain.cdl
-- Created:     Mon Dec  4 12:02:24 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWBoxDomain from RWStepShape

	---Purpose : Read & Write Module for BoxDomain

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     BoxDomain from StepShape,
     EntityIterator from Interface

is

	Create returns RWBoxDomain;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable BoxDomain from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : BoxDomain from StepShape);

	Share(me; ent : BoxDomain from StepShape; iter : in out EntityIterator);

end RWBoxDomain;
