-- File:        CompositeText.cdl
-- Created:     Mon Dec  4 12:02:24 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWCompositeText from RWStepVisual

	---Purpose : Read & Write Module for CompositeText

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     CompositeText from StepVisual,
     EntityIterator from Interface

is

	Create returns RWCompositeText;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable CompositeText from StepVisual);

	WriteStep (me; SW : in out StepWriter; ent : CompositeText from StepVisual);

	Share(me; ent : CompositeText from StepVisual; iter : in out EntityIterator);

end RWCompositeText;
