-- Created on: 1993-03-03
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Update:      fma


class Datum3D from PTopLoc inherits Persistent from Standard

	---Purpose: An  elementary local coordinate system. It  may be
	--          shared in the Database.

uses
    Trsf from gp

raises
    ConstructionError from Standard

is
    Create(T : Trsf from gp) returns mutable Datum3D from PTopLoc
	---Purpose: Creates a   local coordinate  system    with   the
	--          transformation.  An   error   is raised  if    the
	--          transformation is not rigid.
	---Level: Internal 
    raises
    	ConstructionError from Standard;
	
    Transformation(me) returns Trsf from gp
    	---Purpose: Returns the transformation defining the coordinate
    	--          system.
	---Level: Internal 
    is static;
    
fields

    myTrsf : Trsf from gp;

end Datum3D;
