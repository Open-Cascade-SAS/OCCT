-- File:	Blend_AppFunction.cdl
-- Created:	Mon Sep 13 16:54:05 1993
-- Author:	Jacques GOUSSARD
--		<jag@topsn2>
---Copyright:	 Matra Datavision 1993


deferred class AppFunction from Blend

inherits FunctionSetWithDerivatives from math

    ---Purpose: Deferred class for a function used to compute a blending
    --          surface between two surfaces, using a guide line.
    --          The vector <X> used in Value, Values and Derivatives methods
    --          has to be the vector of the parametric coordinates U1,V1,
    --          U2,V2, of the extremities of a section on the first and
    --          second surface.

uses Vector from math,
     Matrix from math,
     Pnt    from gp,
     Shape  from GeomAbs,
     Point  from Blend,
     Array1OfPnt     from TColgp,
     Array1OfVec     from TColgp,
     Array1OfPnt2d   from TColgp,
     Array1OfVec2d   from TColgp,
     Array1OfReal    from TColStd,
     Array1OfInteger from TColStd



raises DomainError from Standard

is

	
    NbVariables(me)
	---Purpose: returns the number of variables of the function.
    	returns Integer from Standard
	is deferred;

    NbEquations(me)
    	---Purpose: returns the number of equations of the function.
    	returns Integer from Standard
	is deferred;

    Value(me: in out; X: Vector; F: out Vector)
    	---Purpose: computes the values <F> of the Functions for the 
    	--          variable <X>.
    	--          Returns True if the computation was done successfully, 
    	--          False otherwise.

    	returns Boolean from Standard
	is deferred;
    
    
    Derivatives(me: in out; X: Vector; D: out Matrix)
    	---Purpose: returns the values <D> of the derivatives for the 
    	--          variable <X>.
    	--          Returns True if the computation was done successfully, 
    	--          False otherwise.

    returns Boolean from Standard
    is deferred;
    
    
    Values(me: in out; X: Vector; F: out Vector; D: out Matrix)
    	---Purpose: returns the values <F> of the functions and the derivatives
    	--          <D> for the variable <X>.
    	--          Returns True if the computation was done successfully, 
    	--          False otherwise.

    returns Boolean from Standard
    is deferred;
    
 
    Set(me: in out; Param: Real from Standard)
    
	---Purpose: Sets the value of the parameter along the guide line.
	--          This determines the plane in which the solution has
	--          to be found.

    	is deferred;
	
    Set(me: in out; First, Last: Real from Standard)
    
	---Purpose: Sets the bounds of the parametric interval on 
	--          the guide line.
	--          This determines the derivatives in these values if the
	--          function is not Cn.
    	is deferred;    


    GetTolerance(me; Tolerance: out Vector from math; Tol: Real from Standard)
    
	---Purpose: Returns in the vector Tolerance the parametric tolerance
	--          for each of the 4 variables;
	--          Tol is the tolerance used in 3d space.
    
    	is deferred;


    GetBounds(me; InfBound,SupBound: out Vector from math)
    
	---Purpose: Returns in the vector InfBound the lowest values allowed
	--          for each of the 4 variables.
	--          Returns in the vector SupBound the greatest values allowed
	--          for each of the 4 variables.
    
    	is deferred;


   IsSolution(me: in out; Sol: Vector from math; Tol: Real from Standard)
    	---Purpose: Returns Standard_True if Sol is a zero of the function.
	--          Tol is the tolerance used in 3d space.
	--          The computation is made at the current value of
	--          the parameter on the guide line.
    
    	returns Boolean from Standard
    	is deferred; 
	 
   GetMinimalDistance(me) 
        ---Purpose: Returns   the    minimal  Distance  beetween   two
        --          extremitys of calculed sections.          
   	returns  Real  from  Standard 
	is  deferred; 
	 
   Pnt1(me)
       	---Purpose: Returns the point on the first support.
	---C++: return const &
    	returns Pnt from gp 
    	is deferred;

   Pnt2(me)   
       	---Purpose: Returns the point on the first support.
	---C++: return const &     	
    	returns Pnt from gp 
    	is deferred;

-- Methods for the approximation
-- 
    IsRational(me) returns Boolean
	---Purpose: Returns  if the section is rationnal
    is deferred;
    
    GetSectionSize(me) returns Real
    	---Purpose:  Returns the length of the maximum section
    is deferred;
    
    GetMinimalWeight(me; Weigths  : out Array1OfReal  from TColStd)
    	---Purpose: Compute the minimal value of weight for each poles
    	--          of all sections.
    is deferred;

    NbIntervals(me; S : Shape from GeomAbs) returns Integer
	---Purpose: Returns  the number  of  intervals for  continuity
	--          <S>. May be one if Continuity(me) >= <S>
    is deferred;
    
    Intervals(me; T : in out Array1OfReal from TColStd; 
    	          S : Shape from GeomAbs)
	---Purpose: Stores in <T> the  parameters bounding the intervals
	--          of continuity <S>.
	--          
	--          The array must provide  enough room to  accomodate
	--          for the parameters. i.e. T.Length() > NbIntervals()
--    raises
--    	OutOfRange from Standard 
    is deferred;

    GetShape(me: in out;
                 NbPoles   : out Integer from Standard;
                 NbKnots   : out Integer from Standard;
                 Degree    : out Integer from Standard;
                 NbPoles2d : out Integer from Standard)

    	is deferred;

    GetTolerance(me; 
    	    	 BoundTol, SurfTol, AngleTol : Real;
		 Tol3d : out Vector;
		 Tol1D : out Vector )
	---Purpose: Returns the tolerance to reach in approximation
	--          to respecte
	--          BoundTol error at the Boundary
	--          AngleTol tangent error at the Boundary
	--          SurfTol error inside the surface.
        is deferred;

    Knots(me: in out; TKnots: out Array1OfReal from TColStd)

	is deferred;


    Mults(me: in out; TMults: out Array1OfInteger from TColStd)

	is deferred;


    Section(me: in out; P: Point from Blend;
			Poles    : out Array1OfPnt   from TColgp;
			DPoles   : out Array1OfVec   from TColgp;
    	                Poles2d  : out Array1OfPnt2d from TColgp;
			DPoles2d : out Array1OfVec2d from TColgp;
			Weigths  : out Array1OfReal  from TColStd;
			DWeigths : out Array1OfReal  from TColStd)

	---Purpose: Used for the first and last section 
	--          The method returns Standard_True if the derivatives
	--          are computed, otherwise it returns Standard_False.

    	returns Boolean from Standard

    	is deferred;


    Section(me: in out; P: Point from Blend;
                        Poles    : out Array1OfPnt   from TColgp;
    	                Poles2d  : out Array1OfPnt2d from TColgp;
			Weigths  : out Array1OfReal  from TColStd)
    	is deferred;
	
    Section(me: in out; P: Point from Blend;
			Poles     : out Array1OfPnt   from TColgp;
			DPoles    : out Array1OfVec   from TColgp;
			D2Poles   : out Array1OfVec   from TColgp;
    	                Poles2d   : out Array1OfPnt2d from TColgp;
			DPoles2d  : out Array1OfVec2d from TColgp;
			D2Poles2d : out Array1OfVec2d from TColgp;
			Weigths   : out Array1OfReal  from TColStd;
			DWeigths  : out Array1OfReal  from TColStd;
                        D2Weigths : out Array1OfReal  from TColStd)

	---Purpose: Used for the first and last section 
	--          The method returns Standard_True if the derivatives
	--          are computed, otherwise it returns Standard_False.

    	returns Boolean from Standard

    	is deferred;

    	Resolution(me; 
    	    	   IC2d : Integer from Standard;
		   Tol  : Real from Standard;
		   TolU, TolV : out Real from Standard)
	is deferred;

-- Static function for approx
    Parameter(me; P: Point from Blend)
	---Purpose: Returns  the parameter  of  the point  P. Used  to
	--          impose the parameters in the approximation.
    	returns Real from Standard
	is static;


end AppFunction;
