-- Created on: 1993-03-23
-- Created by: BBL,JLF
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class XWUD from ImageUtility

	---Version: 0.0

	---Purpose: Performs a "xwud -noclick" with a XAlienImage build
	-- 		 from any Image , any AlienImage .

	---Keywords:
	---Warning:
	---References:

uses
	AlienUserImage 	from AlienImage,
	XAlienImage  	from AlienImage,
	File  		from OSD,
	Image 		from Image

raises
	TypeMismatch 	from Standard

is
	XWUD( myclass ; aImage          : in Image from Image; 
			aName           : CString from Standard;
			xwudOptions     : CString from Standard 
						= "-new -noclick" ) ;
	---Level: Internal
	  ---Purpose: Write content of a Image object to aTmpFile and
	  --          execute a Spawn "xwud xwudOptions -in aTmpFile &" .

	XWUD( myclass ; aAlienUserImage : in AlienUserImage from AlienImage; 
			aName           : CString from Standard ;
			xwudOptions     : CString from Standard 
						= "-new -noclick" ) ;
	---Level: Internal
	  ---Purpose: Write content of a  AlienImage object to aTmpFile and
	  --          execute a Spawn "xwud xwudOptions -in aTmpFile &" .

	XWUD( myclass ; aXAlienImage    : in XAlienImage from AlienImage ;
			xwudOptions     : CString from Standard 
						= "-new -noclick" ) ;
	---Level: Internal
	  ---Purpose: Write content of a  XAlienImage object to aTmpFile and
	  --          execute a Spawn "xwud xwudOptions -in aTmpFile &" .

	XWUD( myclass ; aFile           : in File from OSD ;
			xwudOptions     : CString from Standard 
						= "-new -noclick" ) ;
	---Level: Internal
	  ---Purpose: execute a Spawn 
	  --	"xwud -new -noclick -in /aFile.SystemName()/ &" .

	XWUD( myclass ; aFileName       : CString from Standard ;
			xwudOptions     : CString from Standard 
						= "-new -noclick" ) ;
	---Level: Internal
	  ---Purpose: execute a Spawn "xwud xwudOptions -in aFileName &" .



end ;
