-- File:	GeomFill_FunctionDraft.cdl
-- Created:	Mon Apr 27 10:53:22 1998
-- Author:	 Stephanie HUMEAU
--		<shu@sun17>
---Copyright:	 Matra Datavision 1998

private  class FunctionDraft  from  GeomFill   
inherits  FunctionSetWithDerivatives  from  math 

uses   

    Vector from math,  
    Matrix from math, 
    HSurface  from  Adaptor3d, 
    HCurve  from  Adaptor3d, 
    Vec  from  gp, 
    Tensor  from  GeomFill

is
 
    Create(S  :  HSurface  from  Adaptor3d ;  C  :  HCurve  from  Adaptor3d)   
    returns FunctionDraft  from  GeomFill ;

    NbVariables(me)
    	---Purpose: returns the number of variables of the function.

    returns Integer  is  redefined;
    
    
    NbEquations(me)
    	---Purpose: returns the number of equations of the function.

    returns Integer  is redefined;
    
    
    Value(me: in out; X: Vector; F: out Vector)
    	---Purpose: computes the values <F> of the Functions for the 
    	--          variable <X>.
    	--          Returns True if the computation was done successfully, 
    	--          False otherwise.

    returns Boolean  is redefined;
    
    
    Derivatives(me: in out; X: Vector; D: out Matrix)
    	---Purpose: returns the values <D> of the derivatives for the 
    	--          variable <X>.
    	--          Returns True if the computation was done successfully, 
    	--          False otherwise.

    returns Boolean  is redefined;
    
    
    Values(me: in out; X: Vector; F: out Vector; D: out Matrix)
    	---Purpose: returns the values <F> of the functions and the derivatives
    	--          <D> for the variable <X>.
    	--          Returns True if the computation was done successfully, 
    	--          False otherwise.

    returns Boolean  is redefined;
   

    DerivT(me: in out;   
    	   C  :  HCurve  from  Adaptor3d; 
	   Param  :  Real  from  Standard;
	   W  :  Real  from  Standard; 
 	   dN  :  Vec  from  gp; 
    	   teta  :  Real;  
    	   F: out Vector) 
    	---Purpose: returns the values <F> of the T derivatives for
    	--          the parameter Param .
    returns Boolean  is static;
 

    Deriv2T(me: in out;  
    	    C  :  HCurve  from  Adaptor3d; 
	    Param  :  Real  from  Standard;  
       	    W  :  Real  from  Standard;  
 	    d2N  :  Vec  from  gp; 
    	    teta  :  Real;  
    	    F: out Vector)	 
    	---Purpose: returns the values <F> of the T2 derivatives for
    	--          the parameter Param .
    returns Boolean  is static;    
   
  
    DerivTX(me: in out;  
    	    dN  :  Vec  from  gp; 
    	    teta  :  Real;  
    	    D: out Matrix)	 
    	---Purpose: returns the values <D> of  the TX derivatives for
    	--          the parameter Param .
    returns Boolean  is static;        
   
      
    Deriv2X(me: in out;  
    	    X  :  Vector  from  math; 
      	    T: out Tensor)	 
	 ---Purpose: returns the values <T> of  the X2 derivatives for
    	--          the parameter Param .   
    returns Boolean  is static;     
     
     
    
fields   
    TheCurve  :  HCurve  from  Adaptor3d;
    TheSurface  :  HSurface  from  Adaptor3d;

end  FunctionDraft;
