-- Created on: 1991-07-17
-- Created by: Isabelle GRIGNON
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class FunctionSample from math 

	---Purpose: This class gives a default sample (constant difference
	--          of parameter) for a function defined between
	--          two bound A,B.

raises OutOfRange from Standard

is

    Create(A,B: Real; N: Integer)
    
    	returns FunctionSample from math;


    Bounds(me; A,B: out Real) is virtual;
    
	---Purpose: Returns the bounds of parameters.



    NbPoints(me)
    
	---Purpose: Returns the number of sample points.

    returns Integer
    is static;


    GetParameter(me; Index: Integer)
    
	---Purpose: Returns the value of parameter of the point of 
	--          range Index : A + ((Index-1)/(NbPoints-1))*B.
	--          An exception is raised if Index<=0 or Index>NbPoints.

    returns Real
    raises OutOfRange
    is virtual;



fields

    a: Real;
    b: Real;
    n: Integer;

end FunctionSample;
