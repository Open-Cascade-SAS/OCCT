-- Created by: DAUTRY Philippe
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

--      	-------

---Version:	0.0
--Version	Date		Purpose
--		0.0	Mar 13 1997	Creation


package PDF 

	---Purpose: This pakage is the persistent equivalent of
	--          TDF. It describes persistent classes used to store
	--          a TDF structure into a Database.


uses

    Standard,
    PCollection,
    PColStd

is

    class Data;
    
    
    deferred class Attribute;

    class TagSource; 

    class Reference;

    -- Instantiations ---------------------------------------------------

    class HAttributeArray1 from PDF instantiates HArray1 from PCollection
    	(Attribute from PDF);

end PDF;
