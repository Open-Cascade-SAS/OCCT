-- Created on: 1996-08-21
-- Created by: Jacques MINOT
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

--              modified 12-january-98  by  Sergey ZARITCHNY

class DiameterPresentation from DsgPrs
        
    	---Purpose: A framework for displaying diameters in shapes.  
        
        
uses
    Presentation from Prs3d,
    Pnt from gp,
    Circ from gp,
    Drawer from Prs3d,
    ArrowSide from DsgPrs,
    ExtendedString from TCollection
    	
is  
    Add( myclass; aPresentation   : Presentation   from Prs3d;
    	    	  aDrawer         : Drawer         from Prs3d;
		  aText           : ExtendedString from TCollection;
                  AttachmentPoint : Pnt            from gp;
		  aCircle         : Circ           from gp; 
	          ArrowSide: ArrowSide             from DsgPrs;
    	    	  IsDiamSymbol    : Boolean        from Standard );
	---Purpose: Draws the diameter of the circle aCircle displayed in
    	-- the presentation aPresentation and with attributes
    	-- defined by the attribute manager aDrawer. The point
    	-- AttachmentPoint defines the point of contact
    	-- between the circle and the diameter presentation.
    	-- The value of the enumeration ArrowSide controls
    	-- whether arrows will be displayed at either or both
    	-- ends of the length. The text aText labels the diameter.
		   

    Add( myclass; aPresentation   : Presentation   from Prs3d;
    	    	  aDrawer         : Drawer         from Prs3d;
		  aText           : ExtendedString from TCollection;
                  AttachmentPoint : Pnt            from gp;
		  aCircle         : Circ           from gp; 
		  uFirst          : Real           from Standard; 
		  uLast           : Real           from Standard;
	          ArrowSide       : ArrowSide      from DsgPrs; 
    	    	  IsDiamSymbol    : Boolean        from Standard);
	---Purpose: Draws the diameter of the arc anArc displayed in the
    	-- presentation aPresentation and with attributes
    	-- defined by the attribute manager aDrawer. The point
    	-- AttachmentPoint defines the point of contact
    	-- between the arc and the diameter presentation. The
    	-- value of the enumeration ArrowSide controls whether
    	-- arrows will be displayed at either or both ends of the
    	-- length. The parameters uFirst and uLast define the
    	-- first and last points of the arc. The text aText labels the diameter.

end DiameterPresentation;
