-- Created on: 1995-03-08
-- Created by: Mister rmi
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

--Modified by ROB : Add ShapeFilters.
--	      GG  : 5/10/99 BUC60576 Add Cone to TypeOfFace enum


package StdSelect 

	---Purpose: The StdSelect package provides the following services
    	-- -   the definition of selection modes for topological shapes
    	-- -   the definition of several concrete filtertandard
    	--   Selection2d.ap classes
    	-- -   2D and 3D viewer selectors.
    	--  Note that each new Interactive Object must have all
    	-- its selection modes defined.
    	--        Standard Classes is useful to build
	--          3D Selectable Objects, and to process
	--          3D Selections:
	--          
	--          - Implementation of View Selector for dynamic selection
	--            in Views from V3d.
	--          
	--          - Implementation of Tool class to decompose 3D BRep Objects
	--            into sensitive Primitives for every desired mode of selection
	--            (selection of vertex,edges,wires,faces,...)
	--            
	--          -  Implementation of dedicated Sensitives Entities:
	--             Text for 2D Views (linked to Specific 2D projectors.)
uses
    MMgt,
    Standard,
    TCollection,
    TopLoc,
    TopoDS,
    SelectMgr,
    TopAbs,
    TColStd,
    gp,
    Select3D,
    Graphic3d,Visual3d,
    Quantity,
    Prs3d,
    V3d,
    PrsMgr,
    SelectBasics,
    TopTools,
    Bnd,
    Geom, 
    TColgp

is

    enumeration TypeOfResult is TOR_SIMPLE,TOR_MULTIPLE
    end TypeOfResult;
    	---Purpose: Provides values for type of result.
    	-- These are used to specify whether the result is to
    	-- be simple or whether it may be multiple.
        
    enumeration DisplayMode is DM_Wireframe,DM_Shading,DM_HLR
    end DisplayMode;
    
--    enumeration TypeOfFace is AnyFace,Plane,Cylinder,Sphere,Torus,Revol;
    enumeration TypeOfFace is AnyFace,Plane,Cylinder,Sphere,Torus,Revol,Cone;
    	---Purpose: Provides values for different types of faces. These
    	-- values are used to filter faces in frameworks inheriting
    	-- StdSelect_FaceFilter.
    
    enumeration TypeOfEdge is AnyEdge,Line,Circle;
    	---Purpose: Provides values for different types of edges. These
    	-- values are used to filter edges in frameworks
    	-- inheriting StdSelect_EdgeFilter.
    
    enumeration SensitivityMode is SM_WINDOW, SM_VIEW;
    	---Purpose: Selection sensitivity mode. SM_WINDOW mode uses the
    	-- specified pixel tolerance to compute the sensitivity value,
    	-- SM_VIEW mode allows to define the sensitivity manually.


    class ViewerSelector3d;
    	---Purpose: Viewer Selector for a view from V3d
    	--          Accepts Only Sensitive Entities inheriting Select3D entities...
    
    
    
    class BRepSelectionTool;
    	---Purpose: gives standard selections for Shapes

    class BRepOwner;
    	---Purpose: Owner classes for BRep objects 
	--          used by BRepSelectionTool to know which entities
	--          own the sensitive primitives created.
	--          the hilight-unhilight methods are empty and
	--          must be redefined by each User...

    ---Category: Shape Filters

    class EdgeFilter;
    class FaceFilter;
    class ShapeTypeFilter;

    ---Category: Private Classes

    private class Prs;

    private class Shape;

    private class IndexedDataMapOfOwnerPrs instantiates IndexedDataMap from TCollection
    (EntityOwner from SelectBasics,Prs from StdSelect,MapTransientHasher from TColStd);

    GetProjector (aView: View from V3d) returns Projector from Select3D;
    	---Purpose: Returns the 3D projector for the view aView.
    SetDrawerForBRepOwner(aSelection: mutable Selection from SelectMgr;
			  aDrawer   : Drawer from Prs3d);
     	---Purpose: puts The same drawer in every BRepOwner Of SensitivePrimitive
     	--          Used Only for hilight Of BRepOwner...
			

end StdSelect;
