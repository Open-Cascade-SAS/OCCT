-- Created on: 1994-05-31
-- Created by: Christian CAILLET
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DispPerDrawing  from IGESSelect  inherits Dispatch

    ---Purpose : This type of dispatch defines sets of entities attached to
    --           distinct drawings. This information is taken from attached
    --           views which appear in the Directory Part. Also Drawing Frames
    --           are considered when Drawings are part of input list.
    --           
    --           Remaining data concern entities not attached to a drawing.

uses AsciiString from TCollection, EntityIterator, Graph, SubPartsIterator,
     ViewSorter

is

    Create returns DispPerDrawing;
    ---Purpose : Creates a DispPerDrawing

    Label (me) returns AsciiString from TCollection;
    ---Purpose : Returns as Label, "One File per Drawing"

    	    -- --    Evaluation    -- --

    Packets (me; G : Graph; packs : in out SubPartsIterator);
    ---Purpose : Computes the list of produced Packets. Packets are computed
    --           by a ViewSorter (SortDrawings with also frames).

    CanHaveRemainder (me) returns Boolean  is redefined;
    ---Purpose : Returns True, because of entities attached to no view.

    Remainder (me; G : Graph) returns EntityIterator  is redefined;
    ---Purpose : Returns Remainder which is a set of Entities.
    --           It is supposed to be called once Packets has been called.

fields

    thesorter : ViewSorter;

end DispPerDrawing;
