-- Created on: 1997-09-03
-- Created by: Christian CAILLET
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class RealVal  from MoniTool    inherits TShared  from MMgt

    ---Purpose : A Real through a Handle (i.e. managed as TShared)

uses Real

is

    Create (val : Real = 0.0) returns RealVal;

    Value (me) returns Real;

    CValue (me : mutable) returns Real;
    ---C++ : return &

fields

    theval : Real;

end RealVal;
