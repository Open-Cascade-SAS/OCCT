-- Created on: 1998-04-17
-- Created by: Andre LIEUTIER
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class  HPG2Constraint  from  NLPlate  inherits  HPG1Constraint from  NLPlate 
---Purpose: define a PinPoint (no G0)  G2 Constraint used to load a Non
--  Linear Plate
uses
     XY from gp,
     D1  from  Plate,
     D2  from  Plate
     
is
    Create(UV : XY; D1T : D1 from Plate; D2T : D2 from Plate) returns mutable HPG2Constraint;
    -- create a G2 Constraint
    -- 


    ActiveOrder(me)  returns  Integer 
    is   redefined; 
    --  returns the constraint active  order, i.e. the maximum between
    --  -- the initial constraint i.e 2 (for G2 Constraints)
    --  
    -- 

    G2Target(me) returns D2  from  Plate 
    ---C++: return const &
    is   redefined; 

fields
    myG2Target : D2 from Plate;
end;
