-- Created on: 1993-03-17
-- Created by: Laurent BUCHARD
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

generic class PrmPrmSvSurfaces from ApproxInt (
    ThePSurface         as any;
    ThePSurfaceTool     as any;
    TheLine             as Transient)

inherits SvSurfaces from ApproxInt

uses 
    Pnt     from gp,
    Pnt2d   from gp,
    Vec     from gp,
    Vec2d   from gp

    class TheInt2S instantiates Int2S from IntImp(
    	ThePSurface,ThePSurfaceTool);

is 
    Create(Surf1,Surf2: ThePSurface);
    
    Compute(me: in out; 
            u1,v1,u2,v2: in out Real from Standard;
	    Pt: out Pnt from gp;
	    Tg: out Vec from gp;
	    Tguv1,Tguv2: out Vec2d from gp)
	    ---Purpose: returns True if Tg,Tguv1 Tguv2 can be computed.
       returns Boolean from Standard	is static;
       
    Pnt(me: in out;
    	u1,v1,u2,v2: in Real from Standard;
    	P: out Pnt from gp) is static;
	
    Tangency(me: in out;
    	     u1,v1,u2,v2: in Real from Standard;
	     Tg: out Vec from gp)
       returns Boolean from Standard is static;
       
    TangencyOnSurf1(me: in out;
    	            u1,v1,u2,v2: in Real from Standard;
	            Tg: out Vec2d from gp)
       returns Boolean from Standard is static;
       
    TangencyOnSurf2(me: in out;
    	            u1,v1,u2,v2: in Real from Standard;
	            Tg: out Vec2d from gp)
       returns Boolean from Standard is static;   
    
fields
    MyParOnS1            : Pnt2d        from gp;
    MyParOnS2            : Pnt2d        from gp;
    MyPnt                : Pnt          from gp;
    MyTguv1              : Vec2d        from gp;
    MyTguv2              : Vec2d        from gp;
    MyTg                 : Vec          from gp;
    MyIsTangent          : Boolean      from Standard;
    MyHasBeenComputed    : Boolean      from Standard;
    
    MyParOnS1bis            : Pnt2d        from gp;
    MyParOnS2bis            : Pnt2d        from gp;
    MyPntbis                : Pnt          from gp;
    MyTguv1bis              : Vec2d        from gp;
    MyTguv2bis              : Vec2d        from gp;
    MyTgbis                 : Vec          from gp;
    MyIsTangentbis          : Boolean      from Standard;
    MyHasBeenComputedbis    : Boolean      from Standard;
    
    MyIntersectionOn2S   : TheInt2S;
 
end PrmPrmSvSurfaces;



