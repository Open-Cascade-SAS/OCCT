-- Created on: 1992-10-13
-- Created by: Ramin BARRETO
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package MMgt 

---Purpose:
--   The package MMgt provides single class TShared which is second in hierarchy
--   of inheritance from Standard_Transient, kept for historic reasons

uses Standard

is
    deferred class TShared;
    ---Purpose:
    --   Intermediate class between Standard_Transient and descendants.

end MMgt;
