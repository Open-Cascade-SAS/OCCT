-- Created on: 1992-04-07
-- Created by: Christian CAILLET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



deferred class LevelListEntity  from IGESData  inherits IGESEntity

    ---Purpose : defines required type for LevelList in directory part
    --           an effective LevelList entity must inherits it

uses Boolean, Integer

raises OutOfRange

is

    NbLevelNumbers (me) returns Integer  is deferred;
    ---Purpose : Must return the count of levels

    LevelNumber (me; num : Integer) returns Integer
        raises OutOfRange  is deferred;
    ---Purpose : returns the Level Number of <me>, indicated by <num>
    -- raises an exception if num is out of range

    HasLevelNumber (me; level : Integer) returns Boolean;
    ---Purpose : returns True if <level> is in the list

end LevelListEntity;
