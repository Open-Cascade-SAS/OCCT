-- Created on: 1999-07-22
-- Created by: data exchange team
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ClosedFaceDivide from ShapeUpgrade inherits FaceDivide from ShapeUpgrade

	---Purpose: Divides a Face with one or more seam edge to avoid closed faces.
	--          Splitting is performed by U and V direction. The number of 
        --          resulting faces can be defined by user.

uses

    Face    from TopoDS

is
    
    Create returns ClosedFaceDivide from ShapeUpgrade;
    	---Purpose: Creates empty  constructor.
    
    Create (F : Face from TopoDS)
    returns ClosedFaceDivide from ShapeUpgrade;
        --- Purpose : Initialize by a Face.
    
    SplitSurface (me: mutable) 
    returns Boolean is redefined;
    	---Purpose: Performs splitting of surface and computes the shell
	--          from source face.
    
    SetNbSplitPoints(me: mutable; num: Integer);
    	---Purpose: Sets the number of cutting lines by which closed face 
        --          will be splitted. The resulting faces will be num+1.
    
    GetNbSplitPoints(me) returns Integer;
    	---Purpose: Returns the number of splitting points
  
fields

    myNbSplit: Integer;

end ClosedFaceDivide;
