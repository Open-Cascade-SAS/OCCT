-- Created on: 1993-07-06
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class CurveOnSurface from BRep inherits GCurve from BRep

	---Purpose: Representation  of a  curve   by a   curve  in the
	--          parametric space of a surface.

uses
    Pnt                 from gp,
    Pnt2d               from gp,
    Box2d               from Bnd,
    Curve               from Geom2d,
    Surface             from Geom,
    Location            from TopLoc,
    CurveRepresentation from BRep

is

    Create(PC : Curve    from Geom2d; 
    	   S  : Surface  from Geom; 
    	   L  : Location from  TopLoc)
    returns mutable CurveOnSurface from BRep;

    SetUVPoints(me : mutable; P1, P2 : Pnt2d from gp)
	---C++: inline
    is static;

    UVPoints(me; P1, P2 : out Pnt2d from gp)
	---C++: inline
    is static;
    
    D0(me; U : Real; P : out Pnt from gp);
	---Purpose: Computes the point at parameter U.

    IsCurveOnSurface(me) returns Boolean
	---Purpose: Returns True.
    is redefined;
    
    IsCurveOnSurface(me; S : Surface from Geom; L : Location from TopLoc) 
    returns Boolean
	---Purpose: A curve in the parametric space of a surface.
    is redefined;
    
    Surface(me) returns any Surface from Geom
	---C++: return const &
    is redefined;

    PCurve(me) returns any Curve from Geom2d
	---C++: return const &
    is redefined;

    PCurve(me : mutable; C : Curve from Geom2d)
    is redefined;

    Copy(me) returns mutable CurveRepresentation from BRep is virtual;
	---Purpose: Return a copy of this representation.

    Update(me : mutable)
	---Purpose: Recomputes any derived data after a modification.
	--          This is called when the range is modified.
    is redefined;

fields
    
    myPCurve      : Curve from Geom2d;
    mySurface     : Surface from Geom;
    myUV1         : Pnt2d from gp  is protected;
    myUV2         : Pnt2d from gp  is protected;

end CurveOnSurface;
