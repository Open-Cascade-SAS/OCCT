-- Created on: 1999-11-05
-- Created by: Vladislav ROMASHKO
-- Copyright (c) 1999-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Prism from QANewBRepNaming inherits TopNaming from QANewBRepNaming

    ---Purpose: To load the Prism results 

uses 
 
    MakePrism from BRepPrimAPI,
    Label     from TDF,
    Shape     from TopoDS

is
 
    Create returns Prism from QANewBRepNaming;
    
    Create(ResultLabel : Label from TDF) 
    returns Prism from QANewBRepNaming;

    Init(me : in out; ResultLabel : Label from TDF);
    

    Load (me; mkPrism : in out MakePrism from BRepPrimAPI;
	      basis   : in     Shape     from TopoDS);
    ---Purpose: Loads the prism in the data framework

    Bottom (me)
    ---Purpose : Returns the insertion label of the bottom face of the Prism.
    returns Label from TDF;

    Top (me)
    ---Purpose : Returns  the insertion label of the  top face of the Prism.
    returns Label  from TDF;

    Lateral (me)
    ---Purpose: Returns the insertion label of the lateral face of the Prism.
    returns Label from TDF;

    Degenerated (me)
    ---Purpose: Returns the insertion label of the degenerated face of the Prism.
    returns Label from TDF;

    Dangle (me)
    ---Purpose: Returns the insertion label of the degenerated face of the Prism.
    returns Label from TDF;

    Content (me)
    ---Purpose: Returns the insertion label of the degenerated face of the Prism.
    returns Label from TDF;

end Prism;
