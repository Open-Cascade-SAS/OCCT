-- Created on: 1994-10-03
-- Created by: Christian CAILLET
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class TransientListBinder  from Transfer  inherits Binder from Transfer

    ---Purpose : This binder binds several (a list of) Transients with a starting
    --           entity, when this entity itself corresponds to a simple list
    --           of Transients. Each part is not seen as a sub-result of an
    --           independant componant, but as an item of a built-in list

uses CString, Type,
	      HSequenceOfTransient from TColStd

raises TypeMismatch, OutOfRange

is

    Create returns mutable TransientListBinder;

    Create (list : mutable HSequenceOfTransient from TColStd)
    	 returns mutable TransientListBinder;

    IsMultiple (me) returns Boolean  is redefined;
    -- returns True if more than one result

    ResultType (me) returns Type;
    -- returns Standard_Transient

    ResultTypeName (me) returns CString;
    -- returns list(Standard_Transient)

    AddResult (me : mutable; res : Transient);
    ---Purpose : Adds an item to the result list

    Result (me) returns HSequenceOfTransient from TColStd;

    SetResult (me : mutable; num : Integer; res : Transient);
    ---Purpose : Changes an already defined sub-result

    NbTransients (me) returns Integer;

    Transient (me; num : Integer) returns Transient
    	raises OutOfRange;
    ---C++ : return const &


fields

    theres :  HSequenceOfTransient from TColStd;

end TransientListBinder;
