-- Created on: 1996-01-25
-- Created by: LAVNIKOV Alexey & PLOTNIKOV Eugeny
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class GraphicDevice from WNT inherits GraphicDevice from Aspect

    	---Purpose: This class defines Windows NT display device.
    	--          A Graphic Device defines color management. Windows can run in three
    	--          different color modes depending of the installed graphic board:
    	--           - Low color resolution which allows us to use 16 predefined pure
    	--             colors for drawing lines and unlimited number of dithered colors
    	--             for window's background, solid filled areas etc. Here Graphic Device
    	--             will approximate requested colors by existing ones for line colors
    	--             ( really this approximation is doing by Windows ). A dithering
    	--             technique will be used for window's backgrounds, solid fills etc.
    	--             ( this is doing by WIndows also ). A dithering techique will be use 
    	--             for solid fill.
    	--           - Medium color resolution which requires a Windows palette manager.
    	--             This mode takes after X window system's PseudoColor Visual. The
    	--             application can create a LOGICAL PALETTE to represent 20 reserved
    	--             by Windows colors and 236 programmable ones. It's possible to reserve
    	--             odd entries in the palette for highlighting purposes ( but real
    	--             technique is not the same as in X window system - see Windows manual ).
    	--             It's possible to create several logical palettes. To do it create
    	--             other GraphicDevice but in this case color "flicking" is possible.
    	--           - High color resolution. Here 65 536 or 16 777 216 colors are available.
    	--             Any color we like will be exactly displayed on the screen, but
    	--             highlighting technique is not available. This mode often called
    	--             TrueColor but it's not the same as X window TrueColor.
    	--          A Graphic Device also defines physical dimensions of the screen.

 uses

    Color         from Quantity,
    Length        from Quantity,
    ColorMap      from Aspect,
    Handle        from Aspect,
    ColorRef      from WNT,
    HColorTable   from WNT,
    Long          from WNT,
    GraphicDriver from Aspect

 raises

    GraphicDeviceDefinitionError from Aspect,
    BadAccess                    from Aspect

 is

    Create (
     aColorCube  : Boolean from Standard = Standard_False;
     aDevContext : Handle  from Aspect = 0
    )
     returns mutable GraphicDevice from WNT
	---Level:   Public
	---Purpose: Creates a GraphicDevice and logical palette.
	--          Builds an OpenGL colorcube on that palette depending
	--          of the aColorCube flag and hardware. 
	--  Warning: Raises if createion of the logical palette failed.
     raises GraphicDeviceDefinitionError from Aspect;

	Create (
	 aColorCube  : Boolean from Standard;
	 aDevContext : Integer from Standard
	) returns mutable GraphicDevice from WNT
	---Purpose: same as previous one (to provide access form CCL)
	  raises GraphicDeviceDefinitionError from Aspect;

    Destroy ( me : mutable ) is virtual;
	---Level:   Public
	---Purpose: Destroies all ressources attached to the GraphicDevice.
    	---C++:     alias ~

    SetColor (
     me         : mutable;
     aColor     : Color   from Quantity;
     aHighlight : Boolean from Standard = Standard_False
    )
     returns ColorRef from WNT is static;
    	---Level:   Public
    	---Purpose: Returns the color value in form specific to Windows NT.
    	--          Sets the color values in the logical palette if the
    	--          hardware supports it. If in this case there are not
    	--          free cell in the logical palette then this method will
    	--          search for nearest color in the palette.
    	--          If <aHighlight> is True then sets a highlight color.
           
    SetColor (
     me         : mutable;
     aRed       : Integer from Standard;
     aGreen     : Integer from Standard;
     aBlue      : Integer from Standard;
     aHighlight : Boolean from Standard = Standard_False
    )
     returns ColorRef from WNT is virtual;
	---Level:   Public
        ---Purpose: See above

    SetColor ( me : mutable; aPixel : Long from WNT )
     is virtual;
	---Level:   Internal
	---Purpose: Color allocation for images.

    MapColors (
     me          : mutable;
     aColorMap   : ColorMap           from Aspect;
     aColorTable : in out HColorTable from WNT
    ) is static;
    	---Level:   Public
    	---Purpose: Returns the color value in form specific to WIndows NT
    	--          in the <aColorTable>. See SetColor method.
    	--  Warning: The dimensions and index ranges of the <aColorMap> and
    	--          <aColorTable> must be the same; 

    HPalette ( me ) returns Handle from Aspect is static;
	---Level:   Public
	---Purpose: Returns logical palette handle attached to the
	--          GraphicDevice.
    	---C++:     inline

    DisplaySize ( me; aWidth, aHeight : out Integer from Standard ) is static;
	---Level:   Public
	---Purpose: Returns the Display size in PIXEL
        ---C++:     inline

    DisplaySize ( me; aWidth, aHeight : out Length from Quantity ) is static;
	---Level:   Public
	---Purpose: Returns the Display size in working units units
        ---C++:     inline

    IsPaletteDevice ( me ) returns Boolean from Standard is static;
    	---Level:   Public
    	---Purpose: Returns True if hardware is palette-compatible.
        ---C++:     inline

    NumColors ( me ) returns Integer from Standard is static;
    	---Level:   Public
    	---Purpose: Returns number of available colors.
        ---C++:     inline

    HighlightColor ( me ) returns ColorRef from WNT is static;
	---Level:   Public
	---Purpose: Returns highlight color.
        ---C++:     inline

    GraphicDriver ( me ) returns GraphicDriver from Aspect is redefined;
	---Level:   Public
	---Purpose: Dummy method

	Init (
	 me          : mutable; 
     aColorCube  : Boolean from Standard;
     aDevContext : Handle  from Aspect
	) is protected;

 fields

    myMWidth,
    myMHeight         : Length   from Quantity is protected;
    myWidth,
    myHeight,
    myNumColors       : Integer  from Standard is protected;
    myFreeIndex       : Integer  from Standard is protected;
    myPalette         : Handle   from Aspect   is protected;
    myLogPal          : Address  from Standard is protected;
    myHighlightColor  : ColorRef from WNT      is protected;
    myOpenGLPalette   : Boolean  from Standard is protected;

 friends

    class Window from WNT

end GraphicDevice;
