-- Created on: 1998-03-26
-- Created by: Robert COUBLANC
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



private class SortCriterion from SelectMgr 

    ---Purpose: This class provides data and criterion for sorting candidate
    --          entities in the process of interactive selection by mouse click

is
    Create returns SortCriterion from SelectMgr;

    Create(thePriority: Integer from Standard;
    	   theDepth, theMinDist, theTol: Real from Standard;
    	   PreferClosest: Boolean from Standard)
    returns SortCriterion from SelectMgr;
    ---Purpose: Defines parameters of selection criterion:
    -- - Priority: selection priority
    -- - Depth: distance from the view plane to the entity
    -- - MinDist: distance from the clicked point to the entity on the view plane
    -- - Tol: tolerance used for selecting candidates
    -- - PreferClosest: specify whether closest object is preferred even if 
    --                  if has less priority

    SetPriority (me : in out; P:Integer from Standard);
    ---C++: inline
    SetDepth    (me : in out; D:Real from Standard);
    ---C++: inline
    SetMinDist  (me : in out; D:Real from Standard);
    ---C++: inline
    SetTol (me : in out; T:Real from Standard);
    ---C++: inline

    Priority(me) returns Integer from Standard;
    ---C++: inline
    Depth(me) returns Real from Standard;
    ---C++: inline
    MinDist(me) returns Real from Standard;
    ---C++: inline
    Tol(me) returns Real from Standard;
    ---C++: inline


    IsGreater(me;anOtherCriterion:SortCriterion from SelectMgr)
    returns Boolean from Standard;
    ---C++: alias operator >

    IsLower(me;anOtherCriterion:SortCriterion from SelectMgr)
    returns Boolean from Standard;
    ---C++: alias operator <


fields
    myPrior: Integer from Standard;
    myDepth: Real    from Standard;
    myDist : Real    from Standard;
    myTol  : Real    from Standard;
    myPreferClosest: Boolean from Standard;
    
end SortCriterion;
