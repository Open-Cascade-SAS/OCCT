-- Created on: 2002-12-12
-- Created by: data exchange team
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class SurfaceSectionFieldVarying from StepElement
inherits SurfaceSectionField from StepElement

    ---Purpose: Representation of STEP entity SurfaceSectionFieldVarying

uses
    HArray1OfSurfaceSection from StepElement

is
    Create returns SurfaceSectionFieldVarying from StepElement;
	---Purpose: Empty constructor

    Init (me: mutable; aDefinitions: HArray1OfSurfaceSection from StepElement;
                       aAdditionalNodeValues: Boolean);
	---Purpose: Initialize all fields (own and inherited)

    Definitions (me) returns HArray1OfSurfaceSection from StepElement;
	---Purpose: Returns field Definitions
    SetDefinitions (me: mutable; Definitions: HArray1OfSurfaceSection from StepElement);
	---Purpose: Set field Definitions

    AdditionalNodeValues (me) returns Boolean;
	---Purpose: Returns field AdditionalNodeValues
    SetAdditionalNodeValues (me: mutable; AdditionalNodeValues: Boolean);
	---Purpose: Set field AdditionalNodeValues

fields
    theDefinitions: HArray1OfSurfaceSection from StepElement;
    theAdditionalNodeValues: Boolean;

end SurfaceSectionFieldVarying;
