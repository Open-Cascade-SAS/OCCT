-- File:	GeomToStep_MakeConicalSurface.cdl
-- Created:	Mon Jun 14 16:05:32 1993
-- Author:	Martine LANGLOIS
--		<mla@mastox>
---Copyright:	 Matra Datavision 1993

class MakeConicalSurface from GeomToStep inherits Root from GeomToStep

    ---Purpose: This class implements the mapping between class
    --          ConicalSurface from Geom and the class
    --          ConicalSurface from StepGeom which describes a
    --          conical_surface from Prostep
  
uses ConicalSurface from Geom,
     ConicalSurface from StepGeom
     
raises NotDone from StdFail
     
is 



Create ( CSurf : ConicalSurface from Geom ) returns MakeConicalSurface;

Value (me) returns ConicalSurface from StepGeom
    raises NotDone
    is static;
    ---C++: return const&

fields

    theConicalSurface : ConicalSurface from StepGeom;
    	-- The solution from StepGeom
    	
end MakeConicalSurface;


