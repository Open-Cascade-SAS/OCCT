-- File:	STEPControl.cdl
-- Created:	Tue Apr  9 10:33:36 1996
-- Author:	Christian CAILLET
--		<cky@paris1>
---Copyright:	 Matra Datavision 1996


package STEPControl

    ---Purpose : This package provides external access and control for STEP,
    --           especially to deal with Shapes

uses 
    Standard, 
    gp,
    TColStd, 
    TCollection,
    Interface, 
    Transfer, 
    IFSelect, 
    XSControl,
    TopoDS, 
    TopTools, 
    StepBasic, 
    StepData, 
    StepGeom, 
    StepShape, 
    StepRepr,
    STEPConstruct,
    TransferBRep,
    StepToTopoDS, -- Non-manifold topology: STEP -> TopoDS (ssv; 13.11.2010)
    MoniTool -- Non-manifold topology: TopoDS -> STEP (ssv; 13.11.2010)
is

    enumeration StepModelType is
    	AsIs,
    	ManifoldSolidBrep,
	BrepWithVoids,
	FacetedBrep,
	FacetedBrepAndBrepWithVoids,
	ShellBasedSurfaceModel,
	GeometricCurveSet,
	Hybrid
    end StepModelType;
        ---Purpose:  Gives you the choice of translation mode for an Open
--   CASCADE shape that is being translated to STEP.
--   - STEPControl_AsIs translates an Open CASCADE shape to its
--   highest possible STEP representation.
--   - STEPControl_ManifoldSolidBrep translates an Open CASCADE shape
--   to a STEP manifold_solid_brep or brep_with_voids entity.
--   - STEPControl_FacetedBrep translates an Open CASCADE shape
--   into a STEP faceted_brep entity.
-- -  STEPControl_ShellBasedSurfaceModel translates an Open CASCADE shape
--   into a STEP shell_based_surface_model entity.
--   - STEPControl_GeometricCurveSet
--   translates an Open CASCADE shape into a STEP geometric_curve_set entity.

    class Controller;

    class Reader;
    class Writer;

    class ActorRead;
    class ActorWrite;

end STEPControl;
