-- Created on: 2001-12-19
-- Created by: Sergey KUUL
-- Copyright (c) 2001-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MTHasher from MoniTool

	---Purpose: 
	-- The auxiliary class provides hash code for mapping objects   

is

    HashCode(myclass; Str : CString; Upper : Integer) returns Integer;
	---C++: inline
	---Purpose: Returns a HasCode value for the CString <Str>  in the
	-- range 0..Upper.
	-- Default ::HashCode(Str,Upper)
	
    IsEqual(myclass; Str1, Str2 : CString) returns Boolean;
	---C++: inline
	---Purpose: Returns True  when the two CString are the same. Two
	-- same strings must have the same hashcode, the
	-- contrary is not necessary.
	-- Default Str1 == Str2
	
end MTHasher;
