-- Created on: 1993-01-09
-- Created by: CKY / Contract Toubro-Larsen ( Deepak PRABHU )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


package IGESDefs

        ---Purpose : To embody general definitions of Entities
        --           (Parameters, Tables ...)

uses

        Standard,
        TCollection,
	TColStd,
	Message,
        Interface,
        IGESData,
        IGESBasic,
        IGESGraph

is

        class   AssociativityDef;
        -- Type 302, Form 5001-9999
        ---Purpose : This class permits the preprocessor to define an
        --           associativity schema. i.e., by using it preprocessor
        --           defines the type of relationship.

        class   MacroDef;
        -- Type 306, Form 0
        ---Purpose : This Class specifies the action of a specific MACRO.
        --           After specification MACRO can be used as necessary
        --           by means of MACRO class instance entity.

        class   UnitsData;
        -- Type 316, Form 0
        ---Purpose : This class stores data about a model's
        --           fundamental units.

        class   AttributeDef;
        -- Type 322, Form 0,1,2
        ---Purpose : This is class is used to support the concept of well
        --           defined collection of attributes, whether it is a table
        --           or a single row of attributes.

        class   TabularData;
        -- Type 406,  Form 11
        ---Purpose : This Class is used to provide a Structure to accomodate
        --           point form data.

        class   GenericData;
        -- Type 406,  Form 27
        ---Purpose : This Class is used to communicate information which is
        --           defined by the system operator while creating the model.
        --           The information is system specific and does not map into
        --           one of the predefined properties or associativities.
        --           Properties and property values can be defined by multiple
        --           instances of this property.

        class   AttributeTable;
        -- Type 422, Form 0,1
        ---Purpose : This class is used to represent an occurence of
        --           Attribute Table. This Class may be independent
        --           or dependent or pointed at by other Entities.

    	--    Tools for Entities    --

        class ToolAssociativityDef;
        class ToolMacroDef;
        class ToolUnitsData;
        class ToolAttributeDef;
        class ToolTabularData;
        class ToolGenericData;
        class ToolAttributeTable;

	-- Definition and Exploitation of Entities defined in this Package

        class Protocol;
	class ReadWriteModule;
	class GeneralModule;
	class SpecificModule;

        -- Instantiations

     class  Array1OfTabularData instantiates  Array1 from TCollection(TabularData);

     class HArray1OfTabularData instantiates HArray1 from TCollection
    	(TabularData,Array1OfTabularData);
     class HArray1OfHArray1OfTextDisplayTemplate instantiates
    --	HArray1 (HArray1OfTextDisplayTemplate,Array1OfHArray1OfTextDisplayTemplate);
      JaggedArray from Interface (HArray1OfTextDisplayTemplate from IGESGraph);

        -- Package Methods

    Init;
    ---Purpose : Prepares dynamic data (Protocol, Modules) for this package

    Protocol  returns Protocol from IGESDefs;
    ---Purpose : Returns the Protocol for this Package

end IGESDefs;
