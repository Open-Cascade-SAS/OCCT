-- Created on: 1991-07-24
-- Created by: Michel CHAUVAT
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

private generic class FuncExtCC from Extrema 
(Curve1    as any;
 Tool1     as any;-- as ToolCurve(Curve1);
 Curve2    as any;
 Tool2     as any;-- as ToolCurve(Curve2);
 POnC      as any;
 Pnt       as any;
 Vec       as any )
 
 
inherits FunctionSetWithDerivatives from math
    ---Purpose: Function allows finding extrema of the distance between 2 curves.

uses    Vector            from math,
	Matrix            from math,
	SequenceOfReal    from TColStd

raises  OutOfRange from Standard

private class SeqPOnC instantiates Sequence from TCollection(POnC);

is

    Create (thetol: Real = 1.0e-10) returns FuncExtCC;
    ---Purpose:

    Create (C1: Curve1; C2: Curve2; thetol: Real = 1.0e-10) returns FuncExtCC;
    ---Purpose:

    SetCurve (me: in out; theRank: Integer; C1: Curve1);
    ---Purpose:

    SetTolerance (me: in out; theTol: Real);
    ---C++: inline
    ---Purpose:

    NbVariables (me) returns Integer is redefined;
    ---C++: inline

    NbEquations (me) returns Integer is redefined;
    ---C++: inline

    Value (me: in out; UV: Vector; F: out Vector) returns Boolean is redefined;
    	---Purpose: Calculate Fi(U,V).

    Derivatives (me: in out; UV: Vector; DF: out Matrix)
    	returns Boolean;
    	---Purpose: Calculate Fi'(U,V).

    Values (me: in out; UV: Vector; F: out Vector; DF: out Matrix)
    	returns Boolean;
    	---Purpose: Calculate Fi(U,V) and Fi'(U,V).

    GetStateNumber (me: in out) returns Integer
    	---Purpose: Save the found extremum.
    	is redefined;

    NbExt (me) returns Integer;
        ---C++: inline
    	---Purpose: Return the number of found extrema.

    SquareDistance (me; N: Integer) returns Real
        ---C++: inline
    	---Purpose: Return the value of the Nth distance.
    	raises  OutOfRange;
	    	-- if N < 1 or N > NbExt(me).

    Points (me; N: Integer; P1,P2: out POnC)
    	---Purpose: Return the points of the Nth extreme distance.
    	raises  OutOfRange;
	    	-- if N < 1 or N > NbExt(me).

    CurvePtr (me; theRank: Integer) returns Address;
        ---C++: inline
        ---Purpose: Returns a pointer to the curve specified in the constructor
        --          or in SetCurve() method.

    Tolerance (me) returns Real;
        ---C++: inline
        ---Purpose: Returns a tolerance specified in the constructor
        --          or in SetTolerance() method.

    SubIntervalInitialize(me: in out; theUfirst, theUlast: Vector);
    	---Purpose: Determines of boundaries of subinterval for find of root.
    
    SearchOfTolerance(me: in out; C: Address from Standard) returns Real from Standard;
    	---Purpose: Computes a Tol value. If 1st derivative of curve
    	--          |D1|<Tol, it is considered D1=0.      


fields
    myC1    : Address from Standard;
    myC2    : Address from Standard;
    myTol   : Real;
    myU     : Real;        
    myV     : Real;        
    myP1    : Pnt;   -- current point C1(U)
    myP2    : Pnt;   -- current point C2(U)
    myDu    : Vec;   -- current D1 C1(U)
    myDv    : Vec;   -- current D1 C2(V)

    mySqDist: SequenceOfReal from TColStd;
    myPoints: SeqPOnC;

    myTolC1,myTolC2: Real from Standard;  -- toolerance for derivate

--Supremum of search 1st non-zero derivative    
    myMaxDerivOrderC1, myMaxDerivOrderC2: Integer from Standard;
    
--boundaries of subinterval for find of root
    myUinfium, myUsupremum: Real from Standard; -- C1 curve
    myVinfium, myVsupremum: Real from Standard; -- C2 curve


end FuncExtCC;
