-- Created on: 2000-05-18
-- Created by: Peter KURNEV
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

package BOPTest 
---Purpose: 

uses
    gp,
    Draw,
    DBRep, 
    TopAbs,    	     
    TopoDS,
    TopTools, 
    BOPCol,    
    BOPDS,    
    BOPAlgo 
     
is  
    
    class Objects; 
    class DrawableShape; 
    -- 
    AllCommands        (aDI:out Interpretor from Draw);
    BOPCommands        (aDI:out Interpretor from Draw); 
    CheckCommands      (aDI:out Interpretor from Draw); 
    TolerCommands      (aDI:out Interpretor from Draw); 
    LowCommands        (aDI:out Interpretor from Draw); 
    ObjCommands        (aDI:out Interpretor from Draw);
    PartitionCommands  (aDI:out Interpretor from Draw);
    Factory            (aDI:out Interpretor from Draw);
    
end BOPTest;
