-- Created on: 1998-04-02
-- Created by: Christian CAILLET
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SignLevelNumber  from IGESSelect    inherits Signature  from IFSelect

    ---Purpose : Gives D.E. Level Number under two possible forms :
    --           * for counter : "LEVEL nnnnnnn", " NO LEVEL", " LEVEL LIST"
    --           * for selection : "/nnn/", "/0/", "/1/2/nnn/"
    --           
    --           For matching, giving /nn/ gets any entity attached to level nn
    --           whatever simple or in a level list

uses CString, Transient, AsciiString, InterfaceModel

is

    Create (countmode : Boolean) returns SignLevelNumber;
    ---Purpose : Creates a SignLevelNumber
    --           <countmode> True : values are naturally displayed
    --           <countmode> False: values are separated by slashes
    --             in order to allow selection by signature by Draw or C++

    Value   (me; ent : any Transient; model : InterfaceModel) returns CString;
    ---Purpose : Returns the value (see above)

fields

    thecountmode : Boolean;

end SignLevelNumber;
