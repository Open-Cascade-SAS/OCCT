-- Created on: 1998-01-22
-- Created by: Sergey ZARITCHNY
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



deferred class EllipseRadiusDimension from AIS inherits Relation from AIS

	---Purpose: 
    	--  Computes  geometry  (  basis  curve  and  plane  of  dimension)
    	--  for  input  shape  aShape  from  TopoDS
	--  Root  class  for MinRadiusDimension  and  MaxRadiusDimension 
uses
     Shape                 from TopoDS,
     Elips                 from gp,
     Pnt                   from gp, 
     Pln                   from gp, 
     Curve                 from Geom,  
     OffsetCurve           from Geom,
     Ellipse               from Geom,
     Plane                 from Geom, 
     Surface               from Geom,
     ExtendedString        from TCollection,    
     KindOfSurface         from AIS,
     KindOfDimension       from AIS 

is
     Initialize(aShape      :  Shape           from  TopoDS; 
    	    	aText       :  ExtendedString  from  TCollection); 

    	--  Ellipse  radius  dimension  of  a  Shape  which  can  be  Edge 
    	--  or  Face  (planar  or  cylindrical(surface  of  extrusion  or 
    	--  surface  of  offset)) 		 

      

    KindOfDimension(me) returns KindOfDimension from AIS 
    is redefined;

    IsMovable(me) returns Boolean from Standard 
    is redefined;        


--
--     Computation private methods
-- 

    ComputeGeometry( me: mutable ) ;
--     is  private;  
      
    ComputeFaceGeometry(me: mutable)
    is private; 
     
    ComputeCylFaceGeometry(me: mutable;
    	    	     	aSurfType     : KindOfSurface  from  AIS; 
    	    	    	aSurf         : Surface  from  Geom; 
    	    	    	Offset        : Real     from  Standard )
    is private; 
     
    ComputePlanarFaceGeometry(me: mutable)
    is private; 
    
    ComputeEdgeGeometry(me: mutable)
    is private;
    
fields 

    myEllipse     :  Elips        from  gp        is  protected; 
    myFirstPar    :  Real         from  Standard  is  protected; 
    myLastPar     :  Real         from  Standard  is  protected;  
    myIsAnArc     :  Boolean      from  Standard  is  protected; 
    myOffsetCurve  : OffsetCurve  from  Geom      is  protected; 
    myOffset       : Real         from  Standard  is  protected; 
    myIsOffset     : Boolean      from  Standard  is  protected;  
     
end EllipseRadiusDimension;
