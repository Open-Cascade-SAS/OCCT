-- Created on: 1994-06-01
-- Created by: Christian CAILLET
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class UpdateLastChange  from IGESSelect  inherits ModelModifier from IGESSelect

    ---Purpose : Allows to Change the Last Change Date indication in the Header
    --           (Global Section) of IGES File. It is taken from the operating
    --           system (time of application of the Modifier).
    --           The Selection of the Modifier is not used : it simply acts as
    --           a criterium to select IGES Files to touch up.
    --           Remark : IGES Models noted as version before IGES 5.1 are in
    --           addition changed to 5.1

uses AsciiString from TCollection,
     IGESModel, CopyTool, ContextModif

is

    Create returns mutable UpdateLastChange;
    ---Purpose : Creates an UpdateLastChange, which uses the system Date

    Performing (me; ctx : in out ContextModif;
    	        target  : mutable IGESModel;
                TC      : in out CopyTool);
    ---Purpose : Specific action : only <target> is used : the system Date
    --           is set to Global Section Item n0 25. Also sets IGES Version
    --           (Item n0 23) to IGES5 if it was older.

    Label (me) returns AsciiString from TCollection;
    ---Purpose : Returns a text which is
    --           "Update IGES Header Last Change Date"

end UpdateLastChange;
