-- Created on: 1995-04-25
-- Created by: Marie Jose MARTZ
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package BRepToIGESBRep

    ---Purpose : Provides tools in order to transfer CAS.CADE entities
    --         to IGESBRep.

uses 
    Interface,
    IGESData,
    IGESBasic,
    IGESGeom,
    IGESSolid,
    Geom,
    Geom2d,
    GeomAbs,
    GeomToIGES,
    Geom2dToIGES,
    TColStd,
    TopoDS,
    TopTools,
    TopLoc,
    TopAbs,
    Transfer,
    TransferBRep,
    BRep,
    BRepTools, 
    gp,
    TCollection,
    BRepToIGES

is

--  ------------------------------------------------------
--  Package Classes
--  ------------------------------------------------------

    class Entity;


end BRepToIGESBRep;
