-- Created on: 1997-05-13
-- Created by: Fabien REUTER
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package  StlAPI 

    	 ---Purpose : Offers the API for STL data manipulation.
    	 --         

uses 
 
    TopoDS,
    StlMesh
     
is 
    class Writer; 
    class Reader; 
    
    Write(aShape      : in Shape from TopoDS;  
          aFile       : in CString from Standard;
    	  aAsciiMode  : in Boolean from Standard = Standard_True);
	  ---Purpose : Convert and write shape to STL format.
	  --         file is written in binary if aAsciiMode is False
	  --         otherwise it is written in Ascii (by default)

    Read(aShape      : in out Shape from TopoDS;  
          aFile      : CString from Standard);
	  ---Purpose : Create a shape from a STL format.

end  StlAPI;
