-- Created on: 2008-10-31
-- Created by: EPA
-- Copyright (c) 2008-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class FaceAttribute from BRepMesh inherits TShared from MMgt

    ---Purpose: auxiliary class for FastDiscret and FastDiscretFace classes

uses    
    Real          from Standard,
    Address       from Standard,
    ClassifierPtr from BRepMesh

is 

    Create returns mutable FaceAttribute from BRepMesh;

    GetDefFace(me:mutable) returns Real;
       ---C++: return &
       ---C++: inline    

    GetUMin(me:mutable) returns Real;
       ---C++: return &
       ---C++: inline

    GetVMin(me:mutable) returns Real;
       ---C++: return &
       ---C++: inline

    GetUMax(me:mutable) returns Real;
       ---C++: return &
       ---C++: inline

    GetVMax(me:mutable) returns Real;
       ---C++: return &
       ---C++: inline

    GetDeltaX(me:mutable) returns Real;
       ---C++: return &
       ---C++: inline

    GetDeltaY(me:mutable) returns Real;
       ---C++: return &
       ---C++: inline

    GetMinX(me:mutable) returns Real;
       ---C++: return &
       ---C++: inline

    GetMinY(me:mutable) returns Real;
       ---C++: return &
       ---C++: inline
       
    GetClassifier(me:mutable) returns ClassifierPtr from BRepMesh;
       ---C++: return &
       ---C++: inline

fields  
    mydefface   : Real          from Standard;
    myumin      : Real          from Standard;
    myumax      : Real          from Standard;
    myvmin      : Real          from Standard;
    myvmax      : Real          from Standard;
    mydeltaX    : Real          from Standard;
    mydeltaY    : Real          from Standard;
    myminX      : Real          from Standard;
    myminY      : Real          from Standard;
    myclassifier: ClassifierPtr from BRepMesh;

end FaceAttribute;
