-- Created on: 1993-01-09
-- Created by: CKY / Contract Toubro-Larsen ( Kiran )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SplineSurface from IGESGeom  inherits IGESEntity

        ---Purpose: defines IGESSplineSurface, Type <114> Form <0>
        --          in package IGESGeom
        --          A parametric spline surface is a grid of polynomial
        --          patches. Patch could be of the type Linear, Quadratic,
        --          Cubic, Wilson-Fowler, Modified Wilson-Fowler, B-Spline
        --          The M * N grid of patches is defined by the 'u' break
        --          points TU(1), TU(2), ..., TU(M+1) and the 'v' break
        --          points TV(1), TV(2), TV(3) ..., TV(N+1).

uses

        Pnt           from gp,
        HArray1OfReal from TColStd,
        HArray2OfReal from TColStd,
        HArray2OfHArray1OfReal from IGESBasic

raises DimensionMismatch, OutOfRange

is

        Create returns mutable SplineSurface;

        -- Specific Methods pertaining to the class

        Init (me                              : mutable;
           aBoundaryType, aPatchType          : Integer;
           allUBreakpoints, allVBreakpoints   : HArray1OfReal;
           allXCoeffs, allYCoeffs, allZCoeffs : HArray2OfHArray1OfReal)
        raises DimensionMismatch;
        ---Purpose : This method is used to set the fields of the class
        --           SplineSurface
        --       - aBoundaryType   : Type of Spline boundary
        --                           1 = Linear
        --                           2 = Quadratic
        --                           3 = Cubic
        --                           4 = Wilson-Fowler
        --                           5 = Modified Wilson-Fowler
        --                           6 = B-spline
        --       - aPatchType      : Type of patch contained in the grid
        --                           1 = Cartesian Product
        --                           0 = Unspecified
        --       - allUBreakpoints : u values of grid lines
        --       - allVBreakpoints : v values of grid lines
        --       - allXCoeffs      : X coefficients of M x N patches
        --       - allYCoeffs      : Y coefficients of M x N patches
        --       - allZCoeffs      : Z coefficients of M x N patches
        -- raises exception if allXCoeffs, allYCoeffs & allZCoeffs are not
        -- of the same size.
        -- or if the size of each element of the double array is not 16

        NbUSegments(me) returns Integer;
        ---Purpose : returns the number of U segments

        NbVSegments(me) returns Integer;
        ---Purpose : returns the number of V segments

        BoundaryType(me) returns Integer;
        ---Purpose : returns boundary type

        PatchType(me) returns Integer;
        ---Purpose : returns patch type

        UBreakPoint(me; anIndex : Integer) returns Real
        raises OutOfRange;
        ---Purpose : returns U break point of the grid line referred to by anIndex
        -- raises exception if anIndex <= 0 or anIndex > NbUSegments() + 1

        VBreakPoint(me; anIndex : Integer) returns Real
        raises OutOfRange;
        ---Purpose : returns V break point of the grid line referred to by anIndex
        -- raises exception if anIndex <= 0 or anIndex > NbVSegments() + 1

        XPolynomial(me; anIndex1, anIndex2 : Integer) returns HArray1OfReal
        raises OutOfRange;
        ---Purpose : returns X polynomial of patch referred to by anIndex1, anIndex2
        -- raises exception if anIndex1 <= 0 or anIndex1 > NbUSegments()
        --                  or anIndex2 <= 0 or anIndex2 > NbVSegments()

        YPolynomial(me; anIndex1, anIndex2 : Integer) returns HArray1OfReal
        raises OutOfRange;
        ---Purpose : returns Y polynomial of patch referred to by anIndex1, anIndex2
        -- raises exception if anIndex1 <= 0 or anIndex1 > NbUSegments()
        --                  or anIndex2 <= 0 or anIndex2 > NbVSegments()

        ZPolynomial(me; anIndex1, anIndex2 : Integer) returns HArray1OfReal
        raises OutOfRange;
        ---Purpose : returns Z polynomial of patch referred to by anIndex1, anIndex2
        -- raises exception if anIndex1 <= 0 or anIndex1 > NbUSegments()
        --                  or anIndex2 <= 0 or anIndex2 > NbVSegments()

    	Polynomials (me; XCoef, YCoef, ZCoef : out HArray2OfHArray1OfReal);
	---Purpose : returns in one all the polynomial values "in bulk"
	--           usefull for massive treatements

fields

--
-- Class    : IGESGeom_SplineSurface
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class SplineSurface.
--
-- Reminder : A SplineSurface instance is defined by :
--            Spline boundary type, the type of patches in the grid
--            the number of U, V segments, the break points, the X, Y, Z
--            polynomials for each patch.

        theBoundaryType : Integer;
        thePatchType    : Integer;
        theUBreakPoints : HArray1OfReal;
        theVBreakPoints : HArray1OfReal;
        theXCoeffs      : HArray2OfHArray1OfReal;
            -- each element of the HArray2 is of size 16
            -- the HArray2 is of size MN where M is the number of
            -- U segments and N is the number of V segments
        theYCoeffs      : HArray2OfHArray1OfReal;
            -- each element of the HArray2 is of size 16
            -- the HArray2 is of size MN where M is the number of
            -- U segments and N is the number of V segments
        theZCoeffs      : HArray2OfHArray1OfReal;
            -- each element of the HArray2 is of size 16
            -- the HArray2 is of size  MN where M is the number of
            -- U segments and N is the number of V segments

end SplineSurface;
