-- Created on: 1997-02-12
-- Created by: Alexander BRIVIN
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Rotation from Vrml 

	---Purpose:  defines a Rotation node of VRML specifying matrix and transform properties.
    	--  This  node  defines  a  3D  rotation  about  an  arbitrary  axis  through  the  origin. 
    	--  By  default  :  myRotation  =  (0 0 1 0)

uses
 
    SFRotation  from  Vrml

is
 
    Create returns   Rotation from Vrml;

    Create  (  aRotation  :  SFRotation  from  Vrml ) 
    	returns   Rotation from Vrml;
      
    SetRotation ( me : in out; aRotation : SFRotation  from  Vrml );
    Rotation ( me )  returns  SFRotation  from  Vrml;

    Print  ( me;  anOStream: in out OStream from Standard) returns OStream from Standard;
    ---C++:  return  & 

fields
 
    myRotation  :  SFRotation  from  Vrml; -- Rotation

end Rotation;
