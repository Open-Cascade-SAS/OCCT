-- Created on: 1995-02-22
-- Created by: Mister rmi
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

--Modified by Rob Jan 13 th  98 : Compute Depth on EyeLine for
--                                Each Kind of SensitiveEntity. 
--                                (Deferred Method to be implemented)


package Select3D 

	---Purpose: The Select3D package provides the following services
    	-- -   definition of standard   3D sensitive primitives such as points, curves and faces.
    	-- -   recovery of the bounding boxes in the 2D graphic selection space, if required.
    	-- -   a 3D-2D projector.

uses
    Standard,
    TCollection,
    TColStd,
    TColgp,
    gp,
    Bnd,
    Poly,
    TopLoc,
    Geom,
    SelectBasics,
    V3d

is
    
    ---Category: sensitive entities

    enumeration TypeOfSensitivity is TOS_INTERIOR,TOS_BOUNDARY,TOS_EXTERIOR
    end TypeOfSensitivity;
    	---Purpose: Provides values for type of sensitivity in 3D.
    	-- These are used to specify whether it is the interior,
    	-- the boundary, or the exterior of a 3D sensitive entity which is sensitive.

    deferred class SensitiveEntity;
    
    deferred class SensitivePoly;

    class SensitivePoint;

    class SensitiveSegment;

    class SensitiveCircle;

    class SensitiveCurve;

    class SensitiveTriangle; 

    class SensitiveTriangulation;

    class SensitiveFace;

    class SensitiveBox;

    class SensitiveWire;

    class SensitiveGroup;

    class SensitiveEntitySequence instantiates Sequence from TCollection 
    	(SensitiveEntity from Select3D);

    ---Category: selectors/projectors

    class Projector;


    class ListOfSensitiveTriangle instantiates List from TCollection
    (SensitiveTriangle from Select3D);

    class ListOfSensitive instantiates List from TCollection
    (SensitiveEntity from Select3D);

    imported Pnt;
    imported Pnt2d;
    imported Box2d;
    imported PointData;

end Select3D;
