-- Created on: 1993-10-19
-- Created by: Gerard GRAS
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

--		corrections MFA 21 Oct 94

class GraphicDevice from Xw inherits GraphicDevice from Aspect

	---Purpose: This class defines an X11 Graphic Device 
	--  Warning: An Graphic Device is defined by :
	--		- a connection "host:server.screen"
	--		- a colormap mapping of type Xw_TOM_xxxxx
	--		- a "UseDefault" flag which permits the use of the 
	--			DefaultColormap if possible.
	--	    The connection can be specified directly
	--	    or extracted from an existing Window.
	--	    All Xw_Windows may share the same Graphic Device if
	--	    you don't want to have any side effects on the stations
	--	    which have only one hardware pseudo-colormap .
	--	    Four kind of mapping are possible :
	--	    1) Xw_TOM_SIMPLERAMP
	--	       Allocates the number of required colors in the
	--	       colormap.
	--	       The number of user colors depends directly on
	--	       the hardware colormap size if UseDefault is False,
	--	       or on the remainding free colors in the hardware colormap
	--	       if UseDefault is True.
	--	    2) Xw_TOM_BESTRAMP
	--	       Allocates the number of required colors in the
	--	       colormap but leaves the Odd color indexes free
	--	       if possible for highlight color management.
        --	       (plane 0 is reserved for this usage)
	--	       The number of user colors depends directly on
	--	       the hardware colormap size if UseDefault is False,
	--	       or on the remainding free colors in the hardware colormap
	--	       if UseDefault is True.
	--	    3) Xw_TOM_COLORCUBE (the default)
	--	       Allocates the maximum available colors in the colormap
	--	       and builds a colorcube at this place.
	--	       Any user color will be approximate and will be chosen as
	--	       the nearest of the set of available colorcube colors.
	--	       In this case the number of user colors can be unlimited.
	--	    4) Xw_TOM_HARDWARE
	--	       May do serious damage to the color system.
	--	       Must be used for maintenance only.
	--	    5) Xw_TOM_READONLY
	--	       Allocates the number of required read only colors in the
	--	       default colormap.
	--	       The number of user colors depends directly on
	--	       the hardware colormap size. 

	---References:

uses

	AsciiString	from TCollection,
	Length		from Quantity,
	GraphicDriver	from Aspect,
	ColorMap	from Xw,
	TypeMap		from Xw,
	WidthMap	from Xw,
	FontMap		from Xw,
	MarkMap		from Xw,
	TypeOfVisual	from Xw,
	TypeOfMapping	from Xw,
	Handle		from Aspect

raises

	GraphicDeviceDefinitionError	from Aspect,
	BadAccess			from Aspect

is

	Create
	returns mutable GraphicDevice from Xw is protected ;

	Create (Connection	: CString from Standard ;
		Mapping		: TypeOfMapping from Xw = Xw_TOM_COLORCUBE ;
		Ncolors		: Integer from Standard = 0 ;
		UseDefault	: Boolean from Standard = Standard_True )
	returns mutable GraphicDevice from Xw
	---Level: Public
	---Purpose: Create an Graphic Device on the specified Connection
	--	    by using ALL screen defaults if possible
	--	    (i.e:Default Colormap)
	--  Warning: Raises if the Device is Badly defined
	raises GraphicDeviceDefinitionError from Aspect ;

	---------------------------------------------------
	-- Category: methods to modify the class definition
	---------------------------------------------------

	Destroy ( me : mutable )
	---Level: Public
	---Purpose: Destroies all ressources attached to the GraphicDevice
	--	    (Windows, Colormaps, ....)
	--  Warning: Raises if the Device is Badly defined
	raises BadAccess from Aspect is virtual;
	---C++: alias ~
	---Category: methods to modify the class definition

	InitMaps ( me : mutable ; Connection : CString from Standard ;
				  Mapping   : TypeOfMapping from Xw ;
				  Ncolors   : Integer from Standard ;
				  UseDefault: Boolean from Standard )
	---Level: Public
	---Purpose: Initializes all ressources attached to the GraphicDevice
	--  Category: methods to modify the class definition
	--  Warning: Raises if the Device is Badly defined
	raises GraphicDeviceDefinitionError from Aspect
	is static protected ;

	----------------------------
	-- Category: Inquire methods
	----------------------------

	ColorMap2D ( me )
	returns ColorMap from Xw is static;
	---Level: Internal
	---Purpose: Returns the 2D oriented Device color map.
	---Category: Inquire methods

	VisualClass2D ( me )
	returns TypeOfVisual from Xw is static;
	---Level: Internal
	---Purpose: Returns the 2D oriented Visual Class.
	---Category: Inquire methods

	OverlayVisualClass2D ( me )
	returns TypeOfVisual from Xw is static;
	---Level: Internal
	---Purpose: Returns the 2D oriented overlay Visual Class.
	---Category: Inquire methods

	ExtendedColorMap2D ( me )
	returns Address from Standard
	is static protected ;
	---Level: Internal
	---Purpose: Returns extended data colormap 2D structure pointer.
	---Category: Inquire methods

	ExtendedOverlayColorMap2D ( me )
	returns Address from Standard
	is static protected ;
	---Level: Internal
	---Purpose: Returns extended data overlay colormap 2D structure pointer.
	---Category: Inquire methods

	ColorMap3D ( me )
	returns ColorMap from Xw is static;
	---Level: Internal
	---Purpose: Returns the 3D oriented Device color map.
	---Category: Inquire methods

	VisualClass3D ( me )
	returns TypeOfVisual from Xw is static;
	---Level: Internal
	---Purpose: Returns the 3D oriented Visual Class.
	---Category: Inquire methods

	OverlayVisualClass3D ( me )
	returns TypeOfVisual from Xw is static;
	---Level: Internal
	---Purpose: Returns the 3D oriented overlay Visual Class.
	---Category: Inquire methods

	ExtendedColorMap3D ( me )
	returns Address from Standard
	is static protected ;
	---Level: Internal
	---Purpose: Returns extended data colormap 3D structure pointer.
	---Category: Inquire methods

	ExtendedOverlayColorMap3D ( me )
	returns Address from Standard
	is static protected ;
	---Level: Internal
	---Purpose: Returns extended data overlay colormap 3D structure pointer.
	---Category: Inquire methods

	TypeMap ( me )
	returns TypeMap from Xw is static;
	---Level: Internal
	---Purpose: Returns the Device Type map.
	---Category: Inquire methods

	ExtendedTypeMap ( me )
	returns Address from Standard
	is static protected ;
	---Level: Internal
	---Purpose: Returns extended data typemap structure pointer.
	---Category: Inquire methods

	WidthMap ( me )
	returns WidthMap from Xw is static;
	---Level: Internal
	---Purpose: Returns the Device Width map.
	---Category: Inquire methods

	ExtendedWidthMap ( me )
	returns Address from Standard
	is static protected ;
	---Level: Internal
	---Purpose: Returns extended data widthmap structure pointer.
	---Category: Inquire methods

	FontMap ( me )
	returns FontMap from Xw is static;
	---Level: Internal
	---Purpose: Returns the Device Font map.
	---Category: Inquire methods

	ExtendedFontMap ( me )
	returns Address from Standard
	is static protected ;
	---Level: Internal
	---Purpose: Returns extended data fontmap structure pointer.
	---Category: Inquire methods

	MarkMap ( me )
	returns MarkMap from Xw is static;
	---Level: Internal
	---Purpose: Returns the Device Mark map.
	---Category: Inquire methods

	ExtendedMarkMap ( me )
	returns Address from Standard
	is static protected ;
	---Level: Internal
	---Purpose: Returns extended data markmap structure pointer.
	---Category: Inquire methods

	Display ( me )
	returns CString from Standard is static;
	---Level: Internal
	---Purpose: Returns the Device connection string.
	---Category: Inquire methods

	XDisplay ( me )
	returns Address from Standard is static;
	---Level: Internal
	---Purpose: Returns the Device Display Address.
	---Category: Inquire methods

	ExtendedDisplay ( me )
	returns Address from Standard
	is static protected ;
	---Level: Internal
	---Purpose: Returns extended data display structure pointer.
	---Category: Inquire methods

	DisplaySize ( me ; Width, Height : out Integer from Standard )
	---Level: Public
	---Purpose: Returns the Display size in PIXEL
	--  Warning: Raises if the connection is not defined properly
	raises BadAccess from Aspect is static;

	DisplaySize ( me ; Width, Height : out Length from Quantity )
	---Level: Public
	---Purpose: Returns the Display size in METER
	--  Warning: Raises if the connection is not defined properly
	raises BadAccess from Aspect is static;

	PlaneLayer ( me ; aVisualID : Integer from Standard )
	returns Integer from Standard
	---Level: Public
	---Purpose: Returns the plane layer ID from a visual ID
	--  Warning: Raises if the connection is not defined properly
	raises BadAccess from Aspect is static;

	GraphicDriver ( me )
		returns GraphicDriver from Aspect
		is redefined;

fields

	MyDisplay 		: AsciiString from TCollection ;
	MyColorMap2D		: ColorMap from Xw ;
	MyColorMap3D		: ColorMap from Xw ;
	MyTypeMap		: TypeMap from Xw ;
	MyWidthMap		: WidthMap from Xw ;
	MyFontMap		: FontMap from Xw ;
	MyMarkMap		: MarkMap from Xw ;
	MyExtendedDisplay	: Address from Standard is protected ;

friends

	class Window from Xw

end GraphicDevice from Xw ;
