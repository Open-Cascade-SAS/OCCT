-- Created on: 1994-11-30
-- Created by: Frederic MAUPAS
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MakeStepVertex from TopoDSToStep 
    inherits Root from TopoDSToStep

    ---Purpose: This class implements the mapping between classes 
    --          Vertex from TopoDS and TopologicalRepresentationItem from
    --          StepShape. 
  
uses Vertex                        from TopoDS,
     TopologicalRepresentationItem from StepShape,
     Tool                          from TopoDSToStep,
     MakeVertexError               from TopoDSToStep,
     FinderProcess                 from Transfer
          
raises NotDone from StdFail
     
is 

    Create returns MakeStepVertex;
    
    Create (V : Vertex from TopoDS;
    	    T : in out Tool from TopoDSToStep;
	   FP : mutable FinderProcess from Transfer)
         returns MakeStepVertex;
    
    Init(me : in out;
     	 V  : Vertex from TopoDS;
     	 T  : in out Tool from TopoDSToStep;
         FP : mutable FinderProcess from Transfer);

	    
    Value (me) returns TopologicalRepresentationItem from StepShape
    	raises NotDone
    	is static;
    	---C++: return const&
        
    Error(me) returns MakeVertexError from TopoDSToStep;

fields

    myResult : TopologicalRepresentationItem from StepShape;

    myError  : MakeVertexError from TopoDSToStep;
    
end MakeStepVertex;


