-- File:	GeomPlate_MakeApprox.cdl
-- Created:	Wed Mar  5 11:49:39 1996
-- Author:	Joelle CHAUVET
--		<jct@sgi38>
---Copyright:	 Matra Datavision 1996

class MakeApprox from GeomPlate
---Purpose:
-- Allows you to convert a GeomPlate surface into a BSpline.
uses

    Surface        from GeomPlate,
    BSplineSurface from Geom, 
    Shape          from GeomAbs,
    Criterion      from AdvApp2Var


is
    Create(SurfPlate: Surface from GeomPlate;
    	   PlateCrit: Criterion from AdvApp2Var;
    	   Tol3d: Real;
    	   Nbmax: Integer; 
    	   dgmax: Integer; 
     	   Continuity:  Shape  from  GeomAbs  =  GeomAbs_C1;
	   EnlargeCoeff : Real from Standard = 1.1)
    returns MakeApprox;
    ---Purpose:  Converts SurfPlate into a Geom_BSplineSurface with
    --  n Bezier pieces (n<=Nbmax) of degree <= dgmax 
    --  and an approximation error < Tol3d if possible
    --  the criterion CritPlate is satisfied if possible
    
    Create(SurfPlate: Surface from GeomPlate;
    	   Tol3d: Real;
    	   Nbmax: Integer; 
    	   dgmax: Integer;
    	   dmax : Real;
    	   CritOrder: Integer = 0; 
           Continuity:  Shape  from  GeomAbs  =  GeomAbs_C1;
	   EnlargeCoeff : Real from Standard = 1.1)
    returns MakeApprox;
    ---Purpose:  Converts SurfPlate into a Geom_BSplineSurface with
    --  n Bezier pieces (n<=Nbmax) of degree <= dgmax 
    --  and an approximation error < Tol3d if possible
    --  if CritOrder = -1 , no criterion is used
    --  if CritOrder = 0 , a PlateG0Criterion is used with max value > 10*dmax
    --  if CritOrder = 1 , a PlateG1Criterion is used with max value > 10*dmax
    --  WARNING : for CritOrder = 0 or 1, only the constraints points of SurfPlate
    --            are used to evaluate the value of the criterion
    
    Surface(me) returns BSplineSurface from Geom;
    ---Purpose: Returns the BSpline surface extracted from the
    --          GeomPlate_MakeApprox object.   
    
    ApproxError(me) returns Real;
    ---Purpose: Returns the error in computation of the approximation
    --          surface. This is the distance between the entire target
    --          BSpline surface and the entire original surface
    --          generated by BuildPlateSurface and converted by GeomPlate_Surface.    
    CriterionError(me) returns Real;
    ---Purpose: Returns the criterion error in computation of the
    --          approximation surface. This is estimated relative to the
    --          curve and point constraints only.
fields

    myPlate : Surface from GeomPlate;
    mySurface : BSplineSurface from Geom;
    myAppError,myCritError : Real;

end;
