-- File:        ConversionBasedUnitAndLengthUnit.cdl
-- Created:     Mon Dec  4 12:02:37 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWConversionBasedUnitAndLengthUnit from RWStepBasic

	---Purpose : Read & Write Module for ConversionBasedUnitAndLengthUnit

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     ConversionBasedUnitAndLengthUnit from StepBasic,
     EntityIterator from Interface

is

	Create returns RWConversionBasedUnitAndLengthUnit;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable ConversionBasedUnitAndLengthUnit from StepBasic);

	WriteStep (me; SW : in out StepWriter; ent : ConversionBasedUnitAndLengthUnit from StepBasic);

	Share(me; ent : ConversionBasedUnitAndLengthUnit from StepBasic; iter : in out EntityIterator);

end RWConversionBasedUnitAndLengthUnit;
