-- Created on: 1993-03-24
-- Created by: JCV
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class VectorWithMagnitude from Geom2d inherits Vector from Geom2d

        --- Purpose :
        --  Defines a vector with magnitude.
        --  A vector with magnitude can have a zero length.

uses Pnt2d     from gp,
     Trsf2d    from gp,
     Vec2d     from gp,
     Geometry  from Geom2d

raises ConstructionError from Standard

is


  Create (V : Vec2d) returns mutable VectorWithMagnitude;
        --- Purpose : Creates a persistent copy of V.


  Create (X, Y : Real)   returns mutable VectorWithMagnitude;
        --- Purpose : Creates a vector with two cartesian coordinates. 


  Create (P1, P2 : Pnt2d)   returns mutable VectorWithMagnitude;
        --- Purpose :
        --  Creates a vector from the point P1 to the point P2.
        --  The magnitude of the vector is the distance between P1 and P2



  SetCoord (me : mutable; X, Y : Real);
        --- Purpose :  Set <me> to X, Y coordinates.


  SetVec2d (me : mutable; V : Vec2d);
        -- Purpose : Set <me> to V.X(), V.Y() coordinates.


  SetX (me : mutable; X : Real);
        --- Purpose : Changes the X coordinate of <me>.


  SetY (me : mutable; Y : Real);
        --- Purpose :  Changes the Y coordinate of <me>


  Magnitude (me)  returns Real;
        --- Purpose : Returns the magnitude of <me>.


  SquareMagnitude (me)  returns Real;
        --- Purpose : Returns the square magnitude of <me>.


  Add (me : mutable; Other : Vector);
        --- Purpose :
        --  Adds the Vector Other to <me>.
        ---C++: alias operator +=


  Added (me; Other : Vector)  returns mutable VectorWithMagnitude
        --- Purpose :
        --  Adds the vector Other to <me>.
        ---C++: alias operator +
     is static;


  Crossed (me; Other : Vector)  returns Real;
        --- Purpose :
        --  Computes the cross product  between <me> and Other 
        --  <me> ^ Other. A new vector is returned.
        ---C++: alias operator ^


  Divide (me : mutable; Scalar : Real);
        --- Purpose : Divides <me> by a scalar.
        ---C++: alias operator /=


  Divided (me; Scalar : Real)  returns mutable VectorWithMagnitude
        --- Purpose :
        --  Divides <me> by a scalar. A new vector is returned.
        ---C++: alias operator /
     is static;


  Multiplied (me; Scalar : Real)  returns mutable VectorWithMagnitude
        --- Purpose :
        --  Computes the product of the vector <me> by a scalar.
        --  A new vector is returned.
        --  
        --  -C++: alias operator * 
        --  Collision with same operator defined for the class Vector!
     is static;


  Multiply (me : mutable; Scalar : Real);
        --- Purpose : 
        --  Computes the product of the vector <me> by a scalar.
        ---C++: alias operator *=


  Normalize (me : mutable)
        --- Purpose : Normalizes <me>.
     raises ConstructionError;
        --- Purpose : 
        --  Raised if the magnitude of the vector is lower or equal to
        --  Resolution from package gp.


  Normalized (me)  returns mutable VectorWithMagnitude
        --- Purpose : Returns a copy of <me> Normalized.
     raises ConstructionError
        --- Purpose :
        --  Raised if the magnitude of the vector is lower or equal to
        --  Resolution from package gp.
     is static;


  Subtract (me : mutable; Other : Vector);
        --- Purpose : Subtracts the Vector Other to <me>.
        ---C++: alias operator -=


  Subtracted (me; Other : Vector)  returns mutable VectorWithMagnitude
        --- Purpose :
        --  Subtracts the vector Other to <me>. A new vector is returned.
        ---C++: alias operator -
     is static;



  Transform (me: mutable; T : Trsf2d);
    	---Purpose: Applies the transformation T to this vector.


  Copy (me)  returns mutable like me;
    	--- Purpose: Creates a new object which is a copy of this vector.    
end;


