-- Created on: 1993-01-20
-- Created by: Laurent PAINNOT
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred generic class MLineTool from AppParCurves (MLine  as any)

    ---Purpose: Template which defines all the services relative to
    --          a MultiLine for approximation algorithms.


uses Pnt           from gp,
     Pnt2d         from gp,
     Vec           from gp,
     Vec2d         from gp,
     Array1OfPnt   from TColgp,
     Array1OfPnt2d from TColgp,
     Array1OfVec   from TColgp,
     Array1OfVec2d from TColgp

is
    
    
    FirstPoint(myclass; ML: MLine) returns Integer;
    	---Purpose: Returns the first index of multipoints of the MLine.


    LastPoint(myclass; ML: MLine) returns Integer;
    	---Purpose: Returns the last index of multipoints of the MLine.



    NbP2d(myclass; ML: MLine) returns Integer;
    	---Purpose: Returns the number of 2d points of a MLine.


    NbP3d(myclass; ML: MLine) returns Integer;
    	---Purpose: Returns the number of 3d points of a MLine.



    Value(myclass; ML: MLine; MPointIndex: Integer; tabPt: out Array1OfPnt);
    	---Purpose: returns the 3d points of the multipoint <MPointIndex>
    	--          when only 3d points exist.


    Value(myclass; ML: MLine; MPointIndex: Integer; 
          tabPt2d: out Array1OfPnt2d);
    	---Purpose: returns the 2d points of the multipoint <MPointIndex>
    	--          when only 2d points exist.


    Value(myclass; ML: MLine; MPointIndex: Integer; 
          tabPt: out Array1OfPnt; tabPt2d: out Array1OfPnt2d);
    	---Purpose: returns the 3d and 2d points of the multipoint 
    	--          <MPointIndex>.


    Tangency(myclass; ML: MLine; MPointIndex: Integer; tabV: out Array1OfVec)
    returns Boolean;
    	---Purpose: returns the 3d points of the multipoint <MPointIndex>
    	--          when only 3d points exist.


    Tangency(myclass; ML: MLine; MPointIndex: Integer; 
          tabV2d: out Array1OfVec2d)
    returns Boolean;
    	---Purpose: returns the 2d tangency points of the multipoint 
    	--          <MPointIndex> only when 2d points exist.


    Tangency(myclass; ML: MLine; MPointIndex: Integer; 
             tabV: out Array1OfVec; tabV2d: out Array1OfVec2d)
    returns Boolean;
    	---Purpose: returns the 3d and 2d points of the multipoint 
    	--          <MPointIndex>.





end MLineTool;    
