-- File:        PresentationStyleSelect.cdl
-- Created:     Fri Dec  1 11:11:11 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993



class PresentationStyleSelect from StepVisual inherits SelectType from StepData

	-- <PresentationStyleSelect> is an EXPRESS Select Type construct translation.
	-- it gathers : PointStyle, CurveStyle, SurfaceStyleUsage, SymbolStyle, FillAreaStyle, TextStyle
	-- Rev4 : only remain PointStyle, CurveStyle, SurfaceStyleUsage

uses

	PointStyle,
	CurveStyle,
	SurfaceStyleUsage
--	SymbolStyle,
--	FillAreaStyle,
--	TextStyle
is

	Create returns PresentationStyleSelect;
	---Purpose : Returns a PresentationStyleSelect SelectType

	CaseNum (me; ent : Transient) returns Integer;
	---Purpose: Recognizes a PresentationStyleSelect Kind Entity that is :
	--        1 -> PointStyle
	--        2 -> CurveStyle
	--        3 -> SurfaceStyleUsage
	--        4 -> SymbolStyle
	--        5 -> FillAreaStyle
	--        6 -> TextStyle
	--        0 else

	PointStyle (me) returns any PointStyle;
	---Purpose : returns Value as a PointStyle (Null if another type)

	CurveStyle (me) returns any CurveStyle;
	---Purpose : returns Value as a CurveStyle (Null if another type)

	SurfaceStyleUsage (me) returns any SurfaceStyleUsage;
	---Purpose : returns Value as a SurfaceStyleUsage (Null if another type)

end PresentationStyleSelect;

