-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

---Version:	 1.2 

--  Version	Date		Purpose
--         	Feb  3 1995	Creation
--         	Dec  15 1996    Version CSFDB

package ObjMgt 

---Purpose: This package defines services to manage the storage grain of data 
--          produced by applications and those classes to manage persistent 
--          extern reference.

uses

    PCollection,
    Storage,
    CDM,PCDM, TCollection

is

    --deferred class RetrievalDriver;
    ---Purpose: to retrieve ExternShareable objects in the framework.
 

    deferred class ExternShareable;
    ---Purpose: Defines the root persistent object which can be persistent 
    --          extern reference.

    private class ExternRef;
    ---Purpose: Defines (objet-relais) to implement extern reference.

    private class PSeqOfExtRef instantiates HSequence from 
    	    PCollection (ExternRef from ObjMgt);

end ObjMgt;
