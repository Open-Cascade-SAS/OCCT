-- Created on: 1993-01-20
-- Created by: Laurent PAINNOT
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MyLineTool from AppDef

uses MultiLine     from AppDef,
     Pnt           from gp,
     Pnt2d         from gp,
     Vec           from gp,
     Vec2d         from gp,
     Array1OfPnt   from TColgp,
     Array1OfPnt2d from TColgp,
     Array1OfVec   from TColgp,
     Array1OfVec2d from TColgp,
     Status        from Approx

is
    
    
    FirstPoint(myclass; ML: MultiLine) returns Integer;
    	---Purpose: Returns the first index of multipoints of the MultiLine.


    LastPoint(myclass; ML: MultiLine) returns Integer;
    	---Purpose: Returns the last index of multipoints of the MultiLine.



    NbP2d(myclass; ML: MultiLine) returns Integer;
    	---Purpose: Returns the number of 2d points of a MultiLine.


    NbP3d(myclass; ML: MultiLine) returns Integer;
    	---Purpose: Returns the number of 3d points of a MultiLine.


    Value(myclass; ML: MultiLine; MPointIndex: Integer; 
          tabPt: out Array1OfPnt);
    	---Purpose: returns the 3d points of the multipoint <MPointIndex>
    	--          when only 3d points exist.


    Value(myclass; ML: MultiLine; MPointIndex: Integer; 
          tabPt2d: out Array1OfPnt2d);
    	---Purpose: returns the 2d points of the multipoint <MPointIndex>
    	--          when only 2d points exist.


    Value(myclass; ML: MultiLine; MPointIndex: Integer; 
          tabPt: out Array1OfPnt; tabPt2d: out Array1OfPnt2d);
    	---Purpose: returns the 3d and 2d points of the multipoint 
    	--          <MPointIndex>.


    Tangency(myclass; ML: MultiLine; MPointIndex: Integer; 
             tabV: out Array1OfVec) returns Boolean;
    	---Purpose: returns the 3d points of the multipoint <MPointIndex>
    	--          when only 3d points exist.


    Tangency(myclass; ML: MultiLine; MPointIndex: Integer; 
          tabV2d: out Array1OfVec2d) returns Boolean;
    	---Purpose: returns the 2d tangency points of the multipoint 
    	--          <MPointIndex> only when 2d points exist.


    Tangency(myclass; ML: MultiLine; MPointIndex: Integer; 
             tabV: out Array1OfVec; tabV2d: out Array1OfVec2d)
    returns Boolean;
    	---Purpose: returns the 3d and 2d points of the multipoint 
    	--          <MPointIndex>.


    Curvature(myclass; ML: MultiLine; MPointIndex: Integer; 
             tabV: out Array1OfVec) returns Boolean;
    	---Purpose: returns the 3d curvatures of the multipoint <MPointIndex>
    	--          when only 3d points exist.


    Curvature(myclass; ML: MultiLine; MPointIndex: Integer; 
          tabV2d: out Array1OfVec2d) returns Boolean;
    	---Purpose: returns the 2d curvatures of the multipoint 
    	--          <MPointIndex> only when 2d points exist.


    Curvature(myclass; ML: MultiLine; MPointIndex: Integer; 
             tabV: out Array1OfVec; tabV2d: out Array1OfVec2d)
    returns Boolean;
    	---Purpose: returns the 3d and 2d curvatures of the multipoint 
    	--          <MPointIndex>.



    WhatStatus(myclass; ML: MultiLine; I1, I2: Integer) 
    returns Status from Approx;
    	---Purpose:  returns NoPointsAdded
    
    MakeMLBetween(myclass; ML: MultiLine; I1, I2: Integer;
                  NbPMin: Integer) 
    returns MultiLine;
    	---Purpose: Is never called in the algorithms.
    	--          Nothing is done.
    	---C++: return &


end MyLineTool;
