-- Created on: 1991-03-05
-- Created by: Philippe DAUTRY
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package GccAna 

    ---Purpose : This package provides an implementation of analytics 
    --         algorithms (using only non persistant entities) used 
    --         to create 2d lines or circles with geometric constraints.

uses Standard,
     StdFail,
     gp,
     TColStd,
     TColgp,
     GccInt,
     GccEnt
     

is

    -- Exceptions :

exception NoSolution inherits Failure from Standard;

class Lin2dTanPar;
    ---Purpose : Creates a 2d line TANgent to an 2d entity and PARallel 
    --         to another 2d line.

class Lin2dTanPer;
    ---Purpose : Creates a 2d line TANgent to an 2d entity and PERpendicular
    --         to another 2d entity.

class Lin2dTanObl;
    ---Purpose : Creates a 2d line TANgent to an 2d entity and OBLic 
    --         to another 2d entity.

class Lin2d2Tan;
    ---Purpose : Creates a 2d line TANgent to 2 2d entities.

class Lin2dBisec;
    ---Purpose : Creates a 2d line BISECting line of 2 2d lines.

class Circ2dTanCen;
    ---Purpose : Creates a 2d circle TANgent to a 2d entity and CENtered
    --         on a 2d point.

class Circ2d3Tan;
    ---Purpose : Creates a 2d circle TANgent to 3 2d entities.

class Circ2d2TanRad;
    ---Purpose : Creates a 2d circle TANgent to 2 2d entities with 
    --         the given RADius.

class Circ2d2TanOn;
    ---Purpose : Creates a 2d circle TANgent to a 2d entity and centered 
    --         ON a 2d entity (not a point).

class Circ2dTanOnRad;
    ---Purpose : Creates a 2d circle TANgent to a 2d entity and centered 
    --         ON a 2d entity (not a point) with the given radius.

class Pnt2dBisec;
    ---Purpose : Creates a 2d line BISECting line of 2 2d points.

class Circ2dBisec;
    ---Purpose : Creates a 2d line BISECting line of 2 2d circles.

class CircLin2dBisec;
    ---Purpose : Creates a 2d line BISECting line of a 2d circle 
    --         and a 2d line.

class CircPnt2dBisec;
    ---Purpose : Creates a 2d line BISECting line of a 2d circle 
    --         and a 2d point.

class LinPnt2dBisec;
    ---Purpose : Creates a 2d line BISECting line of a 2d line 
    --         and a 2d point.

end GccAna;
