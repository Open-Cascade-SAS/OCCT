-- Created on: 1992-01-24
-- Created by: Remi LEQUETTE
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package TopAbs 
	---Purpose: This package gives resources for Topology oriented
	--          applications such as : Topological Data Structure,
	--          Topological Algorithms.
	--          
	--          It contains :
	--          
	--            * The ShapeEnum   enumeration  to  describe  the
	--            differents topological shapes.
	--            
	--            * The  Orientation  enumeration to  describe the
	--            orientation of a topological shape.
	--            
	--            * The  State    enumeration  to  describes  the
	--            position of a point relative to a Shape.
	--            
	--            * Methods to manage the enumerations.

    ---Level : Public.
    --  All methods of all  classes will be public.

is

    enumeration ShapeEnum is 
    ---Purpose: Identifies various topological shapes. This
    -- enumeration allows you to use dynamic typing of shapes.
    -- The values are listed in order of complexity, from the
    -- most complex to the most simple i.e.
    -- COMPOUND > COMPSOLID > SOLID > .... > VERTEX > SHAPE.
    --  Any shape can contain simpler shapes in its definition.
    -- Abstract topological data structure describes a basic
    -- entity, the shape (present in this enumeration as the
    -- SHAPE value), which can be divided into the following
    -- component topologies:
    -- - COMPOUND: A group of any of the shapes below.
    -- - COMPSOLID: A set of solids connected by their
    --   faces. This expands the notions of WIRE and SHELL to solids.
    -- - SOLID: A part of 3D space bounded by shells.
    -- - SHELL: A set of faces connected by some of the
    --   edges of their wire boundaries. A shell can be open or closed.
    -- - FACE: Part of a plane (in 2D geometry) or a surface
    --   (in 3D geometry) bounded by a closed wire. Its
    --   geometry is constrained (trimmed) by contours.
    -- - WIRE: A sequence of edges connected by their
    --  vertices. It can be open or closed depending on
    --  whether the edges are linked or not.
    -- - EDGE: A single dimensional shape corresponding
    --   to a curve, and bound by a vertex at each extremity.
    -- - VERTEX: A zero-dimensional shape corresponding to a point in geometry.
        COMPOUND,
        COMPSOLID,
        SOLID,
        SHELL,
        FACE,
    	WIRE,
        EDGE,
        VERTEX,
        SHAPE

    end ShapeEnum;

    enumeration Orientation is 
    ---Purpose: Identifies the orientation of a topological shape.
    -- Orientation can represent a relation between two
    -- entities, or it can apply to a shape in its own right.
    -- When used to describe a relation between two
    -- shapes, orientation allows you to use the underlying
    -- entity in either direction. For example on a curve
    -- which is oriented FORWARD (say from left to right)
    -- you can have both a FORWARD and a REVERSED
    -- edge. The FORWARD edge will be oriented from
    -- left to right, and the REVERSED edge from right to
    -- left. In this way, you share the underlying entity. In
    -- other words, two faces of a cube can share an
    -- edge, and can also be used to build compound shapes.
    -- For each case in which an element is used as the
    -- boundary of a geometric domain of a higher
    -- dimension, this element defines two local regions of
    -- which one is arbitrarily considered as the default
    -- region. A change in orientation implies a switch of
    -- default region. This allows you to apply changes of
    -- orientation to the shape as a whole.
        FORWARD,
        REVERSED,
        INTERNAL,
        EXTERNAL

    end Orientation;

    enumeration State is 
    ---Purpose: Identifies the position of a vertex or a set of
    -- vertices relative to a region of a shape.   
    -- The figure shown above illustrates the states of
    -- vertices found in various parts of the edge relative
    -- to the face which it intersects.
	IN,
	OUT,
	ON,
	UNKNOWN

    end State;
    
   
    Compose(Or1  : Orientation from TopAbs;
            Or2  : Orientation from TopAbs)
    returns Orientation from TopAbs;
    ---Purpose: Compose  the Orientation    <Or1>  and  <Or2>.    This
    --          composition is not symmetric (if  you switch <Or1> and
    --          <Or2> the result  is different). It assumes that <Or1>
    --          is the Orientation of a Shape S1 containing a Shape S2
    --          of Orientation   Or2.  The result    is the  cumulated
    --          orientation of S2 in S1.  The composition law is :
    --          
    --             \ Or2     FORWARD  REVERSED INTERNAL EXTERNAL
    --           Or1       -------------------------------------
    --           FORWARD   | FORWARD  REVERSED INTERNAL EXTERNAL
    --                     |
    --           REVERSED  | REVERSED FORWARD  INTERNAL EXTERNAL
    --                     |
    --           INTERNAL  | INTERNAL INTERNAL INTERNAL INTERNAL
    --                     |
    --           EXTERNAL  | EXTERNAL EXTERNAL EXTERNAL EXTERNAL
    --     Note: The top corner in the table is the most important
    -- for the purposes of Open CASCADE topology and shape sharing.      

    Reverse(Or : Orientation from TopAbs)
    returns Orientation from TopAbs;
    ---Purpose: xchanges the interior/exterior status of the two
    -- sides. This is what happens when the sense of
    -- direction is reversed. The following rules apply:
    --          
    --          FORWARD          REVERSED
    --          REVERSED         FORWARD
    --          INTERNAL         INTERNAL
    --          EXTERNAL         EXTERNAL
    --          
    --          Reverse exchange the material sides.
    --          

    Complement(Or : Orientation from TopAbs)
    returns Orientation from TopAbs;
    ---Purpose: Reverses the interior/exterior status of each side of
    -- the object. So, to take the complement of an object
    -- means to reverse the interior/exterior status of its
    -- boundary, i.e. inside becomes outside.
    -- The method returns the complementary orientation,
    -- following the rules in the table below:
    --          FORWARD          REVERSED
    --          REVERSED         FORWARD
    --          INTERNAL         EXTERNAL
    --          EXTERNAL         INTERNAL
    --          
    --          Complement  complements   the  material  side.  Inside
    --          becomes outside.
    --          

    Print(SE  : ShapeEnum  from TopAbs; S  : in out OStream) returns OStream;
    ---Purpose: Prints the name  of Shape  <SEq>  as  a String  on the
    --          Stream <S> and returns <S>.
    --          
    ---C++: return &

    Print(Or  : Orientation  from TopAbs; S  : in out OStream) returns OStream;
    ---Purpose: Prints the name of the Orientation <Or> as a String on
    --          the Stream <S> and returns <S>.
    --          
    ---C++: return &

    Print(St  : State  from TopAbs; S  : in out OStream) returns OStream;
    ---Purpose: Prints the name of the State <St> as a String on
    --          the Stream <S> and returns <S>.
    --          
    ---C++: return &

end TopAbs;
