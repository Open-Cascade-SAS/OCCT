-- Created on: 1997-03-04
-- Created by: Jean-Pierre COMBE
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class OffsetDimension from AIS inherits Relation from AIS

	---Purpose: A framework to display dimensions of offsets.
    	-- The relation between the offset and the basis shape
    	-- is indicated. This relation is displayed with arrows and
    	-- text. The text gives the dsitance between the offset
    	-- and the basis shape.
        
uses
     Shape                 from TopoDS,
     Presentation          from Prs3d,
     Projector             from Prs3d,
    Transformation        from Geom,
     PresentationManager3d from PrsMgr,
     PresentationManager2d from PrsMgr,
     Selection             from SelectMgr,
     GraphicObject         from Graphic2d,
     Dir                   from gp,
     Pnt                   from gp,
     Trsf                  from gp,
     KindOfDimension       from AIS,
     ExtendedString        from TCollection     
     
is
    Create (FistShape, SecondShape : Shape          from TopoDS;
	    aVal                   : Real           from Standard;
	    aText                  : ExtendedString from TCollection)
    returns mutable OffsetDimension from AIS;
    	---Purpose: Constructs the offset display object defined by the
    	-- first shape aFShape, the second shape aSShape, the
    	-- dimension aVal, and the text aText.    

    Compute(me            : mutable;
    	    aPresentationManager: PresentationManager3d from PrsMgr;
    	    aPresentation : mutable Presentation from Prs3d;
    	    aMode         : Integer from Standard= 0) 
    is redefined private;

    Compute(me:mutable;
    	        aProjector: Projector from Prs3d;
                aPresentation: mutable Presentation from Prs3d)
    is redefined static private;     

    Compute(me:mutable;
    	    aPresentationManager: PresentationManager2d from PrsMgr;
            aPresentation: mutable GraphicObject from Graphic2d;
            aMode: Integer from Standard = 0)
    is redefined static private;	
    
    Compute(me            : mutable;
    	    aProjector    : Projector from Prs3d;
    	    aTrsf         : Transformation from Geom;
	    aPresentation : mutable Presentation from Prs3d)
    is redefined;
    	---Purpose: computes the presentation according to a point of view
    	--          given by <aProjector>. 
    	--          To be Used when the associated degenerated Presentations 
    	--          have been transformed by <aTrsf> which is not a Pure
    	--          Translation. The HLR Prs can't be deducted automatically
    	--          WARNING :<aTrsf> must be applied
    	--           to the object to display before computation  !!!

-- Methods from SelectableObject

    ComputeSelection(me         : mutable;
    	    	     aSelection : mutable Selection from SelectMgr;
    	    	     aMode      : Integer from Standard)
    is redefined private;

    KindOfDimension(me)
   	---Purpose:
    	-- Indicates that the dimension we are concerned with is an offset.
        ---C++: inline
    returns KindOfDimension from AIS 
    is redefined;
    
    IsMovable(me) 
       ---C++: inline       
       ---Purpose: Returns true if the offset datum is movable. 
            returns Boolean from Standard 
    is redefined;    
    
    SetRelativePos (me:mutable; aTrsf: Trsf from gp);
        ---C++: inline
    	---Purpose: Sets a transformation aTrsf for presentation and
    	-- selection to a relative position.

    ComputeTwoFacesOffset(me: mutable;
    	    	    	  aPresentation : mutable Presentation from Prs3d;
    	    	    	  aTrsf         : Trsf from gp)
    is private;
    
    ComputeTwoAxesOffset(me: mutable;
    	    	    	  aPresentation : mutable Presentation from Prs3d;
    	    	    	  aTrsf         : Trsf from gp)
    is private;

    ComputeAxeFaceOffset(me: mutable;
    	    	  	  aPresentation : mutable Presentation from Prs3d;
    	    	    	  aTrsf         : Trsf from gp)
    is private;

fields

    myFAttach     : Pnt  from gp;
    mySAttach     : Pnt  from gp;
    myDirAttach   : Dir  from gp;
    myDirAttach2  : Dir  from gp;
    myRelativePos : Trsf from gp;

end OffsetDimension;
