-- Created on: 1992-12-02
-- Created by: Isabelle GRIGNON
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class SelGProps from GProp inherits GProps

    	    ---Purpose: 
    	    --          Computes the global properties of an elementary 
    	    --          surface (surface of the gp package)

uses  Cylinder from gp,
      Cone     from gp,
      Pnt      from gp,
      Sphere   from gp,
      Torus    from gp

is

  Create returns SelGProps;

  Create (S : Cylinder; Alpha1, Alpha2, Z1, Z2 : Real; SLocation : Pnt)   
     returns SelGProps;


  Create (S : Cone; Alpha1, Alpha2, Z1, Z2 : Real; SLocation : Pnt)   
     returns SelGProps;


  Create (S : Sphere from gp; Teta1, Teta2, Alpha1, Alpha2 : Real;
          SLocation : Pnt)   
     returns SelGProps;


  Create (S : Torus from gp; Teta1, Teta2, Alpha1, Alpha2 : Real;
          SLocation : Pnt)   
     returns SelGProps;

  SetLocation(me : in out ;SLocation :Pnt);

  Perform(me : in out;S : Cylinder; Alpha1, Alpha2, Z1, Z2 : Real);

  Perform(me : in out;S : Cone; Alpha1, Alpha2, Z1, Z2 : Real);

  Perform(me : in out;S : Sphere; Teta1, Teta2, Alpha1, Alpha2 : Real);

  Perform(me : in out;S : Torus; Teta1, Teta2, Alpha1, Alpha2 : Real);

end SelGProps;
