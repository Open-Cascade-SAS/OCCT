-- Created on: 1993-08-24
-- Created by: GG
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class TypeMap from Xw inherits Transient

	---Version: 0.0

	---Purpose: This class defines a TypeMap object.

	---Keywords:
	---Warning:
	---References:

uses

	TypeMap		from Aspect,
	TypeMapEntry	from Aspect,
	LineStyle 	from Aspect

raises

	TypeMapDefinitionError	from Aspect,
	BadAccess		from Aspect

is

	Create
	returns mutable TypeMap from Xw
	is protected ;
	---Level: Internal

	Create ( Connexion : CString from Standard ) 
	returns mutable TypeMap from Xw 
	---Level: Public
	---Purpose: Creates a TypeMap with unallocated TypeMapEntry.
	--  Warning: Raises if TypeMap creation failed according
	--	    to the supported hardware
	raises TypeMapDefinitionError from Aspect ;

	SetEntry ( me : mutable ; 
		   Entry : TypeMapEntry from Aspect )
	---Level: Public
	---Purpose: Modifies an entry already defined or Add the Entry
	--	    in the type map <me> if it don't exist.
	--  Warning: Raises if TypeMap size is exceeded,
	--	    or TypeMap is not defined properly,
	--	    or TypeMapEntry Index is out of range according
	--	    to the supported hardware
	raises BadAccess from Aspect is virtual;

	SetEntries ( me : mutable ; 
		     Typemap : TypeMap from Aspect ) 
	---Level: Public
	---Purpose: Modifies all entries from a new Typemap
	--  Warning: Raises if TypeMap size is exceeded,
	--	    or TypeMap is not defined properly,
	--	    or One of new TypeMapEntry Index is out of range according
	--	    to the supported hardware
	raises BadAccess from Aspect is virtual;

	Destroy ( me : mutable ) is virtual;
	---Level: Public
	---Purpose: Destroies the Typemap
	---C++: alias ~

	----------------------------
	-- Category: Inquire methods
	----------------------------

	FreeTypes ( me )
	returns Integer from Standard 
	---Level: Public
	---Purpose: Returns the Number of Free Types in the Typemap
	--	    depending of the HardWare
	--  Warning: Raises if TypeMap is not defined properly
	raises BadAccess from Aspect is static;

	ExtendedTypeMap ( me )
	returns Address from Standard
	is static protected ;
	---Level: Internal
	---Purpose: Returns extended data typemap structure pointer.
	---Category: Inquire methods


fields

	MyExtendedDisplay	: Address from Standard ;
	MyExtendedTypeMap 	: Address from Standard ;

friends

	class GraphicDevice from Xw

end TypeMap ;
