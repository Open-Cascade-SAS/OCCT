-- Created on: 1991-05-27
-- Created by: Laurent PAINNOT
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class IntegerRandom from math
   ---Purpose:
   -- This class implements an integer random number generator.

is

   Create(Lower, Upper: Integer)
   ---Purpose:
   -- creates a Integer random generator between the values Lower and Upper.
    
   returns IntegerRandom;
   
    
   Reset(me:in out)
    	---Purpose: reinitializes the random generator

   is static;

   Next(me: in out)
    ---Purpose: returns the next random number.

   returns Integer
   is static;
   
fields

Low:    Integer;
Up:     Integer;
Dummy:  Integer;

end IntegerRandom;
