-- Created on: 1996-12-05
-- Created by: Philippe MANGIN
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Tensor from  GeomFill 

	---Purpose: used to store the "gradient of gradient"

uses
    Array1OfReal from TColStd,
    Vector from math,
    Matrix from math

raises DimensionError from Standard, 
       RangeError from Standard 

is
    Create(NbRow, NbCol, NbMat : Integer) 
    returns Tensor;
 
    Init(me : in out; InitialValue: Real)
	   ---Purpose:Initialize all the elements of a Tensor to InitialValue.
    is static;
 
    Value(me; Row, Col, Mat: Integer)
    	---Purpose: accesses (in read or write mode) the value of index <Row>,
    	--          <Col> and <Mat> of a Tensor.
    	--          An exception is raised if <Row>, <Col> or <Mat> are not
    	--          in the correct range.
    	---C++: alias operator() 
    	---C++: return const & 
    	---C++: inline
    returns Real
    is static;
    
    ChangeValue(me : in out; Row, Col, Mat: Integer)
    	---Purpose: accesses (in read or write mode) the value of index <Row>,
    	--          <Col> and <Mat> of a Tensor.
    	--          An exception is raised if <Row>, <Col> or <Mat> are not
    	--          in the correct range.
    	---C++: alias operator() 
    	---C++: return & 
    	---C++: inline
    returns Real
    is static;

    Multiply(me; Right: Vector; Product:out Matrix)
    raises DimensionError
    is static;
    

fields
    Tab     : Array1OfReal;
    nbrow   : Integer;
    nbcol   : Integer;
    nbmat   : Integer;
    nbmtcl  : Integer;
end ;
