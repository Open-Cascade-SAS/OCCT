-- Created on: 1994-04-18
-- Created by: Modelistation
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Marker2D from Draw inherits Drawable2D from Draw

	---Purpose: 

uses
    Pnt2d from gp,
    Color from Draw,
    MarkerShape from Draw,
    Display from Draw

is
    Create(P : Pnt2d from gp; T : MarkerShape from Draw; C : Color from Draw; 
    	Size : Integer = 5) returns mutable Marker2D from Draw;
	
    Create(P : Pnt2d from gp; T : MarkerShape from Draw; C : Color from Draw; 
    	RSize : Real) returns mutable Marker2D from Draw;
    
    ChangePos(me : mutable) returns Pnt2d from gp;
    ---C++: return &
    ---Purpose: myPos field

    DrawOn(me; dis : in out Display from Draw);

    PickReject(me; X,Y,Prec : Real) returns Boolean
	---Purpose: Returs always false
    is redefined;
    

fields
    myPos : Pnt2d from gp;
    myCol : Color from Draw;
    myTyp : MarkerShape from Draw;
    mySiz : Integer;

end Marker2D;
