-- File:	QANewBRepNaming_Cylinder.cdl
-- Created:	Fri Aug 22 11:16:27 1997
-- Author:	VAUTHIER Jean-Claude
---Copyright:	 Open CASCADE 2003


class Cylinder from QANewBRepNaming inherits TopNaming from QANewBRepNaming

    ---Purpose: To load the Cylinder results

uses 
 
    MakeCylinder from BRepPrimAPI,
    Label        from TDF,
    TypeOfPrimitive3D from QANewBRepNaming

is

    Create returns Cylinder from QANewBRepNaming;

    Create(ResultLabel : Label from TDF) 
    returns Cylinder from QANewBRepNaming; 
     
    Init(me : in out; ResultLabel : Label from TDF);


    Load (me; mkCylinder : in out MakeCylinder from BRepPrimAPI; Type : TypeOfPrimitive3D from QANewBRepNaming);

    Bottom (me)
    ---Purpose: Returns the label of the bottom
    --          face of the cylinder.
    returns Label from TDF;

    Top (me)
    ---Purpose: Returns the label of the top
    --          face of the cylinder.
    returns Label from TDF;

    Lateral (me)
    ---Purpose: Returns the label of the lateral
    --          face of the cylinder.
    returns Label from TDF;

    StartSide (me)
    ---Purpose: Returns the label of the first
    --          side of the cylinder
    returns Label from TDF;
        
    EndSide (me)
    ---Purpose: Returns the label of the second
    --          side of the cylinder.
    returns Label from TDF;


end Cylinder;



