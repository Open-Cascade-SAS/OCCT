-- File:        AutoDesignDateAndPersonAssignment.cdl
-- Created:     Mon Dec  4 12:02:23 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWAutoDesignDateAndPersonAssignment from RWStepAP214

	---Purpose : Read & Write Module for AutoDesignDateAndPersonAssignment

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     AutoDesignDateAndPersonAssignment from StepAP214,
     EntityIterator from Interface

is

	Create returns RWAutoDesignDateAndPersonAssignment;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable AutoDesignDateAndPersonAssignment from StepAP214);

	WriteStep (me; SW : in out StepWriter; ent : AutoDesignDateAndPersonAssignment from StepAP214);

	Share(me; ent : AutoDesignDateAndPersonAssignment from StepAP214; iter : in out EntityIterator);

end RWAutoDesignDateAndPersonAssignment;
