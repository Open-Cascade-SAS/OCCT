-- Created on: 1993-04-22
-- Created by: Laurent PAINNOT
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



deferred generic class TheLineTool from AppCont(MLine as any)

    ---Purpose: Template for desribing a continuous MultiLine.
    --          The Vectors returned by the methods Tangency are
    --          the derivative values.

uses
     Pnt           from gp,
     Pnt2d         from gp,
     Vec           from gp,
     Vec2d         from gp,
     Array1OfPnt   from TColgp,
     Array1OfPnt2d from TColgp,
     Array1OfVec   from TColgp,
     Array1OfVec2d from TColgp

is
    
    FirstParameter(myclass; ML: MLine) returns Real;
    	---Purpose: returns the first parameter of the Line.

    LastParameter(myclass; ML: MLine) returns Real;
    	---Purpose: returns the last parameter of the Line.

    NbP2d(myclass; ML: MLine) returns Integer;
    	---Purpose: Returns the number of 2d points of a MLine.


    NbP3d(myclass; ML: MLine) returns Integer;
    	---Purpose: Returns the number of 3d points of a MLine.


    Value(myclass; ML: MLine; U: Real; tabPt: out Array1OfPnt);
    	---Purpose: returns the 3d points of the multipoint <MPointIndex>
    	--          when only 3d points exist.


    Value(myclass; ML: MLine; U: Real; tabPt2d: out Array1OfPnt2d);
    	---Purpose: returns the 2d points of the multipoint <MPointIndex>
    	--          when only 2d points exist.


    Value(myclass; ML: MLine; U: Real; 
          tabPt: out Array1OfPnt; tabPt2d: out Array1OfPnt2d);
    	---Purpose: returns the 3d and 2d points of the multipoint 
    	--          <MPointIndex>.


    D1(myclass; ML: MLine; U: Real; tabV: out Array1OfVec)
    returns Boolean;
    	---Purpose: returns the 3d derivative values of the multipoint 
    	--          <MPointIndex> when only 3d points exist.


    D1(myclass; ML: MLine; U: Real; tabV2d: out Array1OfVec2d)
    returns Boolean;
    	---Purpose: returns the 2d derivative values of the multipoint 
    	--          <MPointIndex> only when 2d points exist.


    D1(myclass; ML: MLine; U: Real; 
             tabV: out Array1OfVec; tabV2d: out Array1OfVec2d)
    returns Boolean;
    	---Purpose: returns the 3d and 2d derivative values of the multipoint 
    	--          <MPointIndex>.


end TheLineTool;    
    
