-- File:	StepAP214_ExternallyDefinedGeneralProperty.cdl
-- Created:	Wed May 10 15:09:07 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class ExternallyDefinedGeneralProperty from StepAP214
inherits GeneralProperty from StepBasic

    ---Purpose: Representation of STEP entity ExternallyDefinedGeneralProperty

uses
    HAsciiString from TCollection,
    SourceItem from StepBasic,
    ExternalSource from StepBasic,
    ExternallyDefinedItem from StepBasic

is
    Create returns ExternallyDefinedGeneralProperty from StepAP214;
	---Purpose: Empty constructor

    Init (me: mutable; aGeneralProperty_Id: HAsciiString from TCollection;
                       aGeneralProperty_Name: HAsciiString from TCollection;
                       hasGeneralProperty_Description: Boolean;
                       aGeneralProperty_Description: HAsciiString from TCollection;
                       aExternallyDefinedItem_ItemId: SourceItem from StepBasic;
                       aExternallyDefinedItem_Source: ExternalSource from StepBasic);
	---Purpose: Initialize all fields (own and inherited)

    ExternallyDefinedItem (me) returns ExternallyDefinedItem from StepBasic;
	---Purpose: Returns data for supertype ExternallyDefinedItem
    SetExternallyDefinedItem (me: mutable; ExternallyDefinedItem: ExternallyDefinedItem from StepBasic);
	---Purpose: Set data for supertype ExternallyDefinedItem

fields
    theExternallyDefinedItem: ExternallyDefinedItem from StepBasic; -- supertype

end ExternallyDefinedGeneralProperty;
