-- Created on: 2008-05-04
-- Created by: Vladislav ROMASHKO
-- Copyright (c) 2008-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


package Voxel

    ---Purpose: Data structuire and visualization engine for voxel modeling.

uses

    IntCurvesFace,
    TCollection,
    SelectMgr,
    Quantity,
    TopTools,
    TColStd,
    TColgp,
    TopoDS,
    PrsMgr,
    Prs3d,
    Poly,
    V3d,
    AIS,
    Bnd,
    gp

is

    enumeration VoxelDisplayMode is
    	VDM_POINTS,
	VDM_NEARESTPOINTS,
	VDM_BOXES,
	VDM_NEARESTBOXES
    end VoxelDisplayMode;

    enumeration VoxelFileFormat is
    	VFF_ASCII,
	VFF_BINARY
    end VoxelFileFormat;

    -- A base class for all voxels data structures.
    class DS;

	    -- A voxel model keeping a boolean flag for each voxel (1 || 0).
	    class BoolDS;
	    
	    	-- A voxel model keeping a boolean flag for each voxel 
	    	-- with an opportunity to split a voxel into 8 sub-voxels.
	    	class OctBoolDS;

    	    	    -- A voxel model keeping a boolean flag for each voxel 
	    	    -- with an opportunity to split a voxel into 8 sub-voxels
	    	    -- recursively.
    	    	    class ROctBoolDS;
		    	private class SplitData;

	    -- A voxel model keeping 4 bits of information for each voxel (16 colors).
	    class ColorDS;
	    
	    -- A voxel model keeping 4 bytes of information for each voxel (a floating-point value).
	    class FloatDS;


    -- A converter of a shape to voxel model.
    --class Converter;
    
    	-- An internal class searching intersections between a line and a shape.
    	--class ShapeIntersector;
    
    -- An alternative method of conversion of a shape into voxels.
    -- It is faster, but less precise.
    class FastConverter;
    
    --- Converts voxels into triangulation
    --class Triangulator;
    
    -- Interactive object of voxels
    class Prs;

    -- Boolean operations for voxels.
    class BooleanOperation;
    
    -- Collision detection
    class CollisionDetection;

    -- Selection of voxels in the viewer 3d
    class Selector;

    -- Ascii writer/reader of voxels
    class Writer;
    class Reader;
    

end Voxel;
