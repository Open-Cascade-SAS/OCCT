-- Created on: 2000-08-15
-- Created by: data exchange team
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package PXCAFDoc 

	---Purpose: This pakage is the persistent equivalent of
	--          XCAFDoc

uses
    Quantity,
    TopLoc,
    PTopLoc,
    PDF,
    PDataStd,
    gp,
    PCollection,
    PColStd
is
    class Location;
    class Color;
    class Volume;
    class Area;
    class Centroid;
    class ColorTool;
    class ShapeTool;
    class DocumentTool;
    class LayerTool;
    class GraphNode;
    class GraphNodeSequence instantiates HSequence from PCollection
    	(GraphNode from PXCAFDoc);
    class Datum;
    class DimTol;
    class DimTolTool;
    class Material;
    class MaterialTool;

end PXCAFDoc;
