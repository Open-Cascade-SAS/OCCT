--
-- File:	AlienImage_AidaAlienData.cdl
-- Created:	23/03/93
-- Author:	BBL
--
---Copyright:	Matravision 1993
--

class AidaAlienData from AlienImage inherits AlienImageData from AlienImage

	---Version: 0.0

	---Level: Public
	---Purpose: This class defines an Aida Alien image.


uses
	File 			from OSD,
	ColorImage 		from Image,
	PseudoColorImage 	from Image,
	ColorMap 		from Aspect,
	HArray2OfInteger 	from TColStd,
	DitheringMethod 	from Image,
	Image			from Image

raises
	OutOfRange 	from Standard,
	TypeMismatch 	from Standard

is
	Create returns mutable AidaAlienData from AlienImage ;

	Clear( me : in out mutable ) ;
	---Level: Public
	---Purpose: Frees memory allocated by AidaAlienData
	---C++: alias ~

	Read ( me : in out mutable ; afile : in out File from OSD )
	  returns Boolean from Standard ;
	---Level: Public
	  ---Purpose: Read content of a  AidaAlienData object from a file .
	  --          Returns True if file is a Aida file .

	Write( me : in immutable; afile : in out File from OSD )
	  returns Boolean from Standard ;
	---Level: Public
	  ---Purpose: Write content of a  AidaAlienData object to a file .

	ToImage( me : in  immutable) 
	  returns mutable Image from Image 
          raises TypeMismatch from Standard ;
	  ---Purpose : Converts a AidaAlienData object to a Image object.

	FromImage( me : in out mutable ; anImage : in Image from Image )
          raises TypeMismatch from Standard ;
	  ---Purpose : Converts a Image object to a AidaAlienData object.

	SetColorImageDitheringMethod( me : in out mutable ; 
				      aMethod : DitheringMethod from Image;
				      aColorMap : ColorMap from Aspect ) ;

	---Level: Public
	  ---Purpose: Set the ImageDitheringMethod and the ColorMap when
	  --          FromImage is called with a ColorImage .
	  --	      Aida BYTEMAPS file handle only PseudoColorImage .
	  --          Default value is DM_NearestColor,
	  --		ColorCubeColorMap( 40, 5,1, 8,6, 3,54 )


        AllocData( me : in out mutable ; DX,DY : in Integer from Standard ) 
		is private;
	---Level: Internal
	   ---Purpose : Allocate HArray2 to store Image data

    	Pixel   ( me : in immutable ;     X,Y : in Integer from Standard ) 
			returns Integer from Standard
    			raises OutOfRange from Standard is private ;
	---Level: Internal

    	SetPixel( me : in out mutable; X,Y   : in Integer from Standard ;
			Value : in Integer from Standard )
    			raises OutOfRange from Standard is private ;
	---Level: Internal

	FromPseudoColorImage( me      : in out mutable; 
			      anImage : in PseudoColorImage from Image )
		is private ;
	---Level: Internal
	  ---Purpose : convert a Image object to a AidaAlienData object.

	FromColorImage( me : in out mutable;
			anImage : in ColorImage from Image)
		is private ;
	---Level: Internal
	  ---Purpose : convert a Image object to a AidaAlienData object.

fields
	myDitheringMethod   : DitheringMethod from Image is protected ;

	myDitheringColorMap : ColorMap from Aspect  is protected ;

	myColors : ColorMap from Aspect  is protected ;
	myColorsIsDef : Boolean from Standard  is protected ;

			-- AidaColors definition
	myData	 : HArray2OfInteger from TColStd ;
	myDataIsDef : Boolean from Standard  is protected ;

end ;
 
