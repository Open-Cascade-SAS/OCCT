-- Created on: 1997-02-12
-- Created by: Alexander BRIVIN
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Transform from Vrml 

	---Purpose:  defines a Transform of VRML specifying transform
	---          properties.
    	--  This  node  defines  a  geometric  3D  transformation   consisting   of  (in  order) 
    	--  a  (possibly)  non-uniform  scale  about  an  arbitrary  point,  a  rotation  about 
    	--  an arbitrary point  and  axis  and  translation. 
    	--  By  default  : 
	--    myTranslation (0,0,0) 
	--    myRotation  (0,0,1,0)
	--    myScaleFactor (1,1,1)
	--    myScaleOrientation (0,0,1,0)
	--    myCenter (0,0,0)

uses
 
   Vec         from  gp, 
   SFRotation  from  Vrml

is
 
    Create returns  Transform from Vrml; 
 
    Create ( aTranslation      : Vec         from  gp; 
    	     aRotation         : SFRotation  from  Vrml; 
    	     aScaleFactor      : Vec         from  gp; 
    	     aScaleOrientation : SFRotation  from  Vrml; 
             aCenter           : Vec         from  gp )
    	returns  Transform from Vrml; 

    SetTranslation ( me : in out;  aTranslation : Vec  from  gp );
    Translation ( me )  returns Vec  from  gp;

    SetRotation ( me : in out;  aRotation : SFRotation  from  Vrml );
    Rotation ( me )  returns  SFRotation  from  Vrml;

    SetScaleFactor ( me : in out;  aScaleFactor : Vec  from  gp );
    ScaleFactor ( me )  returns Vec  from  gp;

    SetScaleOrientation ( me : in out;  aScaleOrientation : SFRotation  from  Vrml );
    ScaleOrientation ( me  )  returns  SFRotation  from  Vrml;

    SetCenter ( me : in out;  aCenter : Vec  from  gp );
    Center ( me )  returns Vec  from  gp;

    Print  ( me;  anOStream: in out OStream from Standard) returns OStream from Standard;
    ---C++:  return  & 

fields
 
    myTranslation      : Vec         from  gp;   -- Translation vector
    myRotation         : SFRotation  from  Vrml; -- Rotation
    myScaleFactor      : Vec         from  gp;   -- Scale factors
    myScaleOrientation : SFRotation  from  Vrml; -- Defines rotational space for scale
    myCenter           : Vec         from  gp;   -- Center point for scale and rotate

end Transform;
