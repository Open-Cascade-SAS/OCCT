-- Created on: 1993-03-03
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

private class ItemLocation from PTopLoc inherits Persistent

	---Purpose: Provides  support  for  the implementation  of the
	--          class Location.

uses
    Datum3D  from PTopLoc,
    Location from PTopLoc

is
    Create(D : Datum3D from PTopLoc; 
    	   P : Integer from Standard;
	   N : Location from PTopLoc) 
    returns mutable ItemLocation from  PTopLoc;
	---Level: Internal 
    
    Datum3D(me) returns Datum3D from PTopLoc
    is static;
	---Level: Internal 

    Power(me)   returns Integer from Standard
    is static;
	---Level: Internal 
    
    Next(me)    returns Location from PTopLoc
    is static;
	---Level: Internal 
    
fields
    myDatum : Datum3D  from PTopLoc;
    myPower : Integer  from Standard;
    myNext  : Location from PTopLoc;

end ItemLocation;
