-- Created on: 1993-04-07
-- Created by: Laurent BUCHARD
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package IntCurveSurface

    ---Purpose: This package provides algorithmes to intersect a Curve 
    --          and a Surface. 
    --  Level: Internal
    --
    -- All the methods of the classes of this package are Internal.
    -- except the methods of the classes <Intersection,
    --                                    IntersectionPoint,
    --                                    IntersectionSegment>
    --
     

uses Standard, TCollection, TColStd, TColgp, gp, 
     Bnd, Intf, IntAna,
     IntImp, IntSurf, 
     GeomAbs, StdFail ,
     Adaptor3d, Geom,
     math

is    

    --------------------------------------------------
    enumeration TransitionOnCurve is
        Tangent,In,Out;
    ---Purpose:
    --     
    --     
    --                    
    --         \ Uo     ^        \ U1     ^
    --          \       | n       \       | n
    -- Surf  ====\======|===   ====\======|=== 
    --            \     .           \     .
    --             \    .            \    .
    --          U1  \   .          Uo \   .
    -- 
    --        
    --           ( In )            ( Out ) 
    --
    --     
    --     
    --       \           /
    --        \         /
    --         \       /
    --          \     /
    -- Surf =====-----=====
    --                             
    --       ( Tangent ) 
    --    Crb and Surf are  C1 
    --------------------------------------------------
    deferred class Intersection;
    --------------------------------------------------    
    class IntersectionPoint;  
    --------------------------------------------------    
    class IntersectionSegment;
    --------------------------------------------------
    class SequenceOfPnt instantiates 
    	Sequence from TCollection(
	    IntersectionPoint from IntCurveSurface);
    --------------------------------------------------	    
    class SequenceOfSeg instantiates 
    	Sequence from TCollection(
	    IntersectionSegment from IntCurveSurface);
    --------------------------------------------------    
    generic class HCurveTool;
    --------------------------------------------------
    generic class Polygon;
    --------------------------------------------------
    generic class Polyhedron;
    --------------------------------------------------
    generic class PolygonTool;
    --------------------------------------------------
    generic class PolyhedronTool;
    --------------------------------------------------    
    generic class QuadricCurveFunc;
    --------------------------------------------------   
    generic class QuadricCurveExactInter,
                  TheQuadCurvFunc;
    --------------------------------------------------
    generic class Inter, 
                  ThePolygon,
                  ThePolygonTool,
                  ThePolyhedron,
                  ThePolyhedronTool,
                  TheInterference,
		  TheCSFunction,
                  TheExactInter,
                  TheQuadCurvExactInter;
	
    -------------------------------------------------	
    
    --class HCurveTool instantiates 
    --	CurveTool from IntCurveSurface
    --        (HCurve     from Adaptor3d); 

    --class HInter instantiates 
    --    Inter from IntCurveSurface (
    --        HCurve        from Adaptor3d, 
    --        HCurveTool    from IntCurveSurface,
    --        HSurface      from Adaptor3d, 
    --        HSurfaceTool  from IntCurveSurface);


    class TheHCurveTool instantiates 
    	HCurveTool from IntCurveSurface (
	    HCurve from Adaptor3d);

    class HInter instantiates 
        Inter from IntCurveSurface (
            HCurve        from Adaptor3d,
            TheHCurveTool from IntCurveSurface,
            HSurface      from Adaptor3d,
            HSurfaceTool  from Adaptor3d);

end IntCurveSurface;
