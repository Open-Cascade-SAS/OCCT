-- Created on: 1997-05-13
-- Created by: Alexander BRIVIN
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class WFRestrictedFace from VrmlConverter 


    	---Purpose: WFRestrictedFace -     computes     the  wireframe
    	--          presentation  of faces  with   restrictions by  
    	--          displaying   a  given  number    of  U   and/or  V
    	--          isoparametric  curves,  converts this  one into VRML
    	--          objects  and writes  (adds)  into anOStream.
    	--          All requested  properties  of the representation
    	--          are specify in  aDrawer.
    	--          This kind of the presentation is converted into
    	--          IndexedLineSet ( VRML ).

        --          The isoparametric curves are drawn with a fixed
        --          number of points. 

uses
 
    HSurface     from BRepAdaptor,
    Drawer       from VrmlConverter

is
 
    Add(myclass; anOStream: in out OStream from Standard; 
        	 aFace: HSurface from BRepAdaptor;
    	    	 aDrawer: Drawer from VrmlConverter);
		 
    AddUIso(myclass; anOStream: in out OStream from Standard; 
        	     aFace: HSurface from BRepAdaptor;
    	    	     aDrawer: Drawer from VrmlConverter);
		 
    AddVIso(myclass; anOStream: in out OStream from Standard; 
        	     aFace: HSurface from BRepAdaptor;
    	    	     aDrawer: Drawer from VrmlConverter);

    Add(myclass;  anOStream: in out OStream from Standard; 
    	          aFace: HSurface from BRepAdaptor;
		  DrawUIso, DrawVIso: Boolean from Standard;
		  NBUiso,NBViso: Integer from Standard;
		  aDrawer: Drawer from VrmlConverter);
		   
end WFRestrictedFace;
