-- Created on: 2003-12-17
-- Created by: Alexander SOLOVYOV
-- Copyright (c) 2003-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Tool from MeshVS

	---Purpose: This class provides auxiliary methods to create differents aspects

uses
  Boolean from Standard,

  Drawer from MeshVS,

  AspectFillArea3d from Graphic3d,
  AspectLine3d     from Graphic3d,
  AspectMarker3d   from Graphic3d,
  AspectText3d     from Graphic3d,
  MaterialAspect   from Graphic3d,

  Array1OfReal     from TColStd,

  Vec              from gp,
  Dir              from gp

is
  CreateAspectFillArea3d ( myclass; theDr : Drawer; UseDefaults : Boolean = Standard_True ) returns AspectFillArea3d from Graphic3d;
	---Purpose: Creates fill area aspect with values from Drawer according to keys from DrawerAttribute

  CreateAspectFillArea3d ( myclass; theDr : Drawer; Mat : MaterialAspect; UseDefaults : Boolean = Standard_True ) returns AspectFillArea3d from Graphic3d;
	---Purpose: Creates fill aspect with values from Drawer according to keys from DrawerAttribute
        -- and specific material aspect

  CreateAspectLine3d     ( myclass; theDr : Drawer; UseDefaults : Boolean = Standard_True ) returns AspectLine3d from Graphic3d;
	---Purpose: Creates line aspect with values from Drawer according to keys from DrawerAttribute

  CreateAspectMarker3d   ( myclass; theDr : Drawer; UseDefaults : Boolean = Standard_True ) returns AspectMarker3d from Graphic3d;
	---Purpose: Creates marker aspect with values from Drawer according to keys from DrawerAttribute

  CreateAspectText3d     ( myclass; theDr : Drawer; UseDefaults : Boolean = Standard_True ) returns AspectText3d from Graphic3d;
	---Purpose: Creates text aspect with values from Drawer according to keys from DrawerAttribute

  GetNormal( myclass; Nodes : Array1OfReal from TColStd;
                      Norm  : out Vec from gp ) returns Boolean;
	---Purpose: Get one of normals to polygon described by these points.
        --          If the polygon isn't planar, function returns false

  GetAverageNormal( myclass; Nodes : Array1OfReal from TColStd;
                      Norm  : out Vec from gp ) returns Boolean;
	---Purpose: Get an average of normals to non-planar polygon described by these points or compute
        --          normal of planar polygon. If the polygon isn't planar, function returns false

end Tool;
