-- Created on: 1995-04-24
-- Created by: Bruno DUMORTIER
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

private class TrimEdgeTool from BRepFill 

	---Purpose: 

uses

    Bisec         from Bisector,
    Edge          from TopoDS,
    Pnt2d         from gp,
    Curve         from Geom2d,
    Geometry      from Geom2d,	
    SequenceOfPnt from TColgp,
    Curve         from Geom2dAdaptor

is
    Create
    returns TrimEdgeTool from BRepFill;
    
    Create( Bisec   : Bisec    from Bisector;
    	    S1, S2  : Geometry from Geom2d;
    	    Offset  : Real     from Standard)
    returns TrimEdgeTool from BRepFill;
    
    IntersectWith( me : in out;
    	    	   Edge1 , Edge2 :        Edge          from TopoDS;
		   Params        : in out SequenceOfPnt from TColgp)
    is static;

    AddOrConfuse ( me ;
    		   Start         :        Boolean       from Standard;
		   Edge1 , Edge2 :        Edge          from TopoDS;
		   Params  : in out SequenceOfPnt from TColgp)
    is static;		  


    IsInside( me; P : Pnt2d from gp)
    returns Boolean from Standard
    is static;
	      
    	    
		       
fields
    isPoint1 : Boolean from Standard;
    isPoint2 : Boolean from Standard;    
    myP1     : Pnt2d   from gp;
    myP2     : Pnt2d   from gp;    	
    myC1     : Curve   from Geom2d;
    myC2     : Curve   from Geom2d;
    myOffset : Real    from Standard;
    myBisec  : Bisec   from Bisector;
    myBis    : Curve   from Geom2dAdaptor;
end TrimEdgeTool;
