-- Created on: 1993-03-02
-- Created by: Philippe DAUTRY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SurfaceOfRevolution from PGeom inherits SweptSurface from PGeom

        ---Purpose :  This  class defines    a   complete   surface of
        --         revolution.  The surface is  obtained by rotating a
        --         curve  a  complete revolution  about an axis.   The
        --         curve and the axis must be in the same plane.
        --         
	---See Also : SurfaceOfRevolution from Geom.

uses Dir         from gp,
     Pnt         from gp,
     Curve       from PGeom,
     SurfaceForm from GeomAbs,
     Shape       from GeomAbs

is


  Create returns mutable SurfaceOfRevolution from PGeom;
	---Purpose: Creates a SurfaceOfRevolution with default values.
    	---Level: Internal 


  Create (
    	    aBasisCurve : Curve from PGeom;
    	    aDirection  : Dir from gp;
	    aLocation   : Pnt from gp)
     returns mutable SurfaceOfRevolution from PGeom;
	---Purpose: Creates a SurfaceOfRevolution with these values.
    	---Level: Internal 


  Location (me : mutable; aLocation : Pnt from gp);
        ---Purpose : Set the value of the field location with <aLocation>.
    	---Level: Internal 


  Location (me) returns Pnt from gp;
        ---Purpose : Returns the value of the field location.
    	---Level: Internal 


fields

  location  : Pnt from gp;

end;
