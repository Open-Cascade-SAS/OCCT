-- Created on: 1993-09-08
-- Created by: Christian CAILLET
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DefaultSpecific  from IGESData  inherits SpecificModule

    ---Purpose : Specific IGES Services for UndefinedEntity, FreeFormatEntity

uses IGESEntity, IGESDumper,
     Messenger from Message

is

    Create returns mutable DefaultSpecific;
    ---Purpose : Creates a DefaultSpecific and puts it into SpecificLib

    OwnDump (me; CN : Integer; ent : IGESEntity;
    	      dumper : IGESDumper;  S : Messenger from Message; own : Integer);
    ---Purpose : Specific Dump for UndefinedEntity : it concerns only
    --           own parameters, the general data (Directory Part, Lists) are
    --           taken into account by the IGESDumper

end DefaultSpecific;
