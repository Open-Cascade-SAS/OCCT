-- Created on: 1993-07-01
-- Created by: Gerard GRAS
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Driver from Xw inherits WindowDriver from Aspect

	---Version:

	---Purpose: This class defines a X window Driver.
	--  Warning: A Driver is associated with one window and lets you
    	-- draw any primitives with any attributes you choose
    	-- inside that window. All Values and coordinates are
    	-- defined in Device Window Unit (DWU) space, which is
    	-- the Normalized Floating Pixel space limited by the size
    	-- of the window. The Maps Driver must be initialized
    	-- with Aspect_Driver::SetXXXXMap(aMap) where XXXX
    	-- may correspond to Color, Mark, Type, Width and Font.
    
	---References:

uses

	ExtendedString		from TCollection,
	Length			from Quantity,
	Factor			from Quantity,
	Ratio			from Quantity,
	PlaneAngle		from Quantity,
	Array1OfShortReal	from TShort,
	TypeOfResize		from Aspect,
	TypeOfDrawMode		from Aspect,
	TypeOfText		from Aspect,
	TypeOfPrimitive		from Aspect,
	ColorMap		from Aspect,
	TypeMap			from Aspect,
	WidthMap		from Aspect,
	FontMap			from Aspect,
	MarkMap			from Aspect,
	TypeOfVisual		from Xw,
	Window			from Xw,
	HArray1OfInteger        from TColStd,
	HListOfMFTFonts		from Xw,
	HArray1OfShortReal      from TShort,
	TextManager		from Xw

raises

	DriverDefinitionError	from Aspect,
	DriverError		from Aspect

is

	-------------------------
	-- Category: Constructors
	-------------------------

	Create (aWindow: Window from Xw)
	returns mutable Driver from Xw
	raises DriverDefinitionError from Aspect;
	---Level: Public
	---Purpose: Creates the X Window Driver associated to the X window
	--	    <aWindow>.
	--	    Default values :
	--		- DrawMode : TODM_REPLACE

	---------------------------------------------------
	-- Category: Methods to modify the class definition
	---------------------------------------------------

	BeginDraw (me: mutable;
                   DoubleBuffer: Boolean = Standard_True;
                   aRetainBuffer: Integer = 0)
	---Level: Public
        ---Purpose: Begin graphics and drawn directly to the Window or Pixmap if
        --<aRetainBuffer> is 0 or in the retain buffer if > 0.
                raises DriverError from Aspect is virtual;
        ---Trigger: Raises if the retain buffer is not open.
        --         call BufferIsOpen() method before.
	---Category: Methods to modify the class definition

	EndDraw (me: mutable; Synchronize: Boolean = Standard_False) is virtual;
	---Level: Public
	---Purpose: Called by the method Graphic2d_View::Update, this
	--	    method manages the buffer flushing and Wait after up to date
	--	    display when Synchronize is TRUE.
	---Category: Methods to modify the class definition


	ResizeSpace (me : mutable)
	returns TypeOfResize from Aspect
	---Level: Public
	---Purpose: Resizes the WorkSpace depending of the Window size
	--	    MUST be call after a Resize or Move WindowDriver Event
	--	    Returns the TypeOfResize gravity mode .
	--  Trigger: Raises if the type of resizing is unknown.
	raises DriverError from Aspect is virtual;
	---Category: Methods to modify the class definition

	---------------------------------------------
	-- Category: Methods to define the attributes
	---------------------------------------------

	InitializeColorMap (me: mutable;
			    Colormap: ColorMap from Aspect)
	---Level: Public
	---Purpose: Defines the color map.
	--  Level: Public
	--  Trigger: Raises if the definition failed.
	raises DriverError from Aspect is virtual protected;
	---Category: Methods to define the color indices.

	InitializeTypeMap (me: mutable;
			   Typemap: TypeMap from Aspect)
	---Purpose: Defines the line type map.
	--  Level: Public
	--  Trigger: Raises if the definition failed.
	raises DriverError from Aspect is virtual protected;
	---Category: Methods to define the type of line indices.

	InitializeWidthMap (me: mutable;
			    Widthmap: WidthMap from Aspect)
	---Purpose: Defines the width line map.
	--  Level: Public
	--  Trigger: Raises if the definition failed.
	raises DriverError from Aspect is virtual protected;
	---Category: Methods to define the width of line indices.

	InitializeFontMap (me: mutable;
			   Fontmap: FontMap from Aspect)
	---Purpose: Defines the font map.
	--  Level: Public
	--  Trigger: Raises if the definition failed.
	raises DriverError from Aspect is virtual protected;
	---Category: Methods to define the font indices.

	InitializeMarkMap (me: mutable;
			   Markmap: MarkMap from Aspect)
	---Purpose: Defines the mark map.
	--  Level: Public
	--  Trigger: Raises if the definition failed.
	raises DriverError from Aspect is virtual protected;
	---Category: Methods to define the marker indices.

	---------------------------------------------
	-- Category: Methods to set the attributes
	---------------------------------------------

	SetDrawMode (me:mutable; aMode: TypeOfDrawMode from Aspect) is virtual;
	---Level: Advanced
	---Purpose: Defines the draw mode for all primitives drawing.
	--	TypeOfDrawMode is
	--		TODM_REPLACE
	--		TODM_ERASE
	--		TODM_XOR
	--		TODM_XORLIGHT

	SetLineAttrib (me: mutable;
		       ColorIndex: Integer from Standard;
		       TypeIndex: Integer from Standard;
		       WidthIndex: Integer from Standard)
	---Level: Public
	---Purpose: Sets the line attributes.
	--  Category: Methods to set the line attributes
	--  Trigger: Raises if one of the index is out of range.
	raises DriverError from Aspect is virtual;

	SetTextAttrib (me: mutable;
		       ColorIndex: Integer from Standard;
		       FontIndex: Integer from Standard)
	---Level: Public
	---Purpose: Sets the text attributes.
	--  Category: Methods to set the text attributes
	--  Trigger: Raises if one of the index is out of range.
	raises DriverError from Aspect is virtual;

	SetTextAttrib (me: mutable;
		       ColorIndex: Integer from Standard;
		       FontIndex: Integer from Standard;
		       aSlant: PlaneAngle from Quantity;
		       aHScale: Factor from Quantity;
		       aWScale: Factor from Quantity;
		       isUnderlined: Boolean from Standard = Standard_False)
	---Level: Public
	---Purpose: Sets the Extended text attributes.
	--  Category: Methods to set the text attributes
	--  Trigger: Raises if one of the index is out of range.
	raises DriverError from Aspect is virtual;

	SetPolyAttrib (me: mutable;
		       ColorIndex: Integer from Standard;
		       TileIndex: Integer from Standard;
		       DrawEdgeFlag: Boolean from Standard = Standard_False)
	---Level: Public
	---Purpose: Sets the polygon attributes.
	--  Warning:
	-- <ColorIndex> is the background poly color index.
	-- <TileIndex> is the background poly fill rule index.
	-- If <DrawEdgeFlag> is TRUE the edge of the poly is drawn with the
	--  current line attributes.
	--  Category: Methods to set the poly attributes
	--  Trigger: Raises if one of the index is out of range.
	raises DriverError from Aspect is virtual;

	SetMarkerAttrib (me: mutable;
		       ColorIndex: Integer from Standard;
		       EdgeWidthIndex: Integer from Standard;
		       FillMarker: Boolean from Standard = Standard_False)
	---Level: Public
	---Purpose: Sets the marker attributes.
	--  Warning:
	-- <ColorIndex> is the edge or fill marker color index.
	-- <EdgeWidthIndex> is the edge marker thickness index.
	-- If <FillMarker> is TRUE the marker is filled on the first set
	--  of consecutive drawn points.
	--  Category: Methods to set the marker attributes
	--  Trigger: Raises if one of the index is out of range.
	raises DriverError from Aspect is virtual;

	-----------------------------------------
	-- Category: Methods to manage the images
	-----------------------------------------

	IsKnownImage (me: mutable; anImage: Transient from Standard)
	returns Boolean from Standard is virtual;
	---Level: Public
        ---Purpose: Returns Standard_True if the associated driver
	--	    have stored the image and Standard_False if not.
	---Category: Methods to manage the images

	SizeOfImageFile (me; anImageFile: CString from Standard;
			     aWidth,aHeight: out Integer from Standard)
	returns Boolean from Standard is virtual;
	---Level: Public
        ---Purpose: Returns Standard_True and the Image Size in PIXEL 
	--          if the image file exist and can be computed by the driver,
	--          NOTE that only XWD image file type are recognized today. 
	---Category: Methods to manage the images

	ClearImage (me: mutable; anImageId: Transient from Standard) is virtual;
	---Level: Public
	---Purpose: Clears the image in <me>.
	---Category: Methods to manage the images

	ClearImageFile (me: mutable; anImageFile: CString from Standard) 
								is virtual;
	---Level: Public
	---Purpose: Clears the image associated with the image file .
	---Category: Methods to manage the images

	DrawImage (me: mutable; anImageId: Transient from Standard;
		   aX, aY: ShortReal from Standard)
	---Level: Public
	---Purpose: Draws the image in <me>.
	--	    <aX>, <aY> is the center of the image.
	--	    Image center must be defined in DWU space.
	raises DriverError from Aspect is virtual;
	---Trigger: If the anImageId is not found 
	---Category: Methods to manage the images

	DrawImageFile (me: mutable; anImageFile: CString from Standard;
		   aX, aY: ShortReal from Standard;
		   aScale: Factor from Quantity = 1.0)
	---Level: Public
	---Purpose: Draws the image file in <me>.
	--	    <aX>, <aY> is the center of the image.
	--	    <aScale> the scale factor which is apply on this image
	--	    Image center must be defined in DWU space.
        --	    anImageFile must be defined with the full pathname
 	--          of the form /..../xxxxx.ext or $DIR/xxxxxx.ext
	--          with DIR defined in a setenv variable.
	--               xxxxxx the image file name.
	--               ext the image file extension.
	raises DriverError from Aspect is virtual;
	---Trigger: If the anImageFile is not found 
	--          or the Image type is not an XWD.
	---Category: Methods to manage the images

	FillAndDrawImage (me: mutable; anImageId: Transient from Standard;
			  aX, aY: ShortReal from Standard;
			  Width, Height: Integer from Standard;
			  anArrayOfPixels: Address from Standard)
	---Level: Public
	---Purpose: Stores a complete image and draws it in <me>.
	--	    Image size must be defined in DWU space>
	--  Category: Methods to manage the images
	--  Trigger: Raises if the creation of the image failed.
	raises DriverError from Aspect is virtual;

	FillAndDrawImage (me: mutable; anImageId: Transient from Standard;
			  aX, aY: ShortReal from Standard;
			  anIndexOfLine, Width, Height: Integer from Standard;
			  anArrayOfPixels: Address from Standard)
	---Level: Advanced
	---Purpose: Stores a line of an image and draws it in <me>.
	--  Warning: 0<= anIndexOfLine < aHeight
	--	    anIndexOfLine = 0 must be the first call
	--  Category: Methods to manage the images
	--  Trigger: Raises if the creation of the image failed.
	raises DriverError from Aspect is virtual;

	---------------------------------------
	-- Category: Methods to draw primitives
	---------------------------------------

	DrawPolyline (me : mutable;
		      ListX: Array1OfShortReal from TShort;
		      ListY: Array1OfShortReal from TShort)
	---Level: Public
	---Purpose: Draws the polyline depending of SetLineAttrib() attributes.
	--  Warning: Coordinates must be defined in DWU space.
	--  Trigger: Raises if Polyline has too many points (> 1024)
	--	    Raises if the length of <ListX> is not equal to
	--	    the length of <ListY>.
	raises DriverError from Aspect is virtual;
	---Category: Methods to draw primitives

	DrawPolygon (me : mutable;
		     ListX: Array1OfShortReal from TShort;
		     ListY: Array1OfShortReal from TShort)
	---Level: Public
	---Purpose: Draws the polygone depending of SetPolyAttrib() attributes.
	--  Warning: Coordinates must be defined in DWU space.
	--  Trigger:  Raises if Polygone has too many points (> 1024)
	--	    Raises if the length of <ListX> is not equal to
	--	    the length of <ListY>.
	raises DriverError from Aspect is virtual;
	---Category: Methods to draw primitives

	DrawSegment (me : mutable;
		     X1, Y1: ShortReal from Standard;
		     X2, Y2: ShortReal from Standard)
	---Level: Public
	---Purpose: Draws the segment depending of SetLineAttrib() attributes.
	--  Warning: Coordinates must be defined in DWU space.
	raises DriverError from Aspect is virtual;
	---Category: Methods to draw primitives

	DrawText (me : mutable;
		  Text: ExtendedString from TCollection;
		  Xpos, Ypos: ShortReal from Standard;
		  anAngle: ShortReal from Standard = 0.0;
		  aType: TypeOfText from Aspect = Aspect_TOT_SOLID)
	---Level: Public
	---Purpose: Draws the text depending of SetTextAttrib() attributes.
	--  Category: Methods to draw primitives
	--  Warning: Coordinates must be defined in DWU space.
	--  Trigger: Raises if Text has too many chars (> 1024)
	raises DriverError from Aspect is virtual;

	DrawText (me : mutable;
		  Text: CString from Standard;
		  Xpos, Ypos: ShortReal from Standard;
		  anAngle: ShortReal from Standard = 0.0;
		  aType: TypeOfText from Aspect = Aspect_TOT_SOLID)
	---Level: Public
	---Purpose: Draws the text depending of SetTextAttrib() attributes.
	--  Category: Methods to draw primitives
	--  Warning: Coordinates must be defined in DWU space.
	--	    Angle must be defined in RADIAN.
	--  Trigger: Raises if Text has too many chars (> 1024)
	raises DriverError from Aspect is virtual;

        DrawPolyText (me : mutable;
                  aText: ExtendedString from TCollection;
                  Xpos:  ShortReal from Standard;
                  Ypos:  ShortReal from Standard;
                  aMarge: Ratio from Quantity = 0.1;
                  anAngle: ShortReal from Standard = 0.0;
		  aType: TypeOfText from Aspect = Aspect_TOT_SOLID)
        ---Level: Public
        ---Purpose: Draws an framed text depending of the
        -- SetTextAttrib() and SetPolyAttrib() attributes.
        --  Warning: Coordinates must be defined in DWU space.
        --          <aMarge> defines the ratio of the space between the 
        --          polygon borders and the bounding box of the text and 
	--	    depending of the height of the text. 
                raises DriverError from Aspect is virtual;
        ---Trigger: Raises if Text has too many chars (> 1024)
        --          or <aMarge is < 0 or > 1.
        ---Category: Methods to draw primitives

        DrawPolyText (me : mutable;
                aText: CString from Standard;
                Xpos:  ShortReal from Standard;
                Ypos:  ShortReal from Standard;
                aMarge: Ratio from Quantity = 0.1;
                anAngle: ShortReal from Standard = 0.0;
		aType: TypeOfText from Aspect = Aspect_TOT_SOLID)
        ---Level: Public
        ---Purpose: Draws an framed text depending of the
        -- SetTextAttrib() and SetPolyAttrib() attributes.
        --  Warning: Coordinates must be defined in DWU space.
        --          <aMarge> defines the ratio of the space between the 
        --          polygon borders and the bounding box of the text and 
	--	    depending of the height of the text. 
                raises DriverError from Aspect is virtual;
        ---Trigger: Raises if Text has too many chars (> 1024)
        --          or <aMarge is < 0 or > 1.
        ---Category: Methods to draw primitives

        DrawPoint (me : mutable; X, Y: ShortReal from Standard)
        ---Level: Public
        ---Purpose: Draws a 1 PIXEL point depending of the SetMarkerAttrib() 
	--color attribute or add a point depending of the incremental 
	--BeginXxxxxx() primitive used.
	raises DriverError from Aspect is virtual;
	---Category: Methods to draw primitives

	DrawMarker (me : mutable;
		  aMarker: Integer from Standard;
		  Xpos, Ypos: ShortReal from Standard;
		  Width,Height: ShortReal from Standard;
		  Angle: ShortReal from Standard = 0.0)
	---Level: Public
	---Purpose: Draws the previously defined marker depending of 
	-- the SetMarkerAttrib() attributes.
	--  Warning: Coordinates and sizes must be defined in DWU space.
	--	    Angle must be defined in RADIAN.
	--	    A one pixel marker is drawn when aMarker index is undefined.
	raises DriverError from Aspect is virtual;
	---Category: Methods to draw primitives

        DrawArc (me : mutable; X,Y : ShortReal from Standard;
                        aXradius,aYradius : ShortReal from Standard;
                        aStartAngle: ShortReal from Standard = 0.0;
                        anOpenAngle: ShortReal from Standard = 6.283185)
                                                        returns Boolean
        ---Level: Public
        ---Purpose: Draws an Ellipsoid arc of center <X,Y> and Radius
        --  <aXradius,aYradius> of relative angle <anOpenAngle> from
        --  the base angle <aStartAngle>
        --  Warning: Returns FALSE if the hardware can't drawing this
        --  primitive properly,application must to simulate it.
                raises DriverError from Aspect is virtual;
        ---Trigger: Raises if one of <aXradius,aYradius> is <= 0.

        DrawPolyArc (me : mutable; X,Y : ShortReal from Standard;
                        anXradius,anYradius : ShortReal from Standard;
                        aStartAngle: ShortReal from Standard = 0.0;
                        anOpenAngle: ShortReal from Standard = 6.283185)
                                                        returns Boolean
        ---Level: Public
        ---Purpose: Draws an filled Ellipsoid arc of center <X,Y> and Radius
        --  <anXradius,anYradius> of relative angle <anOpenAngle> from
        --  the base angle <aStartAngle> and  depending of the SetPolyAttrib()
	-- attributes.
        --  Warning: Returns FALSE if the hardware can't drawing this
        --  primitive properly,application must to simulate it.
                raises DriverError from Aspect is virtual;
        ---Trigger: Raises if one of <aXradius,aYradius> is <= 0.
 
        BeginPolyline (me : mutable; aNumber : Integer) is virtual;
        ---Level: Public
        ---Purpose: Begin a polyline primitive of <aNumber> of points .
	--  Warning: Points must be added by the DrawPoint() method.
 
        BeginPolygon (me : mutable; aNumber : Integer) is virtual;
        ---Level: Public
        ---Purpose: Begin a polygon primitive of <aNumber> of points .
	--  Warning: Points must be added by the DrawPoint() method.
 
        BeginSegments (me : mutable) is virtual;
        ---Level: Public
        ---Purpose: Begin a set of segments .
	--  Warning: Segments must be added by DrawSegment() method.

        BeginArcs (me : mutable) is virtual;
        ---Level: Public
        ---Purpose: Begin a set of circles or ellips .
        --  Warning: Arcs must be added by the DrawArc() method.
 
        BeginPolyArcs (me : mutable) is virtual;
        ---Level: Public
        ---Purpose: Begin a set of polygon circles or ellips .
        --  Warning: Arcs must be added by the DrawPolyArc() method.
 
        BeginMarkers (me : mutable) is virtual;
        ---Level: Public
        ---Purpose: Begin a set of markers .
        --  Warning: Markers must be added by the DrawMarker() method.
 
        BeginPoints (me : mutable) is virtual;
        ---Level: Public
        ---Purpose: Begin a set of points .
        --  Warning: Points must be added by the DrawPoint() method.
  
        ClosePrimitive (me : mutable)
        ---Level: Public
        ---Purpose: Close the last Begining primitive
                raises DriverError from Aspect is virtual;
        ---Trigger: Raises if no primitive have been opened by BeginXxxxxx().

	---------------------------------------
	-- Category: Methods to Manage buffers
	---------------------------------------

        OpenBuffer (me : mutable; aRetainBuffer: Integer;
                                 aPivotX: ShortReal = 0.0;
                                 aPivotY: ShortReal = 0.0;
				 aWidthIndex: Integer = 0;
				 aColorIndex: Integer = 0;
				 aFontIndex: Integer = 0; 
                                 aDrawMode: TypeOfDrawMode = Aspect_TODM_REPLACE)                                                          
                                        returns Boolean is virtual;
        ---Purpose: Allocate the retain buffer <aRetainBuffer> ,   
        -- Defines the DWU coordinates of the pivot point for all primitives
        --  contains inside.
        -- Defines the buffer color, line width and font index :
        --  the default color is the highlight color of the colormap.
        --  the default font is the default system font of the fontmap. 
        -- The other attributes are fixed :
        --  line type is Solid,
        --  line width is 1 Pixel,
        --  polygon fill mode is Solid,   
        --  Warning: The number of allocated buffers is limited,it's 
        --  recommended to close unused buffers some time!  
        --          The TypeOfDrawMode REPLACE is enabled only if the 
        --          background drawing has been drawn with the DoubleBuffer
        --          flag set to ENABLE at the last BeginDraw time. 
        --          The TypeOfDrawMode XOR is enabled in any case.
        --          The other TypeOfDrawMode are not authorized. 
        -- Returns TRUE if the buffer is allocated and enabled for drawing.
 
        CloseBuffer (me; aRetainBuffer: Integer)
        ---Purpose: Clear & Deallocate the retain buffer <aRetainBuffer>.
                raises DriverError from Aspect is virtual;
        ---Trigger: Raises if the retain buffer is not opened.
        --         call BufferIsOpen() method before.
 
        ClearBuffer (me; aRetainBuffer: Integer)
        ---Purpose: Erase & Clear ALL primitives retains in the buffer <aRetainBuffer>.
                raises DriverError from Aspect is virtual;
        ---Trigger: Raises if the retain buffer is not opened.
        --         call BufferIsOpen() method before.
 
        DrawBuffer (me; aRetainBuffer: Integer)
        ---Purpose: Draw ALL primitives retains in the buffer <aRetainBuffer>.
        --  Warning: Note that the aspect of a retain buffer drawing is mono-colored
        -- with the current buffer attributes and
        -- depending of the DoubleBuffer state flag at the BeginDraw() buffer time,
        -- when DB is TRUE,an XOR method is use for drawing and erasing buffers in the
        -- same way.In this case,some color side effect can occurs depending of the
        -- traversal primitive colors and the supported hardware.
        -- when DB is FALSE and the background drawing has been generated with
        -- DB at TRUE,no color side effect occurs because the DB is used for restoring
        -- the drawing context at EraseBuffer() time,this is more powerfull for the
        -- drawing quality excepted for large buffers (flicking) .
                raises DriverError from Aspect is virtual;
        ---Trigger: Raises if the retain buffer is not opened.
        --         call BufferIsOpen() method before.

        EraseBuffer (me; aRetainBuffer: Integer)
        ---Purpose: Erase ALL primitives retains in the buffer <aRetainBuffer>.
                raises DriverError from Aspect is virtual;
        ---Trigger: Raises if the retain buffer is not opened.
        --         call BufferIsOpen() method before.
 
        MoveBuffer (me; aRetainBuffer: Integer;
                                 aPivotX: ShortReal = 0.0;
                                 aPivotY: ShortReal = 0.0)
        ---Purpose: Erase , Translate and reDraw ALL primitives retains in the buffer
        --<aRetainBuffer>.
        --<aPivotX,aPivotY> are the new DWU attached point absolute coordinates
        --of the buffer pivot point.
                raises DriverError from Aspect is virtual;
        ---Trigger: Raises if the retain buffer is not opened.
        --         call BufferIsOpen() method before.
 
        ScaleBuffer (me; aRetainBuffer: Integer; aScaleX: Factor = 1.0;
                                                          aScaleY: Factor = 1.0)
        ---Purpose: Erase , Scale the buffer from the Pivot point and reDraw ALL primitives
        --retains in the buffer <aRetainBuffer>.
        -- The transformation is relative since the creation time of the buffer.
        --<aScaleX,aScaleY> are the relative scale factors apply on the two axis.
        --  Warning: Note that the scalling of some primitives can provided some bad
        --smoothing side effect (i.e: Circles,...)
                raises DriverError from Aspect is virtual;
        ---Trigger: Raises if the retain buffer is not opened or
        --one of <aScale> factor is <= 0.
        --         call BufferIsOpen() method before.
  
        RotateBuffer (me; aRetainBuffer: Integer; anAngle: PlaneAngle = 0.0)
        ---Purpose: Erase , Rotate the buffer from the Pivot point and reDraw ALL primitives
        --  retains in the buffer <aRetainBuffer>.
        -- The transformation is relative since the creation time of the buffer.
        --  <anAngle> is the relative counter-clockwise rotation angle from the
        --  Horizontal axis.
                raises DriverError from Aspect is virtual;
        ---Trigger: Raises if the retain buffer is not opened.
        --         call BufferIsOpen() method before.

	----------------------------
	-- Category: Inquire methods
	----------------------------

	WorkSpace (me; Width, Heigth: out Length from Quantity) is virtual;
	---Level: Public
	---Purpose: Returns the Available WorkSpace in DWU coordinates
	--  Category: Inquire methods

        TextSize (me; aText: ExtendedString from TCollection;
                      aWidth, aHeight: out ShortReal from Standard;
                      aFontIndex: Integer from Standard = -1)
                raises DriverError from Aspect is virtual;
        ---Level: Public
        ---Purpose: Returns the TEXT size in DWU space depending
        --          of the required FontIndex if aFontIndex is >= 0
        --          or the current FontIndex if < 0 (default).
        ---Category: Inquire methods

        TextSize (me; aText: ExtendedString from TCollection;
                      aWidth, aHeight, anXoffset, anYoffset: out ShortReal from Standard;
                      aFontIndex: Integer from Standard = -1)
                raises DriverError from Aspect is virtual;
        ---Level: Public
        ---Purpose: Returns the extended TEXT size and offsets 
	--	    in DWU space depending
        --          of the required FontIndex if aFontIndex is >= 0
        --          or the current FontIndex if < 0 (default).
        --          NOTE that the text offsets defines the relative position of the
        --         of the text string origin from the lower left corner of the text
        --         boundary limits.
        ---Category: Inquire methods

        TextSize (me; aText: CString from Standard;
                      aWidth, aHeight, anXoffset, anYoffset: out ShortReal from Standard;
                      aFontIndex: Integer from Standard = -1)
                raises DriverError from Aspect is virtual;
        ---Level: Public
        ---Purpose: Returns the ascii TEXT size and offsets 
	--	    in DWU space depending
        --          of the required FontIndex if aFontIndex is >= 0
        --          or the current FontIndex if < 0 (default).
        --          NOTE that the text offsets defines the relative position of the
        --         of the text string origin from the lower left corner of the text
        --         boundary limits.
        ---Category: Inquire methods
 
        FontSize (me; aSlant: out PlaneAngle from Quantity;
                      aSize,aBheight: out ShortReal from Standard;
                      aFontIndex: Integer from Standard = -1)
                                returns CString from Standard
        ---Trigger: Raises if font is not defined.
        	raises DriverError from Aspect is virtual;
        ---Level: Public
        ---Purpose: Returns the font string,slant,size and
        --  baseline height in DWU space depending
        --          of the required FontIndex if aFontIndex is >= 0
        --          or the current FontIndex if < 0 (default).
        ---Category: Inquire methods

	Convert (me; PV: Integer from Standard)
	returns Length from Quantity is virtual;
	---Level: Public
	---Purpose: Returns the DWU value depending of
	--	    the PIXEL value.
	---Category: Inquire methods

	Convert (me; DV: Length from Quantity)
	returns Integer from Standard is virtual;
	---Level: Public
	---Purpose: Returns the PIXEL value depending of
	--	    the DWU value.
	---Category: Inquire methods

	Convert (me; PX, PY: Integer from Standard;
		 DX, DY: out Length from Quantity) is virtual;
	---Level: Public
	---Purpose: Returns the DWU position depending of
	--	    the PIXEL position .
	---Category: Inquire methods

	Convert (me; DX, DY: Length from Quantity;
		 PX, PY: out Integer from Standard) is virtual;
	---Level: Public
	---Purpose: Returns the PIXEL position depending of
	--	    the DWU position .
	---Category: Inquire methods

        BufferIsOpen(me; aRetainBuffer : Integer) returns Boolean is virtual;
        ---Purpose: Returns TRUE if the retain buffer <aRetainBuffer> is enabled
        --for drawing.
 
        BufferIsEmpty(me; aRetainBuffer : Integer) returns Boolean is virtual;
        ---Purpose: Returns TRUE if the retain buffer has not been opened or empty.
        ---         Returns FALSE if a lot of primitives have been stored inside 
	--         because a BeginDraw(..,<aRetainBuffer>) has been done previously.
 
        BufferIsDrawn(me; aRetainBuffer : Integer) returns Boolean is virtual;
        ---Purpose: Returns TRUE if the retain buffer s actually displayed at screen.

        AngleOfBuffer(me; aRetainBuffer : Integer; anAngle: out PlaneAngle)
        ---Purpose: Returns the current buffer rotate angle from the X axis.
                raises DriverError from Aspect is virtual;
        ---Trigger: Raises if the retain buffer is not opened.
        --         call BufferIsOpen() method before.
 
        ScaleOfBuffer(me; aRetainBuffer : Integer; aScaleX,aScaleY: out Factor)
        ---Purpose: Returns the current buffer scale factors.
                raises DriverError from Aspect is virtual;
        ---Trigger: Raises if the retain buffer is not opened.
        --         call BufferIsOpen() method before.
 
        PositionOfBuffer(me; aRetainBuffer : Integer; aPivotX,aPivotY: out ShortReal )
        ---Purpose: Returns the current buffer position.
                raises DriverError from Aspect is virtual;
        ---Trigger: Raises if the retain buffer is not opened.
        --         call BufferIsOpen() method before.

        ColorBoundIndexs(me; aMinIndex,aMaxIndex : out Integer from Standard)
                                                                is virtual;
        ---Level: Advanced
        ---Purpose:
        -- Returns the min and max driver virtual color indexs.
        ---Category: Inquire methods
 
        LocalColorIndex(me; anIndex : Integer from Standard)
                                returns Integer from Standard is virtual;
        ---Level: Advanced
        ---Purpose:
        -- Returns the local colormap hardware index from a virtual driver color       
  -- index or returns -1 if the index is not defined.
        ---Category: Inquire methods
 
        FontBoundIndexs(me; aMinIndex,aMaxIndex : out Integer from Standard)
                                                                is virtual;
        ---Level: Advanced
        ---Purpose:
        -- Returns the min and max driver virtual font indexs.
        ---Category: Inquire methods
 
        LocalFontIndex(me; anIndex : Integer from Standard)
                                returns Integer from Standard is virtual;
        ---Level: Advanced
        ---Purpose:
        -- Returns the associated fontmap hardware index from a virtual driver font
        -- index or returns -1 if the index is not defined.
        ---Category: Inquire methods

        TypeBoundIndexs(me; aMinIndex,aMaxIndex : out Integer from Standard)
                                                                is virtual;
        ---Level: Advanced
        ---Purpose:
        -- Returns the min and max driver virtual type indexs.
        ---Category: Inquire methods
 
        LocalTypeIndex(me; anIndex : Integer from Standard)
                                returns Integer from Standard is virtual;
        ---Level: Advanced
        ---Purpose:
        -- Returns the associated typemap hardware index from a virtual driver type
        -- index or returns -1 if the index is not defined.
        ---Category: Inquire methods
 
        WidthBoundIndexs(me; aMinIndex,aMaxIndex : out Integer from Standard)
                                                                is virtual;
        ---Level: Advanced
        ---Purpose:
        -- Returns the min and max driver virtual width indexs.
        ---Category: Inquire methods
 
        LocalWidthIndex(me; anIndex : Integer from Standard)
                                returns Integer from Standard is virtual;
        ---Level: Advanced
        ---Purpose:
        -- Returns the associated widthmap hardware index from a virtual driver width
        -- index or returns -1 if the index is not defined.
        ---Category: Inquire methods

        MarkBoundIndexs(me; aMinIndex,aMaxIndex : out Integer from Standard)
                                                                is virtual;
        ---Level: Advanced
        ---Purpose:
        -- Returns the min and max driver virtual marker indexs.
        ---Category: Inquire methods
 
        LocalMarkIndex(me; anIndex : Integer from Standard)
                                returns Integer from Standard is virtual;
        ---Level: Advanced
        ---Purpose:
        -- Returns the local markmap hardware index from a virtual driver marker        -- index or returns -1 if the index is not defined.
        ---Category: Inquire methods
  
	----------------------------
	-- Category: Private methods
	----------------------------

	PrintError(myclass) is protected;
	---Purpose: Print last error or raise depending of the error gravity.

	DrawRectangle(me; Xpos,Ypos,Angle,Xoffset,Yoffset,Width,Height: 
				ShortReal from Standard) is private;
	---Purpose: Draw an oriented rectangle

	FillRectangle(me; Xpos,Ypos,Angle,Xoffset,Yoffset,Width,Height: 
				ShortReal from Standard) is private;
	---Purpose: Draw an oriented fill rectangle

fields

	MyVisualClass:		TypeOfVisual from Xw is protected;
	MyExtendedDrawable:	Address from Standard is protected;
	MyExtendedColorMap:	Address from Standard is protected;
	MyExtendedTypeMap:	Address from Standard is protected;
	MyExtendedWidthMap:	Address from Standard is protected;
	MyExtendedFontMap:	Address from Standard is protected;
	MyExtendedMarkMap:	Address from Standard is protected;
	MyImage:		Address from Standard is protected;

	MyLineColor:		Integer from Standard is protected;
	MyLineType:		Integer from Standard is protected;
	MyLineWidth:		Integer from Standard is protected;
	MyPolyColor:		Integer from Standard is protected;
	MyPolyType:		Integer from Standard is protected;
	MyPolyTile:		Integer from Standard is protected;
	MyTextColor:		Integer from Standard is protected;
	MyTextFont:		Integer from Standard is protected;
	MyTextType:		Integer from Standard is protected;
	MyTextHScale:		Real from Standard is protected;
	MyTextWScale:		Real from Standard is protected;
	MyTextHSize:		Real from Standard is protected;
	MyTextWSize:		Real from Standard is protected;
	MyTextSlant:		Real from Standard is protected;
	MyTextMinHeight:	Real from Standard is protected;
	MyTextIsUnderlined:	Boolean from Standard is protected;
	MyMarkerColor:		Integer from Standard is protected;
	MyMarkerType:		Boolean from Standard is protected;
	MyMarkerWidth:		Integer from Standard is protected;

	MyColorIndexs:		HArray1OfInteger from TColStd is protected;
	MyTypeIndexs:		HArray1OfInteger from TColStd is protected;
	MyWidthIndexs:		HArray1OfInteger from TColStd is protected;
	MyFontIndexs:		HArray1OfInteger from TColStd is protected;
	MyMarkerIndexs:		HArray1OfInteger from TColStd is protected;

	MyPrimitiveType:	TypeOfPrimitive from Aspect is protected;
	MyMFTFonts:		HListOfMFTFonts from Xw is protected;
	MyMFTSizes:		HArray1OfShortReal from TShort is protected;
	MyTextManager:		TextManager from Xw is protected;

end Driver from Xw;
