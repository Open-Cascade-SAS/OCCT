-- Created on: 1994-10-25
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PointGeomTool from TopOpeBRep

    ---Purpose: Provide services needed by the Fillers

uses

     VPointInter from TopOpeBRep,         -- Value(), Tolerance()
     Point2d from TopOpeBRep,             -- Value(), Tolerance()
     FaceEdgeIntersector from TopOpeBRep, -- Value(), Tolerance()
     Point from TopOpeBRepDS,
     Point from TopOpeBRepDS,
     Shape from TopoDS

is

    Create returns PointGeomTool from TopOpeBRep;

    MakePoint(myclass; IP : VPointInter from TopOpeBRep)
    returns Point from TopOpeBRepDS;

    MakePoint(myclass; P2D : Point2d from TopOpeBRep)
    returns Point from TopOpeBRepDS;

    MakePoint(myclass; FEI : FaceEdgeIntersector from TopOpeBRep)
    returns Point from TopOpeBRepDS;

    MakePoint(myclass; S : Shape from TopoDS)
    returns Point from TopOpeBRepDS;
		       
    IsEqual(myclass; DSP1,DSP2 : Point from TopOpeBRepDS) 
    returns Boolean from Standard;

end PointGeomTool from TopOpeBRep;
