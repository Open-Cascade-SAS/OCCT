-- Created on: 1996-01-30
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class GluedShape from LocOpe inherits GeneratedShape from LocOpe

	---Purpose: 

uses Shape  from TopoDS,
     Face   from TopoDS,
     Wire   from TopoDS,
     Edge   from TopoDS,
     Vertex from TopoDS,
     ListOfShape         from TopTools,
     MapOfShape          from TopTools,
     DataMapOfShapeShape from TopTools

is

    Create
    
    	returns mutable GluedShape from LocOpe;


    Create(S: Shape from TopoDS)
    
    	returns mutable GluedShape from LocOpe;
    

    Init(me: mutable; S: Shape from TopoDS)
    
    	is static;


    GlueOnFace(me: mutable; F: Face from TopoDS)
    
    	is static;


    MapEdgeAndVertices(me: mutable)
    
    	is static private;


    GeneratingEdges(me: mutable)
    
    	returns ListOfShape from TopTools
	---C++: return const&
	;


    Generated(me: mutable; V: Vertex from TopoDS)
	---Purpose: Returns the  edge  created by  the  vertex <V>. If
	--          none, must return a null shape.
    	returns Edge from TopoDS
	;


    Generated(me: mutable; E: Edge from TopoDS)
	---Purpose: Returns the face created by the edge <E>. If none,
	--          must return a null shape.
    	returns Face from TopoDS
	;


    OrientedFaces(me: mutable)
	---Purpose: Returns  the  list of correctly oriented generated
	--          faces. 
    	returns ListOfShape from TopTools
	---C++: return const&
	;


fields

    myShape  : Shape               from TopoDS;
    myMap    : MapOfShape          from TopTools;
    myGShape : DataMapOfShapeShape from TopTools;

end GluedShape;
