-- Created on: 1992-10-13
-- Created by: Ramin BARRETO
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Updated      J.P. TIRAULT, M. MERCIEN Nov,25 1992
--              Adding classes 
--               - Array1
--               - Array2
-- Updated      R.LEQUETTE Jan 1993
--              Adding of modifying classes 
--               - Sequence, HSequence
--               - Set, HSet
--               - List
--               - Stack
--               - BasicMap, BasicMapIterator
--               - Map, DataMap, DoubleMap, IndexedMap, IndexedDataMap

package TCollection

    	---Purpose: The package <TCollection> provides the services for the 
    	-- transient basic data structures.

uses
    Standard,
    MMgt
is
    class AsciiString;

    class ExtendedString;
    
    class HAsciiString;

    class HExtendedString;
    
    generic class Array1;

    generic class HArray1;
    
    generic class Array2;
    
    generic class HArray2;
    
    generic class Stack, StackNode, StackIterator;
	---Purpose: A stack handled by value.
   
    generic class List, ListNode, ListIterator;
	---Purpose: A single list handled by value.

    class BaseSequence;
    class SeqNode;
    pointer SeqNodePtr to SeqNode from TCollection;
    generic class Sequence,SequenceNode;
	---Purpose: An indexed double list handled by value.
     
    generic class HSequence;
	---Purpose: An indexed double list handle by reference.

    generic class Set, SetIterator, SetList;
	---Purpose: A small set handled by value.

    generic class HSet;
	---Purpose: A small set handled by reference.

    generic class MapHasher;
	---Purpose: A Tool to instantiate Maps. Providing HashCode and
	-- Comparisons on Keys.
    
    private deferred class BasicMap;
    private class MapNode;
    pointer MapNodePtr to MapNode from TCollection;
    ---Purpose: Basic class root of all the Maps.
    
    private deferred class BasicMapIterator;
	---Purpose: Basic class root of all the Iterators on Maps.
    
    generic class Map, MapIterator,StdMapNode;
	---Purpose: A Hashed map to store keys.

    generic class DataMap, DataMapIterator,DataMapNode;
	---Purpose: A Map where data can be stored with the keys.
	
    generic class DoubleMap, DoubleMapIterator, DoubleMapNode;
	---Purpose: A Map to store pair of keys.
	
    generic class IndexedMap,IndexedMapNode;
	---Purpose: A Map where the keys are indexed.
	
    generic class IndexedDataMap,IndexedDataMapNode;
	---Purpose: An Indexed Map where data can be stored with the keys.

    enumeration Side is Left , Right;
    
    deferred generic class Compare ;
        ---Purpose: Defines a comparison operator which can be used by
        -- any ordered structure.   The  way to compare items
        -- has  to be described  in  subclasses, which  herit
        -- from instantiations of Compare.

    private deferred class PrivCompareOfInteger 
            instantiates Compare from TCollection(Integer from Standard); 

    private deferred class PrivCompareOfReal 
            instantiates Compare from TCollection(Real from Standard); 

    class CompareOfInteger;
	
    class CompareOfReal;
    

    NextPrimeForMap(I : Integer) returns Integer;
	---Purpose: Returns a  prime number greater than  <I> suitable
	-- to dimension a Map.  When  <I> becomes great there
	-- is  a  limit on  the  result (today  the  limit is
	-- around 1 000 000). This is not a limit of the number of
	-- items but a limit in the number  of buckets.  i.e.
	-- there will be more collisions  in  the map.

end TCollection;






