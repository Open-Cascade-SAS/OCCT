-- Created on: 1996-09-04
-- Created by: Christian CAILLET
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class FinderProcess  from Transfer  inherits ProcessForFinder

    ---Purpose : Adds specific features to the generic definition :
    --           PrintTrace is adapted

uses InterfaceModel from Interface, 
     Messenger from Message,
     Finder, TransientMapper

is

    Create (nb : Integer = 10000) returns mutable FinderProcess;
    ---Purpose : Sets FinderProcess at initial state, with an initial size

    SetModel (me : mutable; model : InterfaceModel);
    ---Purpose : Sets an InterfaceModel, which can be used during transfer
    --           for instance if a context must be managed, it is in the Model

    Model (me) returns InterfaceModel;
    ---Purpose : Returns the Model which can be used for context

    NextMappedWithAttribute (me; name : CString; num0 : Integer) returns Integer;
    ---Purpose : In the list of mapped items (between 1 and NbMapped),
    --           searches for the first mapped item which follows <num0>
    --           (not included) and which has an attribute named <name>
    --           The considered Attributes are those brought by Finders,i.e.
    --           by Input data.
    --           While NextItemWithAttribute works on Result data (Binders)
    --           
    --           Hence, allows such an iteration
    --           
    --           for (num = FP->NextMappedWithAttribute(name,0);
    --                num > 0;
    --                num = FP->NextMappedWithAttribute(name,num) {
    --                .. process mapped item <num>
    --           }

    TransientMapper (me; obj : Transient) returns TransientMapper;
    ---Purpose : Returns a TransientMapper for a given Transient Object
    --           Either <obj> is already mapped, then its Mapper is returned
    --           Or it is not, then a new one is created then returned, BUT
    --             it is not mapped here (use Bind or FindElseBind to do this)


    PrintTrace (me; start : Finder; S : Messenger from Message)  is redefined;
    ---Purpose : Specific printing to trace a Finder (by its method ValueType)

    PrintStats (me; mode : Integer; S : Messenger from Message);
    ---Purpose : Prints statistics on a given output, according mode

fields

    themodel : InterfaceModel;

end FinderProcess;
