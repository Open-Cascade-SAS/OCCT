-- Created on: 1993-01-09
-- Created by: CKY / Contract Toubro-Larsen ( TCD )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class NominalSize from IGESGraph  inherits IGESEntity

        ---Purpose: defines IGESNominalSize, Type <406> Form <13>
        --          in package IGESGraph
        --
        --          Specifies a value, a name, and optionally a
        --          reference to an engineering standard

uses

        HAsciiString from TCollection

is

        Create returns mutable NominalSize;

        -- Specific Methods pertaining to the class

        Init (me                : mutable;
              nbProps           : Integer;
              aNominalSizeValue : Real;
              aNominalSizeName  : HAsciiString from TCollection;
              aStandardName     : HAsciiString from TCollection);
        ---Purpose : This method is used to set the fields of the class
        --           NominalSize
        --      - nbProps           : Number of property values (2 or 3)
        --      - aNominalSizeValue : NominalSize Value
        --      - aNominalSizeName  : NominalSize Name
        --      - aStandardName     : Name of relevant engineering standard

        NbPropertyValues  (me) returns Integer;
        ---Purpose : returns the number of property values in <me>

        NominalSizeValue (me) returns Real;
        ---Purpose : returns the value of <me>

        NominalSizeName (me) returns HAsciiString from TCollection;
        ---Purpose : returns the name of <me>

        HasStandardName (me) returns Boolean;
        ---Purpose : returns True if an engineering Standard is defined for <me>
        -- else, returns False

        StandardName (me) returns HAsciiString from TCollection;
        ---Purpose : returns the name of the relevant engineering standard of <me>

fields

--
-- Class    : IGESGraph_NominalSize
--
-- Purpose  : Declaration of the variables specific to a Nominal Size.
--
-- Reminder : A Nominal Size is defined by :
--            - Number of property values
--            - Value
--            - Name
--            - Name of relevant engineering standard
--

        theNbPropertyValues : Integer;

        theNominalSizeValue : Real;

        theNominalSizeName  : HAsciiString from TCollection;

        theStandardName     : HAsciiString from TCollection;

end NominalSize;
