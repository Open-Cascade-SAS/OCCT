-- Created on: 1995-08-25
-- Created by: Remi LEQUETTE
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class HCurve from Geom2dAdaptor inherits GHCurve from Geom2dAdaptor

	---Purpose: Provides an interface between the services provided by any
    	-- curve from the package Geom2d and those required
    	-- of the curve by algorithms, which use it.

uses
    Curve from Geom2d,
    Curve from Geom2dAdaptor

raises
    ConstructionError from Standard

is

    Create returns mutable HCurve from Geom2dAdaptor;
    
    Create( AS : Curve from Geom2dAdaptor) returns mutable HCurve from Geom2dAdaptor;

    Create( S : Curve from Geom2d) returns mutable HCurve from Geom2dAdaptor;
    
    Create( S : Curve from Geom2d; UFirst,ULast : Real) 
    returns  mutable HCurve from Geom2dAdaptor
    raises ConstructionError from Standard;
    	---Purpose: ConstructionError is raised if UFirst>ULast or VFirst>VLast

end HCurve;
