-- Created on: 1991-09-06
-- Created by: NW,JPB,CAL
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class ClipPlane from Visual3d inherits TShared

	---Version:

	---Purpose: This class allows the definition and update
	--	    of clipping planes in the space model.

	---Keywords: Clipping Plane, Model Clipping

	---Warning:
	---References:

uses

	CPlane	from Graphic3d

is

	Create ( ACoefA		: Real from Standard;
		 ACoefB		: Real from Standard;
		 ACoefC		: Real from Standard;
		 ACoefD		: Real from Standard )
		returns mutable ClipPlane from Visual3d;
	---Level: Internal
	---Purpose: Creates a clipping plane from the equation :
	--	    <ACoefA>*X + <ACoefB>*Y + <ACoefC>*Z + <ACoefD> = 0.0

	---------------------------------------------------
	-- Category: Methods to modify the class definition
	---------------------------------------------------

	SetPlane ( me		: mutable;
		   ACoefA	: Real from Standard;
		   ACoefB	: Real from Standard;
		   ACoefC	: Real from Standard;
		   ACoefD	: Real from Standard )
		is static;
	---Level: Internal
	---Purpose: Modifies the plane equation.
	---Category: Methods to modify the class definition

	--------------------------
	-- Category: Class methods
	--------------------------

	Limit ( myclass )
		returns Integer from Standard;
	---Level: Internal
	---Purpose: Maximum number of activatable clipping planes.
	---Category: Class methods

	----------------------------
	-- Category: Inquire methods
	----------------------------

	Plane ( me;
		ACoefA	: out Real from Standard;
		ACoefB	: out Real from Standard;
		ACoefC	: out Real from Standard;
		ACoefD	: out Real from Standard )
		is static;
	---Level: Internal
	---Purpose: Returns the values of the clipping plane <me>.
	---Category: Inquire methods

	----------------------------
	-- Category: Private methods
	----------------------------

	Identification ( me )
		returns Integer from Standard
		is static private;
	---Level: Internal
	---Purpose: Returns the plane identification.
	---Category: Private methods

--

fields

--
-- Class	:	Visual3d_ClipPlane
--
-- Purpose	:	Declaration of variables specific to the
--			clipping plane model
--
-- Reminders	:	A clipping plane is defined by its equation
--			Equation : A*X + B*Y + C*Z + D = 0
--

	-- the associated C structure
	MyCPlane	:	CPlane from Graphic3d;

friends

	class View from Visual3d

end ClipPlane;
