-- Created on: 1995-03-22
-- Created by: Christophe MARION
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class VData from HLRTopoBRep

uses
    Real  from Standard,
    Shape from TopoDS

is
    Create returns VData from HLRTopoBRep;
    	---C++: inline
	
    Create (P : Real; V : Shape from TopoDS)
    returns VData from HLRTopoBRep;
	
    Parameter(me) returns Real from Standard
    	---C++: inline
    is static;
	
    Vertex(me) returns Shape from TopoDS
    	---C++: inline
    	---C++: return const &
    is static;

fields
    myParameter : Real  from Standard;
    myVertex    : Shape from TopoDS;

end VData;
