-- Created on: 1995-10-06
-- Created by: Jing Cheng MEI
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ShapeDirPresentation from DsgPrs

	---Purpose: A framework to define display of the normal to the
    	-- surface of a shape.

uses
    Shape  from TopoDS,
    Presentation from Prs3d,
    Drawer from Prs3d
    
is

    Add(myclass; prs: Presentation from Prs3d;
                 aDrawer: Drawer from Prs3d;
    	    	 shape: Shape from TopoDS; 
                 mode: Integer from Standard);
    	---Purpose: Adds the shape shape and the mode mode to the
    	-- presentation object prs.
    	-- The display attributes of the normal are defined by the
    	-- attribute manager aDrawer.
    	-- mode determines whether the first or the last point of
    	-- the normal is given to the presentation object. If the
    	-- first point: 0; if the last point, 1.
        
end ShapeDirPresentation;
