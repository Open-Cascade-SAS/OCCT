-- Created on: 1992-04-13
-- Created by: Isabelle GRIGNON
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package IntImp

	---Purpose: 

uses Standard, TColStd, StdFail, math, gp, IntSurf

is

    enumeration ConstIsoparametric is
                UIsoparametricOnCaro1, VIsoparametricOnCaro1,
                UIsoparametricOnCaro2, VIsoparametricOnCaro2;
		
    deferred generic class PSurfaceTool;

    deferred generic class ISurfaceTool;

    deferred generic class CurveTool;

    deferred generic class CSCurveTool;

    deferred generic class COnSCurveTool;

    generic class ZerImpFunc; -- inherits FunctionSetWithDerivatives
    
    generic class ZerParFunc; -- inherits FunctionSetWithDerivatives

    deferred generic class CSFunction; -- inherits FunctionSetWithDerivatives

    generic class ZerCSParFunc; -- inherits FunctionSetWithDerivatives
    
    generic class ZerCOnSSParFunc; -- inherits FunctionSetWithDerivatives
    
    generic class Int2S,TheFunction;
    
    generic class IntCS;

end IntImp;
