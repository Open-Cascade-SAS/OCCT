-- Created on: 1993-03-08
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Update:      Frederic Maupas


package PTopoDS 

	---Purpose: The package PTopoDS provides persistent classes to
	--          store Topological Data Structures in Data Base.
	--          
	--          The  structure  of  this  persistent  topology  is
	--          similar  to   the  transient  topology   (see  its
	--          documentation for more comprehension of this one).
	--          But some differences occure:
	--          
	--          * The class Model and derivatives disappear;
	--          
	--          * The "free"  information  disappears,  because  a 
	--          TShape stored in the Data Base is always "frozen";
	--          

	--          * The class HShape  inherits  from ExternShareable  from
	--          ObjMgt,  so that an intance of HShape  may be
	--          shared by a TShape even if the HShape is not in the
	--          same Container.
	--          
	--          * The class Shape1 inherits from Storable from
	--          Standard.
	--          
	--          Note that the  use of this topology is managed  by
	--          the package MgtTopoDS.
	--          
	--          About the question of "Location", see the  package
	--          PTopLoc  itself;  about  naming,  referencing  and
	--          using persistent  Shapes outsing  the  topological
	--          world, see the package TopoDB.

uses

    ObjMgt,
    Standard,
    TopAbs,      -- basic enumerations : ShapeEnum, Orientation
    PTopLoc,     -- Persistent local coordinate systems
    PCollection,
    TCollection
    
is

    ---Category: Old version of Shape/TShape.
    --           ============================

    class HShape;

    deferred class TShape;

    deferred class TVertex;

    class Vertex;

    deferred class TEdge;

    class Edge;

    class TWire;

    class Wire;

    class TFace;

    class Face;

    class TShell;

    class Shell;

    class TSolid;

    class Solid;

    class TCompSolid;

    class CompSolid;

    class TCompound;

    class Compound;


    class HArray1OfHShape instantiates HArray1 from PCollection
    	(HShape from PTopoDS);


    ---Category: New version of Shape/TShape.
    --           ============================

    class Shape1;

    deferred class TShape1;

    deferred class TVertex1;

    deferred class TEdge1;

    class TWire1;

    class TFace1;

    class TShell1;

    class TSolid1;


    class TCompSolid1;

    class TCompound1;

    class HArray1OfShape1 instantiates HArray1 from PCollection
    	(Shape1 from PTopoDS);

end PTopoDS;
