-- Created on: 1992-03-09
-- Created by: Isabelle GRIGNON
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



deferred generic class PathPointTool from IntWalk 
    (PathPoint as any)

	---Purpose: Template class to describe the necessary ressources 
	--          for a point used as a starting point for a marching
	--          algorithm.
	--          The 'marching algorithm' determines the intersection 
	--          between an implicit surface and a parametrized surface.
	--          these points are necessary on an arc of the surface

uses Pnt from gp,
     Vec from gp,
     Dir2d from gp

raises OutOfRange from Standard,
       UndefinedDerivative from StdFail

is

    Value3d(myclass; PStart: PathPoint)
    
      	---Purpose: Returns the 3d coordinates of the starting point.

    	returns Pnt from gp;


    Value2d(myclass; PStart: PathPoint; U, V: out Real from Standard);
    
	---Purpose: Returns the <U, V> parameters which are associated 
	--          with <P>
	--          it's the parameters which start the marching algorithm


    IsPassingPnt(myclass; PStart: PathPoint)
    
    	---Purpose: Returns True if the point is a point on a non-oriented
    	--          arc, which means that the intersection line does not
    	--          stop at such a point but just go through such a point.
    	--          IsPassingPnt is True when IsOnArc is True 

    	returns Boolean from Standard;


    IsTangent(myclass; PStart: PathPoint )
    
	---Purpose: Returns True if the surfaces are tangent at this point.
	--          IsTangent can be True when IsOnArc is True
	--          if IsPassingPnt is True and IsTangent is True,this point
	--          is a stopped point.

    	returns Boolean from Standard;


    Direction3d(myclass; PStart: PathPoint)
    
        ---Purpose: returns the tangent at the intersection in 3d space
        --          associated to <P>
        --         an exception is raised if IsTangent is true.

    	returns Vec from gp

    	raises UndefinedDerivative from StdFail;


    Direction2d(myclass; PStart: PathPoint)
    
        ---Purpose: returns the tangent at the intersection in the
        --          parametric space of the parametrized surface.This tangent
        --          is associated to the value2d
        --          la tangente a un sens signifiant (indique le sens de chemin
        --          ement)
        --          an exception is raised if IsTangent is true.

    	returns Dir2d from gp

	raises UndefinedDerivative from StdFail;


    Multiplicity(myclass; PStart: PathPoint)
    
    	---Purpose: Returns the multiplicity of the point i-e 
    	--          the number of auxillar parameters associated to the
    	--          point which the principal parameters are given by Value2d 

    	returns Integer from Standard;


    Parameters(myclass; PStart: PathPoint;
               Mult: Integer from Standard;
               U, V: out Real from Standard) 
	       
    	---Purpose: Parametric coordinates associated to the multiplicity.
    	--          An exception is raised if Mult<=0 or Mult>multiplicity.

    	raises OutOfRange from Standard;


end PathPointTool;

