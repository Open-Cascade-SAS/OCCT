-- Created on: 1992-04-30
-- Created by: Remi GILET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package gce

uses gp,
     StdFail

      	--- Level : Public  
      	--  All methods of all  classes will be public.



is

enumeration ErrorType is Done, ConfusedPoints, NegativeRadius, ColinearPoints,
    	    	      IntersectionError, NullAxis, NullAngle, NullRadius,
    	    	      InvertAxis,BadAngle,InvertRadius,NullFocusLength,
    	    	      NullVector,BadEquation;
    	--- Purpose: Indicates the outcome of a construction, i.e.
    	-- whether it is successful or not, as explained below.
    	-- gce_Done: Construction was successful.
    	-- gce_ConfusedPoints: Two points are coincident.
    	-- gce_NegativeRadius: Radius value is negative.
    	-- gce_ColinearPoints: Three points are collinear.
    	-- gce_IntersectionError: Intersection cannot be computed.
    	-- gce_NullAxis: Axis is undefined.
    	-- gce_NullAngle: Angle value is invalid (usually null).
    	-- gce_NullRadius: Radius is null.
    	-- gce_InvertAxis: Axis value is invalid.
    	-- gce_BadAngle: Angle value is invalid.
    	-- gce_InvertRadius: Radius value is incorrect
    	-- (usually with respect to another radius).
    	-- gce_NullFocusLength: Focal distance is null.
    	-- gce_NullVector: Vector is null.
    	-- gce_BadEquation: Coefficients are
    	-- incorrect (applies to the equation of a geometric object).


private deferred class Root;

class MakeDir2d;

class MakeLin2d;
	
class MakeCirc2d;

class MakeHypr2d;

class MakeElips2d;

class MakeParab2d;

---------------------------------------------------------------------------
    --- Constructions of Trsf2d from gp.
---------------------------------------------------------------------------

class MakeTranslation2d;

class MakeMirror2d;

class MakeRotation2d;
 
class MakeScale2d;

---------------------------------------------------------------------------
    --- Constructions of 3d geometrical elements from gp.
---------------------------------------------------------------------------

class MakeDir;

class MakeLin;
	
class MakeCirc;

class MakeHypr;

class MakeElips;

class MakeParab;

---------------------------------------------------------------------------
    --- Constructions of planes from gp.
---------------------------------------------------------------------------

class MakePln;

---------------------------------------------------------------------------
    --- Construction of surfaces from gp.
---------------------------------------------------------------------------

class MakeCylinder;
 
class MakeCone;

---------------------------------------------------------------------------
    --- Constructions of Trsf from gp.
---------------------------------------------------------------------------

class MakeTranslation;

class MakeMirror;

class MakeRotation;
 
class MakeScale;
 
end gce;



