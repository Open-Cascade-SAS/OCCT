-- Created on: 1993-02-03
-- Created by: Gilles DEBARBOUILLE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class RealParameter from Dynamic

inherits

    Parameter from Dynamic
	---Purpose: This  inherited class from Parameter describes all
	--          the parameters, which  are characterized by a real
	--          value.

uses

    OStream from Standard,
    CString from Standard,
    Real    from Standard


is

    Create(aparameter : CString from Standard )
    
    ---Level: Public 
    
    ---Purpose: Creates a RealParameter with <aparameter> as name.
    
    returns mutable RealParameter from Dynamic;

    Create(aparameter : CString from Standard ; avalue : Real from Standard) 
    
    ---Level: Public 
    
    ---Purpose: With  the name  of the Parameter  <aparameter> and the
    --          real <avalue>, creates an instance of RealParameter.
    
    returns mutable RealParameter from Dynamic;
    
    Value(me) returns Real from Standard
    
    ---Level: Public 
    
    ---Purpose: Returns the value of the parameter which is a real.
    
    is static;

    Value (me : mutable ; avalue : Real from Standard)
    
    ---Level: Public 
    
    --- Purpose: Sets the real <avalue> in <me>.

    is static;
    
    Dump(me ; astream : in out OStream from Standard)
    
    ---Level: Internal 
    
    ---Purpose: Useful for debugging.

    is redefined;
    
fields

    thevalue : Real from Standard;

end RealParameter;
