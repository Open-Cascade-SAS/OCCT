-- Created on: 2000-08-15
-- Created by: data exchange team
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Location from XCAFDoc inherits Attribute from TDF

	---Purpose: 

uses
    Location from TopLoc,
    Label from TDF,
    RelocationTable from TDF

is
    Create returns Location from XCAFDoc;
    
    ---Purpose: class methods
    --          =============

    GetID (myclass)   
    	---C++: return const &  
    returns GUID from Standard;

    Set (myclass; label : Label from TDF; Loc : Location from TopLoc)
    ---Purpose: Find, or create, a Location attribute and set it's value
    --          the Location attribute is returned.
    returns Location from XCAFDoc;

    ---Purpose: Location methods
    --          ===============
    
    Set (me : mutable; Loc : Location from TopLoc);
    
    Get (me)
    returns Location from TopLoc;
        ---C++: return const & 

    --IsCaptured(me) returns Boolean;
	---Purpose: Returns True if there is a reference on the same label

    ---Category: methodes de TDF_Attribute
    --           =========================
    
    ID (me)
    	---C++: return const & 
    returns GUID from Standard;

    Restore (me: mutable; With : Attribute from TDF);

    NewEmpty (me)
    returns mutable Attribute from TDF;

    Paste (me; Into : mutable Attribute from TDF;
	       RT   : mutable RelocationTable from TDF);    

--    Dump(me; anOS : in out OStream from Standard)
--    	returns OStream from Standard
--    	is redefined;
--	-C++: return &

fields
    myLocation : Location from TopLoc;
    
end Location;
