-- Created on: 1991-03-28
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



package IntWalk

	---Purpose: This package defines the "walking" (marching) algorithmes
	--          for the intersection between two surfaces.
	--          One of the surfaces is a parametric one.
	--          If the other is an implicit one, the "IWalking" class will
	--          be used.
	--          If both surfaces are parametric, the "PWalking" class will
	--          be used.

        ---Level: Internal
        --
        -- All the methods of the classes of this package are Internal.
	-- 
uses   
     Standard, MMgt, TCollection, TColStd, gp, math, StdFail, IntSurf, IntImp

is

    enumeration StatusDeflection is 
                PasTropGrand, PointConfondu, ArretSurPointPrecedent,
                ArretSurPoint, OK;

-- StepTooGreat, ConfusedPoint, StopOnPreviousPoint, StopOnPoint, OK
		
-- class for definition of ressources on a biparametric surface

    deferred generic class PSurfaceTool;    


-- classes for definition of marching algorithm on a
-- biparametric surface

    deferred generic class PathPointTool;  

    deferred generic class LoopPointTool;  
    
    deferred generic class IWFunction;

    generic class Iterator;
    
    
--class of result objects marching on a biparametric surface

    generic class IWLine;
    
    
--algorithm marching/solution

    generic class IWalking, TheIWLine, SequenceOfIWLine;
    
    imported VectorOfWalkingData;
    ---Purpose: Defines a dynamic vector of work data.
    
    imported VectorOfInteger;
    ---Purpose: Defines a dynamic vector of integer.

    
--algorithm/solution for a marching on intersection between
-- 2 biparametric surfaces

    generic class PWalking, TheInt2S;


end IntWalk;
