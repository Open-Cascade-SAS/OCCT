-- File:	Dynamic_CompositMethod.cdl
-- Created:	Fri Aug 26 10:30:08 1994
-- Author:	Gilles DEBARBOUILLE
--		<gde@watson>
---Copyright:	 Matra Datavision 1994


class CompositMethod from Dynamic

inherits

    MethodDefinition from Dynamic    
	---Purpose: A composite method is  defined as a collection  of
	--          method instances. This collection describes a more
	--          complex    program   or a  network  of  elementary
	--          functions.   The order of  the method instances is
	--          not significant.  It   is  the references to   the
	--          variables  which    define the  signature  of  the
	--          composite  method which  define  the precedence of
	--          one method in relation with another.
   
uses

    OStream from Standard,
    Integer from Standard,
    CString from Standard,
    Method            from Dynamic, 
    SequenceOfMethods from Dynamic


is

    Create(aname : CString from Standard) returns mutable CompositMethod from Dynamic;
    
    ---Level: Advanced 
    
    ---Purpose: Creates a composit method with <aname> as name.
    
    Method(me : mutable ; amethod : Method from Dynamic)
    
    ---Level: Advanced 
    
    ---Purpose: Adds <amethod>, which  is an elementary or  a composit
    --          method to <me>.
    
    is static;
    
    NumberOfMethods(me) returns Integer from Standard
    
    ---Level: Advanced 
    
    ---Purpose: Returns the   number  of methods   referenced  by  the
    --          composit method <me>.
    
    is static;
    
    Method(me ; anindex : Integer from Standard) returns any Method from Dynamic
    
    ---Level: Advanced 
    
    ---Purpose: Returns the method of range <anindex>.
    
    is static;

    Dump(me ; astream : in out OStream from Standard)
    
    ---Level: Internal 
    
    ---Purpose: Useful for debugging.

    is redefined;
    
fields

    thesequenceofmethods : SequenceOfMethods from Dynamic;

end CompositMethod;
