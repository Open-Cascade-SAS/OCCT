-- Created on: 2003-06-04
-- Created by: Galina KULIKOVA
-- Copyright (c) 2003-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class RWDerivedShapeAspect from RWStepRepr

    ---Purpose: Read & Write tool for DerivedShapeAspect

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    DerivedShapeAspect from StepRepr

is
    Create returns RWDerivedShapeAspect from RWStepRepr;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : DerivedShapeAspect from StepRepr);
	---Purpose: Reads DerivedShapeAspect

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: DerivedShapeAspect from StepRepr);
	---Purpose: Writes DerivedShapeAspect

    Share (me; ent : DerivedShapeAspect from StepRepr;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWDerivedShapeAspect;
