-- File:	AIS_ConcentricRelation.cdl
-- Created:	Thu Dec  5 10:28:03 1996
-- Author:	Flore Lantheaume/Odile Olivier
--		<odl@sacadox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1996




class ConcentricRelation from AIS inherits Relation from AIS

	---Purpose: A framework to define a constraint by a relation of
    	-- concentricity between two or more interactive datums.
    	-- The display of this constraint is also defined.
    	-- A plane is used to create an axis along which the
    	-- relation of concentricity can be extended.

uses

    PresentationManager3d from PrsMgr,
    Presentation          from Prs3d,
    Selection             from SelectMgr,
    Shape                 from TopoDS,
    Pnt                   from gp,
    Dir                   from gp,
    Projector             from Prs3d,
    Transformation        from Geom,
    PresentationManager2d from PrsMgr,
    GraphicObject         from Graphic2d ,   
    Plane                 from Geom
    
is
    Create (aFShape     : Shape          from TopoDS;
    	    aSShape     : Shape          from TopoDS;
	    aPlane      : Plane          from Geom)
	 ---Purpose: Constructs the display object for concentric relations
    	 -- between shapes.
    	 -- This object is defined by the two shapes, aFShape
    	 -- and aSShape and the plane aPlane.
    	 -- aPlane is provided to create an axis along which the
    	 -- relation of concentricity can be extended. 
    returns mutable ConcentricRelation from AIS;

    -- Methods from PresentableObject
    
    Compute(me            : mutable;
  	    aPresentationManager: PresentationManager3d from PrsMgr;
    	    aPresentation : mutable Presentation from Prs3d;
    	    aMode         : Integer from Standard= 0) 
    is redefined static private;
    
    Compute(me:mutable;
    	        aProjector: Projector from Prs3d;
                aPresentation: mutable Presentation from Prs3d)
    is redefined static private;     

    Compute(me:mutable;
    	    aPresentationManager: PresentationManager2d from PrsMgr;
            aPresentation: mutable GraphicObject from Graphic2d;
            aMode: Integer from Standard = 0)
    is redefined static private;	        
    
    Compute(me            : mutable;
    	    aProjector    : Projector from Prs3d;
    	    aTrsf         : Transformation from Geom;
	    aPresentation : mutable Presentation from Prs3d)
    is redefined;
	 ---Purpose: computes the presentation according to a point of view
	 --          given by <aProjector>. 
         --          To be Used when the associated degenerated Presentations 
	 --          have been transformed by <aTrsf> which is not a Pure
	 --          Translation. The HLR Prs can't be deducted automatically
	 --          WARNING :<aTrsf> must be applied
	 --           to the object to display before computation  !!!

    ComputeTwoEdgesConcentric(me:mutable;
    	    	    	      aPresentationManager: Presentation from Prs3d)
    is private;	
			      
    ComputeEdgeVertexConcentric(me:mutable;
    	    	    	        aPresentationManager: Presentation from Prs3d)
    is private;	
    
    ComputeTwoVerticesConcentric(me:mutable;
    	    	    	         aPresentationManager: Presentation from Prs3d)
    is private;	
    
    -- Methods from SelectableObject
   
    ComputeSelection(me         : mutable;
    	    	     aSelection : mutable Selection from SelectMgr;
    	    	     aMode      : Integer from Standard)
    is redefined private;
    
fields
    
    myCenter    : Pnt   from gp;
    myRad       : Real  from Standard;
    myDir       : Dir   from gp;
    myPnt       : Pnt   from gp;

end ConcentricRelation;
