-- Created on: 2000-05-10
-- Created by: Andrey BETENEV
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1

class ObjectRole from StepBasic
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity ObjectRole

uses
    HAsciiString from TCollection

is
    Create returns ObjectRole from StepBasic;
	---Purpose: Empty constructor

    Init (me: mutable; aName: HAsciiString from TCollection;
                       hasDescription: Boolean;
                       aDescription: HAsciiString from TCollection);
	---Purpose: Initialize all fields (own and inherited)

    Name (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Name
    SetName (me: mutable; Name: HAsciiString from TCollection);
	---Purpose: Set field Name

    Description (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Description
    SetDescription (me: mutable; Description: HAsciiString from TCollection);
	---Purpose: Set field Description
    HasDescription (me) returns Boolean;
	---Purpose: Returns True if optional field Description is defined

fields
    theName: HAsciiString from TCollection;
    theDescription: HAsciiString from TCollection; -- optional
    defDescription: Boolean; -- flag "is Description defined"

end ObjectRole;
