-- Created on: 1997-04-17
-- Created by: Christophe MARION
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class AreaLimit from HLRBRep inherits TShared from MMgt 

    ---Purpose: The  private  nested class AreaLimit represents   a --
    --          vertex on  the Edge with the  state on the left and --
    --          the right.
	
uses
    Orientation  from TopAbs,
    State        from TopAbs,
    Intersection from HLRAlgo

is

Create(V            : Intersection from HLRAlgo;
       Boundary     : Boolean      from Standard;
       Interference : Boolean      from Standard;
       StateBefore  : State        from TopAbs;
       StateAfter   : State        from TopAbs;
       EdgeBefore   : State        from TopAbs;
       EdgeAfter    : State        from TopAbs)
returns mutable AreaLimit from HLRBRep;
    ---Purpose: The previous and next field are set to NULL.
    
StateBefore(me : mutable; St : State from TopAbs)
is static;

StateAfter(me : mutable; St : State from TopAbs)
is static;

EdgeBefore(me : mutable; St : State from TopAbs)
is static;

EdgeAfter(me : mutable; St : State from TopAbs)
is static;
	
Previous(me : mutable; P : AreaLimit from HLRBRep)
is static;

Next(me : mutable; N : AreaLimit from HLRBRep)
is static;

Vertex(me) returns Intersection from HLRAlgo
    ---C++: return const &
is static;
	    
IsBoundary(me) returns Boolean from Standard
is static;
	
IsInterference(me) returns Boolean from Standard
is static;
	
StateBefore(me) returns State from TopAbs
is static;

StateAfter(me) returns State from TopAbs
is static;
	
EdgeBefore(me) returns State from TopAbs
is static;

EdgeAfter(me) returns State from TopAbs
is static;

Previous(me) returns mutable AreaLimit from HLRBRep
is static;

Next(me) returns mutable AreaLimit from HLRBRep
is static;
	
Clear(me : mutable)
is static;

fields
    myVertex       : Intersection from HLRAlgo;
    myBoundary     : Boolean      from Standard;
    myInterference : Boolean      from Standard;
    myStateBefore  : State        from TopAbs;
    myStateAfter   : State        from TopAbs;
    myEdgeBefore   : State        from TopAbs;
    myEdgeAfter    : State        from TopAbs;
    myPrevious     : AreaLimit    from HLRBRep;
    myNext         : AreaLimit    from HLRBRep;
	
end AreaLimit;
