-- Created on: 1996-12-23
-- Created by: Alexander BRIVIN
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SFRotation from Vrml 

	---Purpose: defines SFRotation type of VRML field types.
    	--          The  4  values  represent  an  axis  of  rotation  followed  by  amount  of 
	--          right-handed  rotation  about  the  that  axis, in  radians. 
is
 
    Create returns SFRotation from Vrml;

    Create ( aRotationX, aRotationY, aRotationZ : Real from Standard;
             anAngle : Real from Standard )   
    returns SFRotation from Vrml;

    SetRotationX ( me : in out; aRotationX : Real from Standard );
    RotationX ( me )  returns Real from Standard;

    SetRotationY ( me : in out; aRotationY : Real from Standard );
    RotationY ( me )  returns Real from Standard;

    SetRotationZ ( me : in out; aRotationZ : Real from Standard );
    RotationZ ( me )  returns Real from Standard;

    SetAngle ( me : in out; anAngle : Real from Standard );
    Angle ( me )  returns  Real from Standard;

fields

    myRotationX : Real from Standard;
    myRotationY : Real from Standard;
    myRotationZ : Real from Standard;
    myAngle     : Real from Standard;

end SFRotation;

