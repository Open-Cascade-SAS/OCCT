-- File:        PresentedItemRepresentation.cdl
-- Created:     Mon Dec  4 12:02:28 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWPresentedItemRepresentation from RWStepVisual

	---Purpose : Read & Write Module for PresentedItemRepresentation

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     PresentedItemRepresentation from StepVisual,
     EntityIterator from Interface

is

	Create returns RWPresentedItemRepresentation;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable PresentedItemRepresentation from StepVisual);

	WriteStep (me; SW : in out StepWriter; ent : PresentedItemRepresentation from StepVisual);

	Share(me; ent : PresentedItemRepresentation from StepVisual; iter : in out EntityIterator);

end RWPresentedItemRepresentation;
