-- File:	IGESGraph_ToolLineFontDefTemplate.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolLineFontDefTemplate  from IGESGraph

    ---Purpose : Tool to work on a LineFontDefTemplate. Called by various
    --           Modules (ReadWriteModule, GeneralModule, SpecificModule)

uses LineFontDefTemplate from IGESGraph,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolLineFontDefTemplate;
    ---Purpose : Returns a ToolLineFontDefTemplate, ready to work


    ReadOwnParams (me; ent : mutable LineFontDefTemplate;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : LineFontDefTemplate;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : LineFontDefTemplate;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a LineFontDefTemplate <ent>, from
    --           its specific (own) parameters

    DirChecker (me; ent : LineFontDefTemplate) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : LineFontDefTemplate;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : LineFontDefTemplate; entto : mutable LineFontDefTemplate;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : LineFontDefTemplate;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolLineFontDefTemplate;
