-- File:	GeomToStep_MakeSphericalSurface.cdl
-- Created:	Mon Jun 14 16:15:22 1993
-- Author:	Martine LANGLOIS
--		<mla@mastox>
---Copyright:	 Matra Datavision 1993

class MakeSphericalSurface from GeomToStep inherits Root from GeomToStep

    ---Purpose: This class implements the mapping between class
    --          SphericalSurface from Geom and the class
    --          SphericalSurface from StepGeom which describes a
    --          spherical_surface from Prostep
  
uses SphericalSurface from Geom,
     SphericalSurface from StepGeom
     
raises NotDone from StdFail
     
is 



Create ( CSurf : SphericalSurface from Geom ) returns MakeSphericalSurface;

Value (me) returns SphericalSurface from StepGeom
    raises NotDone
    is static;
    ---C++: return const&
 
fields

    theSphericalSurface : SphericalSurface from StepGeom;
    	-- The solution from StepGeom
    	
end MakeSphericalSurface;


