-- Created on: 1994-09-19
-- Created by: Gilles DEBARBOUILLE
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

generic class Node from Dynamic (Item as Transient)

	---Purpose: This generic class    is a light  way  to  store a
	--          persistent   homogeneous  collection  of   objects
	--          inside another persistent object.

inherits

    TShared from MMgt
    

is

    Create returns mutable Node from Dynamic;
    
    ---Level: Advanced 
    
    ---Purpose: Returns an empty instance of this class.

    Create(anitem : any Item) returns mutable Node from Dynamic;
    
    ---Level: Advanced 
    
    ---Purpose: Returns an instance  of  this class  initialized  with
    --          <anitem> as object.

    Object(me : mutable ; anitem : any Item)
    
    ---Level: Advanced 
    
    ---Purpose: Sets to <me> the object <anitem>.
    
    is static;
    
    Object(me) returns any Item
    
    ---Level: Advanced 
    
    ---Purpose: Returns the object into <me>.
    
    is static;
    
    Next(me : mutable ; anode : Node from Dynamic)
    
    ---Level: Advanced 
    
    ---Purpose: Links to <me> the node <anode>.
    
    is static;
    
    Next(me) returns any Node from Dynamic
    
    ---Level: Advanced 
    
    ---Purpose: Returns the node linked to <me>.
    
    is static;
    
fields

    thenextnode : Node from Dynamic;
    theitem     : Item;

end Node;



