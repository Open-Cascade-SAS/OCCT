-- Created on: 1993-02-24
-- Created by: Laurent PAINNOT
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ConstraintCouple from AppParCurves
	    ---Purpose: associates an index and a constraint for an object.
    	    -- This couple is used by AppDef_TheVariational when performing approximations.
uses Constraint from AppParCurves

is 

    Create returns ConstraintCouple;
    	---Purpose: returns an indefinite ConstraintCouple.

    Create(TheIndex: Integer; Cons: Constraint)
    	---Purpose: Create a couple the object <Index> will have the 
    	--          constraint <Cons>.

    returns ConstraintCouple;


    Index(me)
    	---Purpose: returns the index of the constraint object.

    returns Integer
    is static;
    

    Constraint(me) 
    	---Purpose: returns the constraint of the object.

    returns Constraint
    is static;
    

    SetIndex(me: in out; TheIndex: Integer)
    	---Purpose: Changes the index of the constraint object.
    
    is static;
    
    
    SetConstraint(me: in out; Cons: Constraint)
    	---Purpose: Changes the constraint of the object.
    
    is static;
    
    
fields

myIndex:      Integer;
myConstraint: Constraint from AppParCurves;

end ConstraintCouple;
