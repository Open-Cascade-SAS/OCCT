-- Created on: 1993-01-21
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Intersection from IntPatch

  ---Purpose: This class provides a generic algorithm to intersect
	--          2 surfaces.

uses
     HVertex         from Adaptor3d,
     HCurve2d        from Adaptor2d,
     HSurface        from Adaptor3d,
     Point           from IntPatch,
     SequenceOfPoint from IntPatch,
     TopolTool       from Adaptor3d,
     SequenceOfLine  from IntPatch,
     Line            from IntPatch,
     SurfaceType     from GeomAbs,
     ListOfPntOn2S   from IntSurf
 
raises NotDone           from StdFail,
       OutOfRange        from Standard,
       DomainError       from Standard,
       ConstructionError from Standard

is
    Create
    
    	returns Intersection from IntPatch;


    Create (S1: HSurface from Adaptor3d; D1: TopolTool from Adaptor3d;
            S2: HSurface from Adaptor3d; D2: TopolTool from Adaptor3d;
            TolArc,TolTang: Real from Standard)
	    
      returns Intersection from IntPatch
	    raises ConstructionError from Standard;

    Create (S1: HSurface from Adaptor3d; D1: TopolTool from Adaptor3d;
            TolArc,TolTang: Real from Standard)
	    
      returns Intersection from IntPatch
      raises ConstructionError from Standard;


    SetTolerances(me       : in out;
                  TolArc   : Real from Standard;
                  TolTang  : Real from Standard;
                  UVMaxStep: Real from Standard;
                  Fleche   : Real from Standard)
		  
      ---Purpose: Set the tolerances used by the algorithms:
      --          --- Implicit   - Parametric  
      --          --- Parametric - Parametric 
      --          --- Implicit   - Implicit 
      --         
      --          TolArc   is  used  to   compute  the intersections
      --          between the restrictions   of  a  surface   and  a
      --          walking line.
      --          
      --          TolTang is used to compute the points on a walking
      --          line, and in geometric algorithms.
      --          
      --          Fleche  is  a  parameter   used in    the  walking
      --          algorithms to provide small curvatures on a line.
      --          
      --          UVMaxStep is  a  parameter   used in  the  walking
      --          algorithms  to    compute the  distance between to
      --          points in their respective parametrtic spaces.
      --
      
      is static;

    Perform (me: in out;
             S1: HSurface from Adaptor3d; D1: TopolTool from Adaptor3d;
             S2: HSurface from Adaptor3d; D2: TopolTool from Adaptor3d;
             TolArc,TolTang: Real from Standard;
             isGeomInt : Boolean from Standard = Standard_True;
             theIsReqToKeepRLine: Boolean from Standard = Standard_False)   	     

      ---Purpose: Flag theIsReqToKeepRLine has been enterred only for
      --          compatibility with TopOpeBRep package. It shall be deleted
      --          after deleting TopOpeBRep.
      --          When intersection result returns IntPatch_RLine and another
      --          IntPatch_Line (not restriction) we (in case of theIsReqToKeepRLine==TRUE)
      --          will always keep both lines even if they are coincided.
             
      raises ConstructionError from Standard    
      is static;
    
      --amv
    Perform ( me: in out;
              S1: HSurface from Adaptor3d; D1: TopolTool from Adaptor3d;
              S2: HSurface from Adaptor3d; D2: TopolTool from Adaptor3d;
              TolArc,TolTang: Real from Standard;
              LOfPnts: in out ListOfPntOn2S from IntSurf;
              RestrictLine: Boolean from Standard = Standard_True;
              isGeomInt : Boolean from Standard = Standard_True)
              
      ---Purpose: If isGeomInt == Standard_False, then method 
      --          Param-Param intersection will be used.
      
      raises ConstructionError from Standard
      is static;

    Perform ( me: in out;
              S1: HSurface from Adaptor3d; D1: TopolTool from Adaptor3d;
              S2: HSurface from Adaptor3d; D2: TopolTool from Adaptor3d;
              U1,V1,U2,V2 : Real from Standard;
              TolArc,TolTang: Real from Standard)
              
      raises ConstructionError from Standard
      is static;

    Perform (me: in out;
             S1: HSurface from Adaptor3d; D1: TopolTool from Adaptor3d;
             TolArc,TolTang: Real from Standard)
      
      raises ConstructionError from Standard
      is static;
  
    ParamParamPerfom( me: in out;
                      S1: HSurface from Adaptor3d; D1: TopolTool from Adaptor3d;
                      S2: HSurface from Adaptor3d; D2: TopolTool from Adaptor3d;
                      TolArc,TolTang: Real from Standard;
                      LOfPnts: in out ListOfPntOn2S from IntSurf;
                      RestrictLine: Boolean from Standard;
                      typs1, typs2: SurfaceType from GeomAbs)

      is private;
      
    GeomGeomPerfom( me: in out;
                    S1: HSurface from Adaptor3d; D1: TopolTool from Adaptor3d;
                    S2: HSurface from Adaptor3d; D2: TopolTool from Adaptor3d;
                    TolArc,TolTang: Real from Standard;
                    LOfPnts: in out ListOfPntOn2S from IntSurf;
                    RestrictLine: Boolean from Standard;
                    typs1, typs2: SurfaceType from GeomAbs;
                    theIsReqToKeepRLine: Boolean from Standard = Standard_False)
                    
      ---Purpose: Flag theIsReqToKeepRLine has been enterred only for
      --          compatibility with TopOpeBRep package. It shall be deleted
      --          after deleting TopOpeBRep.
      --          When intersection result returns IntPatch_RLine and another
      --          IntPatch_Line (not restriction) we (in case of theIsReqToKeepRLine==TRUE)
      --          will always keep both lines even if they are coincided.

      is private;
      
    GeomGeomPerfomTrimSurf( me: in out;
                            S1: HSurface from Adaptor3d; D1: TopolTool from Adaptor3d;
                            S2: HSurface from Adaptor3d; D2: TopolTool from Adaptor3d;
                            TolArc,TolTang: Real from Standard;
                            LOfPnts: in out ListOfPntOn2S from IntSurf;
                            RestrictLine: Boolean from Standard;
                            typs1, typs2: SurfaceType from GeomAbs;
                            theIsReqToKeepRLine: Boolean from Standard = Standard_False)
                            
      ---Purpose: Flag theIsReqToKeepRLine has been enterred only for
      --          compatibility with TopOpeBRep package. It shall be deleted
      --          after deleting TopOpeBRep.
      --          When intersection result returns IntPatch_RLine and another
      --          IntPatch_Line (not restriction) we (in case of theIsReqToKeepRLine==TRUE)
      --          will always keep both lines even if they are coincided.
      
      is private;
                    
    GeomParamPerfom(me: in out;
                    S1: HSurface from Adaptor3d; D1: TopolTool from Adaptor3d;
                    S2: HSurface from Adaptor3d; D2: TopolTool from Adaptor3d;
                    isNotAnalitical: Boolean from Standard;
                    typs1, typs2: SurfaceType from GeomAbs)
      
      is private;
      
    IsDone(me)
    
    	---Purpose: Returns True if the calculus was succesfull.

    	returns Boolean from Standard
      ---C++: inline
      
    	is static;


    IsEmpty(me)
      ---Purpose: Returns true if the is no intersection.
      ---C++: inline
      returns Boolean from Standard
      raises NotDone from StdFail
      is static;


    TangentFaces(me)
      ---Purpose: Returns True if the two patches are considered as
      --          entierly tangent, i-e every restriction arc of one
      --          patch is inside the geometric base of the other patch.
      ---C++: inline
      
      returns Boolean from Standard
      raises NotDone from StdFail
      is static;
      
    OppositeFaces(me)
      ---Purpose: Returns True when the TangentFaces returns True and the
      --          normal vectors evaluated at a point on the first and the
      --          second surface are opposite. 
      --          The exception DomainError is raised if TangentFaces
      --          returns False.
      ---C++: inline

    	returns Boolean from Standard
      raises  NotDone     from StdFail,
              DomainError from Standard
      is static;


    NbPnts(me)
      ---Purpose: Returns the number of "single" points.
      ---C++: inline

    	returns Integer from Standard
    	raises NotDone from StdFail
    	is static;


    Point(me; Index: Integer from Standard)
    
    	---Purpose: Returns the point of range Index.
    	--          An exception is raised if Index<=0 or Index>NbPnt.
      ---C++: return const&
      ---C++: inline

    	returns Point from IntPatch
    	raises  NotDone    from StdFail,
              OutOfRange from Standard

    	is static;


    NbLines(me)
      ---Purpose: Returns the number of intersection lines.
      ---C++: inline
      
      returns Integer from Standard
      raises NotDone from StdFail
      is static;
      
    Line(me; Index: Integer from Standard)
      ---Purpose: Returns the line of range Index.
    	--          An exception is raised if Index<=0 or Index>NbLine.
      ---C++: return const&
      ---C++: inline

    	returns Line from IntPatch
    	raises  NotDone    from StdFail,
              OutOfRange from Standard
              
      is static;
      
    SequenceOfLine(me)
      ---C++: return const&
      
      returns SequenceOfLine from IntPatch
      raises NotDone    from StdFail
      is static;
	
    Dump(me; Mode : Integer from Standard;
             S1   : HSurface from Adaptor3d; D1: TopolTool from Adaptor3d;
             S2   : HSurface from Adaptor3d; D2: TopolTool from Adaptor3d) 
    	---Purpose: Dump of each result line. 
    	---         Mode for more accurate dumps. 
    	--          
    	is static;

fields

    done       : Boolean         from Standard;
    empt       : Boolean         from Standard;
    tgte       : Boolean         from Standard;
    oppo       : Boolean         from Standard;
    spnt       : SequenceOfPoint from IntPatch;
    slin       : SequenceOfLine  from IntPatch;
    myTolArc   : Real from Standard;
    myTolTang  : Real from Standard;
    myUVMaxStep: Real from Standard;
    myFleche   : Real from Standard;
    myIsStartPnt: Boolean from Standard;
    myU1Start  : Real from Standard;
    myV1Start  : Real from Standard;
    myU2Start  : Real from Standard;
    myV2Start  : Real from Standard;

end Intersection;
