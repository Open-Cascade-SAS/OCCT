-- File:	QADBMReflex.cdl
-- Created:	Mon Oct  7 14:55:32 2002
-- Author:	QA Admin
--		<qa@russox>
---Copyright:	 Matra Datavision 2002

package QADBMReflex
     uses Draw,
          TopoDS,
          AIS,
          PrsMgr,
          Prs3d,
          SelectMgr,
	  Quantity,
	  Graphic3d
is

    class OCC749Prs;
    class OCC749PrsUseVertexC;
    class OCC749PrsUseVertex;
    class OCC749PrsUseVertexCABV;
    class OCC749PrsUseVertexABV;
    Commands(DI : in out Interpretor from Draw);
end;
