-- Created on: 1996-04-09
-- Created by: Yves FRICAUD
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Collect from BRepBuilderAPI 

	---Purpose: 

uses
    Shape                     from TopoDS,
    DataMapOfShapeListOfShape from TopTools,
    MapOfShape                from TopTools,
    MakeShape                 from BRepBuilderAPI
    
is

    Create returns Collect from BRepBuilderAPI;
    
    Add  (me : in out; SI  : Shape            from TopoDS  ;
		       MKS : in out MakeShape from BRepBuilderAPI );
    	---Purpose: 
   
    AddGenerated  (me : in out; S   : Shape from TopoDS  ;  
		                 Gen : Shape from TopoDS  );
       ---Purpose:

    AddModif  (me : in out; S      : Shape from TopoDS  ;  
		             Mod    : Shape from TopoDS  ); 
       ---Purpose: 
		   
    Filter     (me : in out; SF : Shape from TopoDS  );
	---Purpose: 

    Modification (me) returns DataMapOfShapeListOfShape from TopTools;
    ---C++: return const &

    Generated    (me) returns DataMapOfShapeListOfShape from TopTools;
    ---C++: return const &
    
    
fields
    myInitialShape : Shape from TopoDS;
    myDeleted      : MapOfShape from TopTools;
    myMod          : DataMapOfShapeListOfShape from TopTools;
    myGen          : DataMapOfShapeListOfShape from TopTools;
end Collect;
