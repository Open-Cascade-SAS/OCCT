-- Created on: 1992-08-26
-- Created by: Remi GILET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MakeLin from gce inherits Root from gce

    ---Purpose : This class implements the following algorithms used 
    --           to create a Lin from gp.
    --           * Create a Lin parallel to another and passing 
    --             through a point.
    --           * Create a Lin passing through 2 points.
    --           * Create a lin from its axis (Ax1 from gp).
    --           * Create a lin from a point and a direction.

uses Pnt  from gp,
     Lin  from gp,
     Ax1  from gp,
     Dir  from gp,
     Real from Standard

raises NotDone from StdFail

is

Create (A1 : Ax1 from gp)  returns MakeLin;
    --- Purpose : Creates a line located along the axis A1.


Create (P : Pnt from gp; 
    	V : Dir from gp) returns MakeLin;
    --- Purpose : 
    --  <P> is the location point (origin) of the line and
    --  <V> is the direction of the line.

Create(Lin    :     Lin from gp;
       Point  :     Pnt from gp) returns MakeLin;
    ---Purpose : Make a Lin from gp <TheLin> parallel to another 
    --           Lin <Lin> and passing through a Pnt <Point>.

Create(P1     :     Pnt from gp;
       P2     :     Pnt from gp) returns MakeLin;
    ---Purpose : Make a Lin from gp <TheLin> passing through 2 
    --           Pnt <P1>,<P2>.
    --           It returns false if <p1> and <P2> are confused.

Value(me) returns Lin from gp
    raises NotDone
    is static;
    ---C++: return const&
    --- Purpose: Returns the constructed line.
    -- Exceptions StdFail_NotDone is raised if no line is constructed.

Operator(me) returns Lin from gp
    is static;
    ---C++: return const&
    ---C++: alias "Standard_EXPORT operator gp_Lin() const;"

fields

    TheLin : Lin from gp;
    --The solution from gp.
    
end MakeLin;
