-- Created on: 1993-03-03
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Update:      fma


package PTopLoc 

	---Purpose: The  PTopLoc     package      describes persistent
	--          structures for 3D local coordinate systems.
	--          
	--          The  class Datum3D describes  an  elementary local
	--          coordinate system.   It is a linear transformation
	--          (Trsf  from  gp).   The  transformation  is  rigid
	--          (Rotation +  Translation).
	--          
	--          The private    class  ItemLocation represents   an
	--          elementary  local   coordinate   system  (Datum3D)
	--          raised to  an Integer power  elevation. It is used
	--          to link coordinate systems in a Location.
	--          
	--          The  class Location  describes a local  coordinate
	--          system.   It   is  a  chain   of  elementary local
	--          coordinate systems raised to power elevations. The
	--          Location keeps track  of how the coordinate system
	--          was built.

uses

    Standard,
    gp

is
    class Datum3D;
    -- inherits Persistent from Standard
	---Purpose: Persistent elementary local coordinate system.
	
    private class ItemLocation;
    -- inherits Persistent from Standard
	---Purpose: Persistent class  used to  implement Locations.
	
    class Location;
    -- inherits Storable from Standard
	---Purpose: Storable composite local coordinate system.

end PTopLoc;
