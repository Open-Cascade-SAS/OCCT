-- Created on: 1999-03-10
-- Created by: data exchange team
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class OrganizationItem from StepAP214 
inherits ApprovalItem from StepAP214
	

uses

	AppliedOrganizationAssignment from StepAP214,   	
    	Approval from StepBasic
is

    Create returns OrganizationItem;
	---Purpose : Returns a OrganizationItem SelectType

    CaseNum (me; ent : Transient) returns Integer is redefined;
	---Purpose: Recognizes a OrganizationItem Kind Entity that is :
    	
    	--        1 -> AppliedOrganizationAssignment
    	--        2 -> Approval  
    	--        3 -> AssemblyComponentUsageSubstitute
	--        4 -> DocumentFile
    	--        5 -> MaterialDesignation
    	--        6 -> MechanicalDesignGeometricPresentationRepresentation
	--        7 -> PresentationArea
    	--        8 -> Product
	--        9 -> ProductDefinition
    	--        10 -> ProductDefinitionFormation
	--        11 -> ProductDefinitionRelationship
	--        12 -> PropertyDefinition
    	--        13 -> ShapeRepresentation
    	--        14 -> SecurityClassification 
	--        0 else
	
    AppliedOrganizationAssignment (me) returns any AppliedOrganizationAssignment;
	---Purpose : returns Value as a AppliedOrganizationAssignment (Null if another type)
	
    Approval (me) returns any Approval;
    	---Purpose : returns Value as a Approval (Null if another type)
	
	
end OrganizationItem;
