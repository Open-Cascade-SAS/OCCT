-- Created on: 1995-01-30
-- Created by: Mister rmi
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class SensitiveCircle from Select2D 
inherits SensitiveEntity from Select2D

	---Purpose: A framework to define sensitive Areas for a Circle
	--           Radius and center, or a geometric circle is given.

uses

    Circ2d from gp,
    TypeOfSelection,
    EntityOwner from SelectBasics,
    ListOfBox2d from SelectBasics
is

    Create (OwnerId      : EntityOwner from SelectBasics;
    	    TheCirc      : Circ2d from gp;
    	    TheType      : TypeOfSelection = Select2D_TOS_BOUNDARY)
    returns mutable SensitiveCircle ;
    	--- Purpose: Constructs a sensitive circle object defined by the
    	-- owner OwnerId, the circle Circle, and the selection type Type.
    	-- Type can be:
    	-- -   interior
    	-- -   boundary.   
    
    Areas (me:mutable ; aresul : in out ListOfBox2d from SelectBasics) is static;
    	---Level: Public 
    	---Purpose: returns the sensitive areas for a circle...    
    
    Matches (me  : mutable ;
             X,Y : Real from Standard;
             aTol: Real from Standard;
             DMin: out Real from Standard) 
    returns Boolean is static;     
    	---Purpose: Returns true if the minimum distance DMin
    	--          between the postion x,y and the circle is less than aTol..

    Matches (me  :mutable; 
             XMin,YMin,XMax,YMax : Real from Standard;
             aTol: Real from Standard) 
    returns Boolean
    is static;
		     


    Circle(me) returns Circ2d from gp;
    	---Purpose: Returns the circle used at the time of construction of this object.
        ---C++: inline
        ---C++: return const&

    SetTypeOfSelection(me:mutable;aType : TypeOfSelection);
    	---Purpose: Sets the selection type.
        ---C++: inline

    Selection(me:mutable) returns TypeOfSelection from Select2D;
    	---Purpose: Returns the selection type used at the time of construction of this object.
        ---C++: inline

fields

    myCirc  : Circ2d from gp;
    mytype  : TypeOfSelection;   

end SensitiveCircle;
