-- Created on: 1995-10-19
-- Created by: Andre LIEUTIER
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class PinpointConstraint from Plate
---Purpose : define a constraint on the Plate
--         

uses 
   XY from gp, 
   XYZ from gp

is
    Create returns PinpointConstraint;
    Create(point2d : XY ; ImposedValue : XYZ ;
           iu : Integer = 0; iv : Integer = 0) returns PinpointConstraint;

     -- Accessors :
    Pnt2d(me) returns XY from gp;
    ---C++: inline 
    ---C++: return const  &
    
    Idu(me) returns  Integer;
    ---C++: inline
    ---C++: return const &
    
    Idv(me) returns Integer;
    ---C++: inline
    ---C++: return const &
    
    Value(me) returns XYZ from gp;
    ---C++: inline
    ---C++: return const &
  
fields
    
    value : XYZ ;  
    pnt2d : XY ; 
    idu,idv : Integer;
   
end;
