-- Created on: 1992-09-30
-- Created by: Gilles DEBARBOUILLE
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Bisector from MAT

	---Purpose:

inherits

    TShared from MMgt

uses

    ListOfBisector from MAT,
    Edge from MAT

is

    Create

    ---Purpose:

    returns mutable Bisector from MAT;
    
    AddBisector(me ; abisector : any Bisector from MAT)
    
    is static;
    
    List(me) returns any ListOfBisector from MAT
    
    is static;
    
    FirstBisector(me) returns any Bisector from MAT
    
    is static;

    LastBisector(me) returns any Bisector from MAT
    
    is static;

    BisectorNumber(me : mutable ; anumber : Integer)
    
    is static;
    
    IndexNumber(me : mutable ; anumber : Integer)
    
    is static;
    
    FirstEdge(me : mutable ; anedge : any Edge from MAT)
    
    is static;
    
    SecondEdge(me : mutable ; anedge : any Edge from MAT)
    
    is static;
    
    IssuePoint(me : mutable ; apoint : Integer)
    
    is static;
    
    EndPoint(me : mutable ; apoint : Integer)
    
    is static;

    DistIssuePoint(me : mutable ; areal : Real)
    
    is static;
    
    FirstVector(me : mutable ; avector : Integer)
    
    is static;
    
    SecondVector(me : mutable ; avector : Integer)
    
    is static;
    
    Sense(me : mutable ; asense : Real)
    
    is static;
    
    FirstParameter(me : mutable ; aparameter : Real)
    
    is static;
    
    SecondParameter(me : mutable ; aparameter : Real)
    
    is static;
    
    BisectorNumber(me) returns Integer
    
    is static;
    
    IndexNumber(me) returns Integer
    
    is static;
    
    FirstEdge(me) returns any Edge from MAT
    
    is static;
    
    SecondEdge(me) returns any Edge from MAT
    
    is static;
    
    IssuePoint(me) returns Integer
    
    is static;
    
    EndPoint(me) returns Integer
    
    is static;

    DistIssuePoint(me) returns Real
    
    is static;
			    
    FirstVector(me) returns Integer
    
    is static;
    
    SecondVector(me) returns Integer
    
    is static;
    
    Sense(me) returns Real
    
    is static;
    
    FirstParameter(me) returns Real
    
    is static;
    
    SecondParameter(me) returns Real
    
    is static;
    
    Dump(me ; ashift , alevel : Integer)
    
    is static;
    
fields

    thebisectornumber  : Integer;
    theindexnumber     : Integer;
    thefirstedge       : Edge from MAT;
    thesecondedge      : Edge from MAT;
    thelistofbisectors : ListOfBisector from MAT;
    theissuepoint      : Integer;
    theendpoint        : Integer;
    thefirstvector     : Integer;
    thesecondvector    : Integer;
    thesense           : Real;
    thefirstparameter  : Real;
    thesecondparameter : Real;
    distissuepoint     : Real;
end Bisector;
