-- Created on: 1992-03-06
-- Created by: Isabelle GRIGNON
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred generic class PSurfaceTool from IntImp
    (Surface as any)          
                                   

	---Purpose: Template class for a tool on a bi-parametrised surface.
	--          It is possible to implement this tool with an
	--          instantiation of the SurfaceTool from Adaptor3d.

uses Pnt from gp,
     Vec from gp
 
is

    UIntervalFirst(myclass ; S: Surface)
	   
	---Purpose: Returns the first U parameter of the surface.

    	returns Real from Standard;
    
    
    VIntervalFirst(myclass ; S: Surface)
	   
	---Purpose: Returns the first V parameter of the surface.

    	returns Real from Standard;
    
    
    UIntervalLast(myclass ; S: Surface)
	   
	---Purpose: Returns the last U parameter of the surface.

    	returns Real from Standard;
    
    
    VIntervalLast(myclass ; S: Surface)
	   
	---Purpose: Returns the last V parameter of the surface.

    	returns Real from Standard;
    
    
    Value (myclass ; S: Surface; U,V : Real from Standard)
    
    	---Purpose: Returns the point of parameter (U,V) on the surface.

    	returns Pnt from gp;


    D1(myclass; S: Surface; U,V: Real from Standard; 
                P: out Pnt from gp; D1U,D1V: out Vec from gp);
		
	---Purpose: Returns the point of parameter (U,V) on the surface,
	--          and the first derivatives in the directions u and v.

    
    UResolution(myclass; S : Surface; Tol3d: Real from Standard)
    
	---Purpose: Returns the numerical resolution in the U direction,
	--          for a given resolution in 3d space.

    	returns Real from Standard;


    VResolution(myclass; S : Surface; Tol3d: Real from Standard)
    
	---Purpose: Returns the numerical resolution in the V direction,
	--          for a given resolution in 3d space.

    	returns Real from Standard;


end PSurfaceTool;
