-- Created on: 1992-10-13
-- Created by: Ramin BARRETO
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class StackManager from MMgt
---Purpose:
--   The class <StackManager> provides primitive facilities for managing
--   stack-based storage.
--   

uses 
    Integer from Standard
   ,Address from Standard

raises
    OutOfMemory from Standard
   ,ProgramError from Standard

is
    Create returns StackManager;
    ---Purpose:
    --   Constructs a StackManager with an empty free stack.
    --
    ---Level: Advanced
    
    Allocate(me: in out; size: Integer) returns Address
    ---Purpose:
    --   Returns the address of a storage of the given size located on
    --   the top of the free stack.
    ---Level: Advanced
    raises OutOfMemory 
    	   -- If the allocation fails
    is static;
    
    Free(me: in out; aStack: in out Address; aSize: Integer)
    ---Purpose:
    --   Deallocates the storage of the given size from the free stack
    --   and nullify the address.
    ---Level: Advanced
    raises ProgramError  
    	   -- If the storage is not on the top of the stack.
    is static;
    
    ShallowCopy (me) returns StackManager;
    ---Purpose: 
    --   There is no way to have a "ShallowCopy" of a "StackManager"
    ---Level: Advanced
    ---Warning:
    --   A ProgramError will be raised with a message.
    --   
    ---C++:  function call

    Purge(me: in out)
    ---Purpose:
    --   Deallocates the storage associated to stack.
    ---Level: Advanced
    is static private;
    
    ShallowDump (me; S: in out OStream);
    ---Purpose: 
    --   Prints the contents of <me> on the stream <s>. 
    ---Level: Advanced
    ---C++:  function call

    Destructor(me: in out);
    ---Purpose:
    --    Deallocates the storage associated to stack.
    --    Delete <me>.
    ---Level: Advanced
    ---C++: alias ~
    
fields
    myFreeListSize: Integer;
    myFreeList:     Address;

end StackManager;
    
