-- Created on: 1999-11-09
-- Created by: data exchange team
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package StepAP203 

    ---Purpose: Contains implementation of STEP entities specific for AP203

uses
    TCollection,
    StepBasic,
    StepRepr

is

    class ApprovedItem;
    class CcDesignApproval;
    class CcDesignCertification;
    class CcDesignContract;
    class CcDesignDateAndTimeAssignment;
    class CcDesignPersonAndOrganizationAssignment;
    class CcDesignSecurityClassification;
    class CcDesignSpecificationReference;
    class CertifiedItem;
    class Change;
    class ChangeRequest;
    class ChangeRequestItem;
    class ClassifiedItem;
    class ContractedItem;
    class DateTimeItem;
    class PersonOrganizationItem;
    class SpecifiedItem;
    class StartRequest;
    class StartRequestItem;
    class StartWork;
    class WorkItem;

    imported Array1OfApprovedItem;
    imported transient class HArray1OfApprovedItem;

    imported Array1OfCertifiedItem;
    imported transient class HArray1OfCertifiedItem;

    imported Array1OfClassifiedItem;
    imported transient class HArray1OfClassifiedItem;

    imported Array1OfContractedItem;
    imported transient class HArray1OfContractedItem;

    imported Array1OfDateTimeItem;
    imported transient class HArray1OfDateTimeItem;

    imported Array1OfPersonOrganizationItem;
    imported transient class HArray1OfPersonOrganizationItem;

    imported Array1OfSpecifiedItem;
    imported transient class HArray1OfSpecifiedItem;

    imported Array1OfWorkItem;
    imported transient class HArray1OfWorkItem;

    imported Array1OfChangeRequestItem;
    imported transient class HArray1OfChangeRequestItem;

    imported Array1OfStartRequestItem;
    imported transient class HArray1OfStartRequestItem;

end StepAP203;
