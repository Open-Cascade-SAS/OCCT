-- Created on: 2002-04-10
-- Created by: QA Admin
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class  MyText  from  QABugs  inherits  InteractiveObject  from  AIS 
uses 
    ExtendedString from TCollection, 
    Pnt from gp, 
    PresentationManager3d from PrsMgr, 
    Presentation from Prs3d,
    NameOfColor  from  Quantity,
    Selection from SelectMgr
is 
    Create(aText  :ExtendedString  from  TCollection;aPosition  : Pnt  from  gp)
    returns mutable MyText from QABugs;
    Create(aText  :ExtendedString  from  TCollection;aPosition  : Pnt  from  gp;aFont :  CString from Standard; aColor : NameOfColor  from  Quantity; aHeight :Real  from  Standard)
    returns mutable MyText from QABugs;

    NbPossibleSelection(me)
    returns Integer from Standard
    is redefined virtual protected;
    
    Compute(me:mutable;
            aPresentationManager: PresentationManager3d from PrsMgr;
            aPresentation: mutable Presentation from Prs3d;
            aMode: Integer from Standard = 0)
    is redefined virtual protected;

    ComputeSelection(me:mutable; aSelection :mutable Selection from SelectMgr;
                                 aMode      : Integer) is redefined virtual protected;

fields
        myPosition                   : Pnt from gp;
        myText                       : ExtendedString from TCollection;
        myNameOfColor                : NameOfColor from Quantity;
        myNameOfFont                 : CString from Standard;
        myHeight                     : Real from Standard;
end MyText;
    
