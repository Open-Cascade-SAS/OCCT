-- Created on: 2000-08-17
-- Created by: Vincent DELOS
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class AncestorsSeqAndSuccessorsSeq from BooleanOperations 

	---Purpose: provide all the ancestors and  successors of a --
	--          given shape.  Exemple : for  an edge the ancestors
	--           -- are the wires  that hold it and the successors
	--          are -- its vertices.  As  we don't know the number
	--          of -- ancestors of a given shape we first put them
	--           in a -- sequence  of integers (our data structure
	--          -- defining      the shapes does not   have   back
	--          pointers). Then  we   transfer these data  in  the
	--          class AncestorsAndSuccessors.

uses
    Orientation from TopAbs,
    SequenceOfInteger from TColStd,
    AncestorsAndSuccessors from BooleanOperations

is

    Create returns AncestorsSeqAndSuccessorsSeq from BooleanOperations;

      
    Dump (me);
    ---Purpose: to display the fields.


    --------------------
    -- INLINE METHODS --
    --------------------

    GetAncestor   (me; AncestorIndex:    Integer) returns Integer;
    ---C++: inline    
    GetSuccessor  (me; SuccessorIndex:   Integer) returns Integer;
    ---C++: inline    
    GetOrientation(me; OrientationIndex: Integer) returns Orientation;
    ---C++: inline    

    NumberOfAncestors  (me) returns Integer;
    ---C++: inline
    NumberOfSuccessors (me) returns Integer;
    ---C++: inline

    SetNewAncestor   (me:in out; AncestorNumber: Integer);
    ---C++: inline    
    ---Purpose: appends AncestorNumber in the sequence.
    SetNewSuccessor  (me:in out; SuccessorNumber: Integer);
    ---C++:   inline
    ---Purpose: appends SuccessorNumber in the array refering to <mySuccessorsInserted>.
    SetNewOrientation(me:in out; theOrientation: Orientation);
    ---C++:   inline
    ---Purpose: appends SuccessorNumber in the array refering to <mySuccessorsInserted>.


fields

myAncestors: SequenceOfInteger;
---Purpose: the sequence containing all the ancestors of our given shape.

mySuccessors: SequenceOfInteger;
---Purpose: the array containing all the successors.

myOrientations:SequenceOfInteger;
---Purpose: the array containing all orientations corresponding to the successors.

end AncestorsSeqAndSuccessorsSeq;
