-- Created on: 1991-01-23
-- Created by: Christophe MARION
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class Datum3D from TopLoc inherits TShared from MMgt

	---Purpose: Describes a coordinate transformation, i.e. a change
-- to an elementary 3D coordinate system, or position in 3D space.
-- A Datum3D is always described relative to the default datum.
-- The default datum is described relative to itself: its
-- origin is (0,0,0), and its axes are (1,0,0) (0,1,0) (0,0,1).

uses
    Trsf   from gp

raises
    ConstructionError from Standard
    
is
    Create returns mutable Datum3D;
    	---Purpose: Constructs a default Datum3D.

    Create(T : Trsf from gp) returns mutable Datum3D from TopLoc
	---Purpose: Constructs a Datum3D form a Trsf from gp. An error is
	--          raised if the Trsf is not a rigid transformation.
    raises 
    	ConstructionError from Standard;
    
    Transformation(me) returns Trsf from gp
    	---Purpose: Returns a gp_Trsf which, when applied to this datum,
    	-- produces the default datum.
    	---C++: inline
    	---C++: return const &
    	is static;
    
    ShallowDump(me; S : in out OStream);
	--- Purpose:
    	-- Writes the contents of this Datum3D to the stream S.
	---C++: function call

fields

    myTrsf : Trsf from gp;

end Datum3D;
