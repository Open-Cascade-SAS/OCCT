-- Created on: 1996-07-05
-- Created by: Design
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

schema ShapeSchema

is


---Category: inheritage and persistence basic tools

    package ObjMgt;

    package PTopLoc;
    package PColgp;
    package PGeom2d;
    package PGeom;
    package PColPGeom;
    package PColPGeom2d;
    package PPoly;
    package PTopoDS;
    package PBRep;

    package PCDMShape; -- class Document from PCDM.

end ShapeSchema;
