-- Created on: 1996-07-24
-- Created by: Herve LOUESSARD
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package LocalAnalysis  

    ---Purpose:
    -- This package gives tools to check the local continuity 
    -- between two  points situated  on two curves or two surfaces. 

uses

    Standard,
    StdFail,
    LProp,
    GeomAbs,
    Geom,
    Geom2d,
    GeomLProp,
    gp
    
is


--  enumeration used to describe the  status error 
   
enumeration  StatusErrorType   is  NullFirstDerivative, NullSecondDerivative, 
                                 TangentNotDefined,NormalNotDefined,
                                 CurvatureNotDefined         
end  StatusErrorType; 

     
    class SurfaceContinuity;

    class CurveContinuity; 
    ---Purpose:
    -- This  class  compute
    -- s  and gives  tools to check  the  local
    -- continuity  between two points situated  on 2  curves) 
    
    
    
   
    Dump( surfconti : SurfaceContinuity from LocalAnalysis;
          o: in out OStream);	
    ---Purpose:
    -- This fonction gives informations  about a  variable CurveContinuity
	  
    Dump( curvconti : CurveContinuity from LocalAnalysis;
          o: in out OStream);	
    ---Purpose:
    -- This fonction gives informations  about a variable SurfaceContinuity 
	  
    	  	  
end LocalAnalysis; 




















