-- Created on: 2014-03-15
-- Created by: Laurent PAINNOT
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class NewtonFunctionRoot from math 
     ---Purpose:
     -- This class implements the calculation of a root of a function of
     -- a single variable starting from an initial near guess using the
     -- Newton algorithm. Knowledge of the derivative is required.


uses Vector from math, Matrix from math,
     FunctionWithDerivative from math,
     OStream from Standard
     
raises NotDone from StdFail

is 

    Create(F: in out FunctionWithDerivative;
    	   Guess, EpsX, EpsF: Real;
	   NbIterations: Integer = 100)
    ---Purpose:
    -- The Newton method is done to find the root of the function F 
    -- from the initial guess Guess.
    -- The tolerance required on the root is given by Tolerance.
    -- The solution is found when :
    --  abs(Xi - Xi-1) <= EpsX and abs(F(Xi))<= EpsF
    -- The maximum number of iterations allowed is given by NbIterations.
    returns NewtonFunctionRoot;


    Create(F: in out FunctionWithDerivative;
    	   Guess, EpsX, EpsF, A, B: Real;
	   NbIterations: Integer = 100)
    ---Purpose:
    -- The Newton method is done to find the root of the function F 
    -- from the initial guess Guess.
    -- The solution must be inside the interval [A, B].
    -- The tolerance required on the root is given by Tolerance.
    -- The solution is found when :
    --  abs(Xi - Xi-1) <= EpsX and abs(F(Xi))<= EpsF
    -- The maximum number of iterations allowed is given by NbIterations.
    returns NewtonFunctionRoot;


    Create(A, B, EpsX, EpsF: Real; 
           NbIterations: Integer = 100)
        ---Purpose: is used in a sub-class to initialize correctly all the fields
        --          of this class.

    returns NewtonFunctionRoot;
    

    Perform(me: in out; F: in out FunctionWithDerivative;
    	    Guess: Real)
        ---Purpose: is used internally by the constructors.

    is static;


    IsDone(me)
    	---Purpose: Returns true if the computations are successful, otherwise returns false.
      	---C++: inline
  returns Boolean
    is static;
    
    
    Root(me)
    	---Purpose: Returns the value of the root of function <F>.
        -- Exception NotDone is raised if the root was not found.
    	---C++: inline

    returns Real
    raises NotDone
    is static;
    

    Derivative(me)
    	---Purpose: returns the value of the derivative at the root.
        -- Exception NotDone is raised if the root was not found.
    	---C++: inline
    returns Real
    raises NotDone
    is static;
    

    Value(me)
    	---Purpose: returns the value of the function at the root.
        -- Exception NotDone is raised if the root was not found.
    	---C++: inline
    returns Real
    raises NotDone
    is static;
    

    NbIterations(me)
        ---Purpose: Returns the number of iterations really done on the 
        -- computation of the Root.
        -- Exception NotDone is raised if the root was not found.
    	---C++: inline
    returns Integer
    raises NotDone
    is static;


    Dump(me; o:in out OStream)
    	---Purpose: Prints information on the current state of the object.

    is static;


fields

Done: Boolean;
X   : Real;
Fx  : Real;
DFx : Real;
It  : Integer;
EpsilonX: Real;
EpsilonF: Real;
Itermax: Integer;
Binf: Real;
Bsup: Real;

end NewtonFunctionRoot;

