-- Created on: 1997-03-28
-- Created by: Christian CAILLET
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class MeasureValueMember  from StepBasic    inherits  SelectReal  from StepData

    ---Purpose : for Select MeasureValue, i.e. :
    --         length_measure,time_measure,plane_angle_measure,
    --         solid_angle_measure,ratio_measure,parameter_value,
    --         context_dependent_measure,positive_length_measure,
    --         positive_plane_angle_measure,positive_ratio_measure,
    --	       area_measure,volume_measure

uses CString

is

    Create returns mutable MeasureValueMember;
    -- starts as case null (no name)

    HasName (me) returns Boolean  is redefined;
    -- returns True is case not null

    Name    (me) returns CString  is redefined;
    --  returns a name according to the case
    --  0 -> void
    --  1 -> LENGTH_MEASURE
    --  2 -> TIME_MEASURE
    --  3 -> PLANE_ANGLE_MEASURE
    --  4 -> SOLID_ANGLE_MEASURE
    --  5 -> RATIO_MEASURE
    --  6 -> PARAMETER_VALUE
    --  7 -> CONTEXT_DEPENDANT_MEASURE
    --  8 -> POSITIVE_LENGTH_MEASURE
    --  9 -> POSITIVE_PLANE_ANGLE_MEASURE
    --  10 -> POSITIVE_RATIO_MEASURE
    --  11 -> AREA_MEASURE
    --  12 ->VOLUME_MEASURE
    --  13 ->MASS_MEASURE
    --  14 ->THERMODYNAMIC_TEMPERATURE_MEASURE
    
    SetName (me : mutable; name : CString)  returns Boolean  is redefined;
    -- checks for one of the names above, and sets the case number
    -- accepts a void name (case 0)

fields

    thecase : Integer;

end MeasureValueMember;
