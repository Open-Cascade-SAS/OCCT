-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class EventManager from Viewer2dTest inherits TShared from MMgt

	---Purpose: 

uses
    View from V2d,
    InteractiveContext from AIS2D

is

    Create(aCtx:InteractiveContext from AIS2D)
    returns mutable EventManager from Viewer2dTest;

    MoveTo(me:mutable; xpix,ypix:Integer;aView:View from V2d) is virtual;

    Select(me:mutable) is virtual;

    ShiftSelect(me:mutable) is virtual;

    Select(me:mutable;xmin,ymin,xmax,ymax:Integer;aView:View from V2d) is virtual;

    ShiftSelect(me:mutable;xmin,ymin,xmax,ymax:Integer;aView:View from V2d) is virtual;

    Context(me) returns InteractiveContext from AIS2D;
    ---C++: return const&

fields

    myCtx : InteractiveContext from AIS2D;

end EventManager;
