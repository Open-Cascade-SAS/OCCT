-- Created on: 1994-03-30
-- Created by: Laurent BUCHARD
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SolidClassifier from BRepClass3d  inherits SClassifier from BRepClass3d
     
     ---Purpose: Provides an algorithm to classify a point in a solid.



uses 
    Pnt           from gp,
    Face          from TopoDS,
    Shape         from TopoDS,
    SolidExplorer from BRepClass3d

raises

    DomainError from Standard
	
is 


    Create
    	---Purpose : empty constructor
    returns SolidClassifier from BRepClass3d;
        
    Load(me:in out; S   :        Shape from TopoDS)
    is static;
    

    Create(S   :        Shape from TopoDS)
    	---Purpose: Constructor from a Shape.
    returns SolidClassifier from BRepClass3d;
    
    
    Create(S   :        Shape from TopoDS; 
           P   :        Pnt from gp;
	   Tol :        Real from Standard)
    	---Purpose: Constructor to classify the point P with the 
    	--          tolerance Tol on the solid S.
    returns SolidClassifier from BRepClass3d;
    

    Perform(me: in out;
            P   :        Pnt from gp;
	    Tol :        Real from Standard)
    	---Purpose: Classify the point P with the 
    	--          tolerance Tol on the solid S.
    is static;

    PerformInfinitePoint(me: in out;
			 Tol :        Real from Standard)
    	---Purpose: Classify an infinite point with the 
    	--          tolerance Tol on the solid S.
    	--          Useful for compute the orientation of a solid. 
    is static;
    
    Destroy(me:in out)
    	---C++: alias ~
    is static;
    

fields
    aSolidLoaded   : Boolean       from Standard;
    explorer       : SolidExplorer from BRepClass3d;
    isaholeinspace : Boolean       from Standard;
end SolidClassifier;
