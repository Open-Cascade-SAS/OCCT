-- Created on: 1999-11-05
-- Created by: Vladislav ROMASHKO
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Revol from QANewBRepNaming inherits TopNaming from QANewBRepNaming 

    ---Purpose: To load the Revol results 

uses 
 
    MakeRevol from BRepPrimAPI, 
    Shape     from TopoDS,
    Label     from TDF

is 
 
    Create returns Revol from QANewBRepNaming;

    Create(ResultLabel : Label from TDF) 
    returns Revol from QANewBRepNaming;

    Init(me : in out; ResultLabel : Label from TDF);


    Load (me; mkRevol : in out MakeRevol from BRepPrimAPI;
	      basis   : in     Shape     from TopoDS);
    ---Purpose: Loads the revol in the data framework 
      
    Start(me)
    ---Purpose: Returns the insertion label of the start face of the Revol.  
    returns Label from TDF;

    End(me) 
    ---Purpose: Returns the insertion label of the end face of the Revol. 
    returns Label from TDF;
       
    Lateral(me) 
    ---Purpose: Returns the insertion label of the lateral faces of the Revol.
    returns Label from TDF; 
    
    Degenerated(me)
    ---Purpose: Returns the label of degenerated edges.
    returns Label from TDF;
    
    Content(me)
    ---Purpose: Returns the label of the content of the result.
    returns Label from TDF;    
    

end Revol;
