-- Created on: 1991-09-05
-- Created by: Philippe COICADAN
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Revised      J.P. TIRAULT
--              New organization of standard Package (August 1992)


class Failure from Standard inherits Transient from Standard 

    ---Purpose: 
    --   Forms the root of the entire exception hierarchy.

uses
    CString from Standard,
    OStream from Standard,
    SStream from Standard

raises
    NoSuchObject from Standard
    
is

    Create returns mutable Failure;
    	---Purpose: 
    	--   Creates a status object of type "Failure".
    	---Level: Advanced
	---C++: alias "Standard_EXPORT Standard_Failure (const Standard_Failure& f);"

    Create (aString: CString) returns mutable Failure;
    	---Purpose: 
    	--   Creates a status object of type "Failure".
        ---Level: Advanced
      	---C++: alias "Standard_EXPORT Standard_Failure& operator= (const Standard_Failure& f);"

    Destroy(me:mutable);
    	---Level: Advanced
      	---C++: alias ~

    Print (me; s: in out OStream);
    	---Purpose: 
    	--   Prints on the stream <s> the exception name followed by 
    	--   the error message.
        --  Level: Advanced
    	--  Warning:
    	--   The operator "OStream& operator<< (Standard_OStream&,
    	--                                      Handle(Standard_Failure)&)"
    	--   is implemented. (This operator uses the method Print)
    	--   
   	---C++: alias operator<< 

    GetMessageString (me) returns CString from Standard;
        ---Purpose: Returns error message
        ---C++: inline
    
    SetMessageString (me: mutable; aMessage: CString);
    	---Purpose: Sets error message

    Reraise (me: mutable);
    Reraise (me: mutable; aMessage: CString);
    Reraise (me: mutable; aReason: SStream);
    	---Purpose: Reraises a caught exception and changes its error message.
        ---Level: Advanced
    
    Raise (myclass; aMessage: CString  = "") ;
    	---Purpose: Raises an exception of type "Failure" and associates
    	--          an error message to it. The message can be printed 
    	--          in an exception handler.
        ---Level: Advanced
	
        
    Raise (myclass; aReason: SStream) ;
    	---Purpose: Raises an exception of type "Failure" and associates
    	--          an error message to it. The message can be constructed
    	--          at run-time.
        ---Level: Advanced
    
    NewInstance(myclass; aMessage: CString) returns mutable Failure;
   	---Purpose: Used to construct an instance of the exception object
	--          as a handle. Shall be used to protect against possible
	--          construction of exception object in C stack -- that is 
	--          dangerous since some of methods require that object
	--          was allocated dynamically.
	
    Jump (me);
   	---Purpose: Used to throw CASCADE exception from C signal handler.
        --          On platforms that do not allow throwing C++ exceptions 
        --          from this handler (e.g. Linux), uses longjump to get to 
        --          the current active signal handler, and only then is 
        --          converted to C++ exception.
        ---Level: Advanced, not for regular use
    
    Caught (myclass) returns mutable Failure raises NoSuchObject;
    	---Purpose: Returns the last caught exception. 
	--          Needed when exceptions are emulated by C longjumps,
        --          in other cases is also provided for compatibility.

    Throw (me) is virtual protected;
	---Purpose: Used only if standard C++ exceptions are used.
	--          Throws exception of the same type as this by C++ throw,
	--          and stores current object as last thrown exception,
	--          to be accessible by method Caught()

fields
    
    myMessage: CString;
    
end Failure from Standard;

