-- Created on: 1995-01-13
-- Created by: GG
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MarkerStyle from Aspect

	---Version:

	---Purpose: This class defines a Marker Style.
	--	    The Style can be Predefined or defined by the user
	--	    A user defined style must be described in the space <-1,+1>

	---Keywords: MarkerStyle 

	---Warning:
	---References:

uses
	TypeOfMarker from Aspect,
	Array1OfReal from TColStd,
	Array1OfBoolean from TColStd,
	HArray1OfBoolean from TColStd,
	Array1OfShortReal from TShort,
	HArray1OfShortReal from TShort

raises
	MarkerStyleDefinitionError from Aspect

is
	Create returns MarkerStyle from Aspect;
	---Level: Public
	---Purpose: Creates a marker style with the default value of
	--	    MarkerStyle type : POINT
	--

	Create ( aType	: TypeOfMarker ) returns MarkerStyle from Aspect ;
	---Level: Public
	---Purpose: Creates the marker style <aType>.

	Create ( aXpoint : Array1OfReal ; 
	         aYpoint : Array1OfReal ) 
					returns MarkerStyle from Aspect
	---Level: Public
	---Purpose: Creates a marker style from a implicit draw point 
	--descriptor .
	-- Each coordinate <aXpoint(i),aYpoint(i)> must be defined 
	--in the space -1,+1.
	raises MarkerStyleDefinitionError;
	---Trigger:
	-- if <aXpoint>,<aYpoint> have different length.
	-- if one coordinate is <-1 or >+1.

	Create ( aXpoint : Array1OfReal ; 
	         aYpoint : Array1OfReal ; 
	  	 aSpoint : Array1OfBoolean )
					returns MarkerStyle from Aspect
	---Level: Public
	---Purpose: Creates a marker style from a move-draw point descriptor .
	-- Each coordinate <aXpoint(i),aYpoint(i)> must be defined 
	--in the space -1,+1.
	-- Each status point <aSpoint(i)> must be TRUE for drawing
	--or FALSE for moving to the last at this point .
	raises MarkerStyleDefinitionError;
	---Trigger:
	-- if <aXpoint>,<aYpoint>,<aSpoint> have different length.
	-- if one coordinate is <-1 or >+1

        ---------------------------------------------------
        -- Category: Methods to modify the class definition
        ---------------------------------------------------
 
        Assign ( me     : in out ;
                 Other  : MarkerStyle from Aspect )
                returns MarkerStyle from Aspect is static;
        ---Level: Public
        ---Purpose: Updates the marker style <me> from the definition of the
        --          marker style <Other>.
        ---Category: Methods to modify the class definition
        ---C++: alias operator =
        ---C++: return &
 
	----------------------------
	-- Category: Inquire methods
	----------------------------

	Type ( me ) returns TypeOfMarker is static;
	---Level: Public
	---Purpose: Returns the type of the marker style <me> 
	---Category: Inquire methods

        Length ( me ) returns Integer is static;
        ---Level: Public
        ---Purpose: Returns the components length of the marker descriptors
        ---Category: Inquire methods

	Values ( me ; aRank : Integer ;
		      aX,aY : out Real ) returns Boolean
	---Level: Public
	---Purpose: Returns the point and status of a marker style 
	--descriptor of rank <aRank>.
	raises MarkerStyleDefinitionError is static;
	---Trigger:
	-- If aRank is < 1 or > Length()
	---Category: Inquire methods

	XValues ( me ) returns Array1OfShortReal is static;
	---Level: Public
	---Purpose: Returns the X vector of a marker style descriptor
	---Category: Inquire methods
	---C++: return const &

	YValues ( me ) returns Array1OfShortReal is static;
	---Level: Public
	---Purpose: Returns the Y vector of a marker style descriptor
	---Category: Inquire methods
	---C++: return const &

	SValues ( me ) returns Array1OfBoolean is static;
	---Level: Public
	---Purpose: Returns the State vector of a marker style descriptor
	---Category: Inquire methods
	---C++: return const &

    	IsEqual(me; Other : MarkerStyle from Aspect) returns Boolean;
	    ---C++: alias operator==

    	IsNotEqual(me; Other : MarkerStyle from Aspect) returns Boolean;
	    ---C++: alias operator!=

	----------------------------
	-- Category: Private methods
	----------------------------

	SetPredefinedStyle ( me : in out ) is static private;
	---Level: Internal
	---Purpose: Set MyMarkerDescriptor with the predefined style values
	--	    according of current type
	---Category: Private methods

--

fields

--
-- Class	:	Aspect_MarkerStyle
--
-- Purpose	:	Declaration of variables specific to marker styles
--

	MyMarkerType		: TypeOfMarker;
	MyXpoint		: HArray1OfShortReal;
	MyYpoint		: HArray1OfShortReal;
	MySpoint		: HArray1OfBoolean;

end MarkerStyle;
