-- Created by: Peter KURNEV
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SetMapHasher from BOPTools 

	---Purpose: 

uses
    Set from BOPTools

--raises

is
    HashCode(myclass;  
    	    aSet  : Set from BOPTools;  
    	    Upper : Integer from Standard)  
    	returns Integer from Standard;
    ---C++: inline 
     
    IsEqual(myclass;  
    	    aSet1 : Set from BOPTools; 
    	    aSet2 : Set from BOPTools) 
    	returns Boolean from Standard;
    ---C++: inline 

--fields

end SetMapHasher;
