-- File:	IGESGeom_ToolCircularArc.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolCircularArc  from IGESGeom

    ---Purpose : Tool to work on a CircularArc. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses CircularArc from IGESGeom,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolCircularArc;
    ---Purpose : Returns a ToolCircularArc, ready to work


    ReadOwnParams (me; ent : mutable CircularArc;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : CircularArc;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : CircularArc;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a CircularArc <ent>, from
    --           its specific (own) parameters

    DirChecker (me; ent : CircularArc) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : CircularArc;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : CircularArc; entto : mutable CircularArc;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : CircularArc;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolCircularArc;
