-- Created on: 1993-04-26
-- Created by: Jean-Louis Frenkel
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

--   GG  : GER61351 17/11/1999 Change SetColor() with a compatible Quantity_Color instead
--				       the restricted NameOfColor.


class LineAspect from Prs3d inherits BasicAspect from Prs3d
    	---Purpose: A framework for defining how a line will be displayed
    	-- in a presentation. Aspects of line display include
    	-- width, color and type of line.
    	-- The definition set by this class is then passed to the
    	-- attribute manager Prs3d_Drawer.
    	-- Any object which requires a value for line aspect as
    	-- an argument may then be given the attribute manager
    	-- as a substitute argument in the form of a field such as myDrawer for example.
uses 

    AspectLine3d from Graphic3d,
    NameOfColor from Quantity,
    Color from Quantity,
    TypeOfLine from Aspect

is

-- 
--  Attributes for the lines.
-- 
    Create (aColor: NameOfColor from Quantity;
	    aType: TypeOfLine from Aspect;
    	    aWidth: Real from Standard)
	    returns mutable LineAspect from Prs3d;
    	---Purpose: Constructs a framework for line aspect defined by
    	-- -   the color aColor
    	-- -   the type of line aType and
    	-- -   the line thickness aWidth.
    	--   Type of line refers to whether the line is solid or dotted, for example.
        
    Create (aColor: Color from Quantity;
	    aType: TypeOfLine from Aspect;
    	    aWidth: Real from Standard)
	    returns mutable LineAspect from Prs3d;
	    
    SetColor (me: mutable; aColor: Color from Quantity) is static;

    SetColor (me: mutable; aColor: NameOfColor from Quantity) 
    	---Purpose: Sets the line color defined at the time of construction.
    	--          Default value: Quantity_NOC_YELLOW
    is static;
    
    SetTypeOfLine (me: mutable; aType: TypeOfLine from Aspect) 
    	---Purpose: Sets the type of line defined at the time of construction.
    	-- This could, for example, be solid, dotted or made up of dashes.
    	--          Default value: Aspect_TOL_SOLID
    is static;
    
    SetWidth  (me: mutable; aWidth: Real from Standard) 
   	---Purpose: Sets the line width defined at the time of construction.
    	--          Default value: 1.
    is static;

    Aspect(me) returns AspectLine3d from Graphic3d 
    is static;
    	--- Purpose: Returns the line aspect. This is defined as the set of
    	-- color, type and thickness attributes.
            
fields

    myAspect: AspectLine3d from Graphic3d;

end LineAspect from Prs3d;
