-- Created on: 2002-12-12
-- Created by: data exchange team
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class ParametricCurve3dElementCoordinateDirection from StepFEA
inherits FeaRepresentationItem from StepFEA

    ---Purpose: Representation of STEP entity ParametricCurve3dElementCoordinateDirection

uses
    HAsciiString from TCollection,
    Direction from StepGeom

is
    Create returns ParametricCurve3dElementCoordinateDirection from StepFEA;
	---Purpose: Empty constructor

    Init (me: mutable; aRepresentationItem_Name: HAsciiString from TCollection;
                       aOrientation: Direction from StepGeom);
	---Purpose: Initialize all fields (own and inherited)

    Orientation (me) returns Direction from StepGeom;
	---Purpose: Returns field Orientation
    SetOrientation (me: mutable; Orientation: Direction from StepGeom);
	---Purpose: Set field Orientation

fields
    theOrientation: Direction from StepGeom;

end ParametricCurve3dElementCoordinateDirection;
