-- Created on: 1993-03-03
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



private class ItemLocation from PTopLoc inherits Persistent

	---Purpose: Provides  support  for  the implementation  of the
	--          class Location.

uses
    Datum3D  from PTopLoc,
    Location from PTopLoc

is
    Create(D : Datum3D from PTopLoc; 
    	   P : Integer from Standard;
	   N : Location from PTopLoc) 
    returns mutable ItemLocation from  PTopLoc;
	---Level: Internal 
    
    Datum3D(me) returns Datum3D from PTopLoc
    is static;
	---Level: Internal 

    Power(me)   returns Integer from Standard
    is static;
	---Level: Internal 
    
    Next(me)    returns Location from PTopLoc
    is static;
	---Level: Internal 
    
fields
    myDatum : Datum3D  from PTopLoc;
    myPower : Integer  from Standard;
    myNext  : Location from PTopLoc;

end ItemLocation;
