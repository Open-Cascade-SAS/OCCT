-- Created on: 1995-12-07
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class GeometricRepresentationContextAndGlobalUnitAssignedContext from StepGeom 

inherits RepresentationContext from StepRepr


	--- This classe is an implementation of EXPRESS
	--  ANDOR Subtype Declaration.
uses

	GeometricRepresentationContext from StepGeom, 
	GlobalUnitAssignedContext from StepRepr, 
	HAsciiString from TCollection, 
	Integer from Standard, 
	HArray1OfNamedUnit from StepBasic,
	NamedUnit from StepBasic
is

	Create returns GeometricRepresentationContextAndGlobalUnitAssignedContext;
	---Purpose: Returns a GeometricRepresentationContextAndGlobalUnitAssignedContext


	Init (me : mutable;
	      aContextIdentifier : HAsciiString from TCollection;
	      aContextType : HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      aContextIdentifier : HAsciiString from TCollection;
	      aContextType : HAsciiString from TCollection;
	      aGeometricRepresentationContext : GeometricRepresentationContext from StepGeom;
	      aGlobalUnitAssignedContext : GlobalUnitAssignedContext from StepRepr) is virtual;

	Init (me : mutable;
	      aContextIdentifier : HAsciiString from TCollection;
	      aContextType : HAsciiString from TCollection;
	      aCoordinateSpaceDimension : Integer from Standard;
	      aUnits : HArray1OfNamedUnit from StepBasic) is virtual;

	-- Specific Methods for Field Data Access --

	SetGeometricRepresentationContext(me : mutable; aGeometricRepresentationContext : GeometricRepresentationContext);
	GeometricRepresentationContext (me) returns GeometricRepresentationContext;
	SetGlobalUnitAssignedContext(me : mutable; aGlobalUnitAssignedContext : GlobalUnitAssignedContext);
	GlobalUnitAssignedContext (me) returns GlobalUnitAssignedContext;

	-- Specific Methods for ANDOR Field Data Access --

	SetCoordinateSpaceDimension(me : mutable; aCoordinateSpaceDimension : Integer);
	CoordinateSpaceDimension (me) returns Integer;

	-- Specific Methods for ANDOR Field Data Access --

	SetUnits(me : mutable; aUnits : HArray1OfNamedUnit);
	Units (me) returns HArray1OfNamedUnit;
	UnitsValue (me; num : Integer) returns NamedUnit;
	NbUnits (me) returns Integer;

fields

	geometricRepresentationContext : GeometricRepresentationContext from StepGeom;
	globalUnitAssignedContext : GlobalUnitAssignedContext from StepRepr;

end GeometricRepresentationContextAndGlobalUnitAssignedContext;
