-- Created on: 1995-12-21
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SolidBuilder from TopOpeBRepBuild 

uses

    Shape from TopoDS,
    
    ShapeSet from TopOpeBRepBuild,
    LoopSet from TopOpeBRepBuild,
    BlockIterator from TopOpeBRepBuild,
    BlockBuilder from TopOpeBRepBuild,

    ShellFaceSet from TopOpeBRepBuild,
    SolidAreaBuilder from TopOpeBRepBuild
    
is

    Create returns SolidBuilder;

    Create(FS : in out ShellFaceSet; ForceClass : Boolean = Standard_False)  
    returns SolidBuilder;
    ---Purpose: Create a SolidBuilder to build the areas on
    -- the shapes (shells, blocks of faces) described by <LS>.

    InitSolidBuilder(me : in out; 
    	    	     FS : in out ShellFaceSet;
    	    	     ForceClass : Boolean) is static;
    
    -- Output methods 
    InitSolid(me : in out) returns Integer from Standard;
    MoreSolid(me) returns Boolean from Standard is static;
    NextSolid(me : in out) is static;
    
    -- Exploration of the wires of the current Solid
    InitShell(me : in out) returns Integer from Standard;
    MoreShell(me) returns Boolean from Standard is static;
    NextShell(me : in out) is static;
    IsOldShell(me) returns Boolean from Standard is static;
    OldShell(me) returns Shape from TopoDS is static;
    ---Purpose: Returns current shell
    -- This shell may be : 
    -- * an old shell OldShell(), which has not been reconstructed;
    -- * a new shell made of faces described by ...NewFace() methods.
    ---C++: return const &

    -- Exploration of the faces of current shell when IsOldShell = False
    InitFace(me : in out) returns Integer from Standard;
    MoreFace(me) returns Boolean from Standard is static;
    NextFace(me : in out) is static;
    Face(me) returns Shape from TopoDS is static;
    ---Purpose: Returns current new face of current new shell.
    ---C++: return const &

    --- private
    MakeLoops(me : in out; SS : in out ShapeSet from TopOpeBRepBuild) 
    is static private;
    
fields

    myLoopSet : LoopSet from TopOpeBRepBuild;
    myBlockIterator : BlockIterator from TopOpeBRepBuild;
    myBlockBuilder : BlockBuilder from TopOpeBRepBuild;

    mySolidAreaBuilder : SolidAreaBuilder from TopOpeBRepBuild;
    
end SolidBuilder;
