-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class CartesianPoint from StepGeom 

inherits Point from StepGeom 

uses

	HArray1OfReal from TColStd, 
	Real from Standard, 
	HAsciiString from TCollection
is

	Create returns mutable CartesianPoint;
	---Purpose: Returns a CartesianPoint


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aCoordinates : mutable HArray1OfReal from TColStd) is virtual;

    	Init2D (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      X,Y : Real);

    	Init3D (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      X,Y,Z : Real);

	-- Specific Methods for Field Data Access --

	SetCoordinates(me : mutable; aCoordinates : mutable HArray1OfReal);
	Coordinates (me) returns mutable HArray1OfReal;
	CoordinatesValue (me; num : Integer) returns Real;
	NbCoordinates (me) returns Integer;

fields

    nbcoord : Integer; -- optimised formula
    coords  : Real[3];
--	coordinates : HArray1OfReal from TColStd;

end CartesianPoint;
