-- Created on: 1992-09-30
-- Created by: Gilles DEBARBOUILLE
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Bisector from MAT

	---Purpose:

inherits

    TShared from MMgt

uses

    ListOfBisector from MAT,
    Edge from MAT

is

    Create

    ---Purpose:

    returns mutable Bisector from MAT;
    
    AddBisector(me ; abisector : any Bisector from MAT)
    
    is static;
    
    List(me) returns any ListOfBisector from MAT
    
    is static;
    
    FirstBisector(me) returns any Bisector from MAT
    
    is static;

    LastBisector(me) returns any Bisector from MAT
    
    is static;

    BisectorNumber(me : mutable ; anumber : Integer)
    
    is static;
    
    IndexNumber(me : mutable ; anumber : Integer)
    
    is static;
    
    FirstEdge(me : mutable ; anedge : any Edge from MAT)
    
    is static;
    
    SecondEdge(me : mutable ; anedge : any Edge from MAT)
    
    is static;
    
    IssuePoint(me : mutable ; apoint : Integer)
    
    is static;
    
    EndPoint(me : mutable ; apoint : Integer)
    
    is static;

    DistIssuePoint(me : mutable ; areal : Real)
    
    is static;
    
    FirstVector(me : mutable ; avector : Integer)
    
    is static;
    
    SecondVector(me : mutable ; avector : Integer)
    
    is static;
    
    Sense(me : mutable ; asense : Real)
    
    is static;
    
    FirstParameter(me : mutable ; aparameter : Real)
    
    is static;
    
    SecondParameter(me : mutable ; aparameter : Real)
    
    is static;
    
    BisectorNumber(me) returns Integer
    
    is static;
    
    IndexNumber(me) returns Integer
    
    is static;
    
    FirstEdge(me) returns any Edge from MAT
    
    is static;
    
    SecondEdge(me) returns any Edge from MAT
    
    is static;
    
    IssuePoint(me) returns Integer
    
    is static;
    
    EndPoint(me) returns Integer
    
    is static;

    DistIssuePoint(me) returns Real
    
    is static;
			    
    FirstVector(me) returns Integer
    
    is static;
    
    SecondVector(me) returns Integer
    
    is static;
    
    Sense(me) returns Real
    
    is static;
    
    FirstParameter(me) returns Real
    
    is static;
    
    SecondParameter(me) returns Real
    
    is static;
    
    Dump(me ; ashift , alevel : Integer)
    
    is static;
    
fields

    thebisectornumber  : Integer;
    theindexnumber     : Integer;
    thefirstedge       : Edge from MAT;
    thesecondedge      : Edge from MAT;
    thelistofbisectors : ListOfBisector from MAT;
    theissuepoint      : Integer;
    theendpoint        : Integer;
    thefirstvector     : Integer;
    thesecondvector    : Integer;
    thesense           : Real;
    thefirstparameter  : Real;
    thesecondparameter : Real;
    distissuepoint     : Real;
end Bisector;
