-- Created on: 1992-12-02
-- Created by: Christian CAILLET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class SelectRootComps  from IFSelect  inherits SelectExtract

    ---Purpose : A SelectRootComps sorts the Entities which are part of Strong
    --           Componants, local roots of a set of Entities : they can be
    --           Single Componants (containing one Entity) or Cycles
    --           This class gives a more secure result than SelectRoots (which
    --           considers only Single Componants) but is longer to work : it
    --           can be used when there can be or there are cycles in a Model
    --           For each cycle, one Entity is given arbitrarily
    --           Reject works as for SelectRoots : Strong Componants defined in
    --           the input list which are not local roots are given

uses AsciiString from TCollection, InterfaceModel, EntityIterator, Graph

is

    Create returns mutable SelectRootComps;
    ---Purpose : Creates a SelectRootComps

    RootResult (me; G : Graph) returns EntityIterator  is redefined;
    ---Purpose : Returns the list of local root strong componants, by one
    --           Entity par componant. It is redefined for a purpose of
    --           effeciency : calling a Sort routine for each Entity would
    --           cost more ressource than to work in once using a Map
    --           RootResult takes in account the Direct status

    HasUniqueResult (me) returns Boolean  is redefined protected;
    ---Purpose : Returns True, RootResult assuring uniqueness

    Sort (me; rank : Integer; ent : Transient; model : InterfaceModel)
    	returns Boolean;
    ---Purpose : Returns always True, because RootResult has done work

    ExtractLabel (me) returns AsciiString from TCollection;
    ---Purpose : Returns a text defining the criterium : "Local Root Componants"

end SelectRootComps;
