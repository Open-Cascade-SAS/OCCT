-- Created on: 1997-12-01
-- Created by: Jean-Louis Frenkel
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class  ReferenceIterator from PCDM inherits Transient from Standard

uses MetaData from CDM,  
    SequenceOfReference from PCDM,  
    Document from CDM, Application from CDM,
    MessageDriver from  CDM
is
    Create (theMessageDriver : MessageDriver from  CDM)
    returns mutable ReferenceIterator from PCDM;
    ---Purpose:  Warning! The constructor does not initialization.


    LoadReferences(me: mutable; aDocument: Document from CDM; aMetaData: MetaData from CDM; anApplication: Application from CDM; UseStorageConfiguration: Boolean from Standard);
    

    Init(me: mutable;aMetaData: MetaData from CDM)
    is virtual;
  
    More(me) returns Boolean from Standard
    is virtual private;

    Next(me: mutable)
    is virtual private;
    
    MetaData(me;UseStorageConfiguration: Boolean from Standard ) 
    returns MetaData from CDM
    is virtual private;


    ReferenceIdentifier(me)  returns Integer from Standard
    is virtual private;

    DocumentVersion(me) returns Integer from Standard
    ---Purpose: returns the version of the document in the reference
    is virtual private;
    
fields
    myReferences: SequenceOfReference from PCDM;
    myIterator: Integer from Standard; 
    myMessageDriver : MessageDriver from CDM; 
   
end ReferenceIterator from PCDM;
