-- Created by: NW,JPB,CAL
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Vertex from Graphic3d

        ---Purpose: This class allows the creation and update of a
	--	    3D point.

	is

	Create
		returns Vertex from Graphic3d;
	---Level: Public
	---Purpose: Creates a point with 0.0, 0.0, 0.0 coordinates.

	Create ( APoint	: Vertex from Graphic3d )
		returns Vertex from Graphic3d;
	---Level: Public
	---Purpose: Creates a point with coordinates identical to <APoint>.
	--
	-- It's just a copy, but this simplifies the management
	-- of the constructors of VertexC, VertexN and VertexNC.

	Create ( AX, AY ,AZ	: Real from Standard )
		returns Vertex from Graphic3d;
	---Level: Public
	---Purpose: Creates a point with <AX>, <AY> and <AZ> coordinates.

	---------------------------------------------------
	-- Category: Methods to modify the class definition
	---------------------------------------------------

	SetCoord ( me			: in out;
		   Xnew, Ynew, Znew	: Real from Standard )
		is static;
	---Level: Public
	---Purpose: Modifies the coordinates of the point <me>.
	---Category: Methods to modify the class definition

	SetXCoord ( me		: in out;
		    Xnew	: Real from Standard )
		is static;
	---Level: Public
	---Purpose: Modifies the X coordinate of the point <me>.
	---Category: Methods to modify the class definition

	SetYCoord ( me		: in out;
		    Ynew	: Real from Standard )
		is static;
	---Level: Public
	---Purpose: Modifies the Y coordinate of the point <me>.
	---Category: Methods to modify the class definition

	SetZCoord ( me		: in out;
		    Znew	: Real from Standard )
		is static;
	---Level: Public
	---Purpose: Modifies the Z coordinate of the point <me>.
	---Category: Methods to modify the class definition

	----------------------------
	-- Category: Inquire methods
	----------------------------

	Coord ( me;
		AX, AY, AZ	: out Real from Standard )
		is static;
	---Level: Public
	---Purpose: Returns the coordinates of the point <me>.
	---Category: Inquire methods

	X ( me )
		returns Real from Standard
		is static;
	---Level: Public
	---Purpose: Returns the X coordinates of the point <me>.
	---Category: Inquire methods

	Y ( me )
		returns Real from Standard
		is static;
	---Level: Public
	---Purpose: Returns the Y coordinate of the point <me>.
	---Category: Inquire methods

	Z ( me )
		returns Real from Standard
		is static;
	---Level: Public
	---Purpose: Returns the Z coordinate of the point <me>.
	---Category: Inquire methods

	--------------------------
	-- Category: Class methods
	--------------------------

	Distance ( myclass;
		   AV1	: Vertex from Graphic3d;
		   AV2	: Vertex from Graphic3d )
		returns Real from Standard;
	---Level: Public
	---Purpose: Returns the distance between <AV1> and <AV2>.
	---Category: Class methods

--

fields

--
-- Class	:	Graphic3d_Vertex
--
-- Purpose	:	Declaration of variables specific to points
--
-- Reminder	:	A point is defined by its coordinates
--
--

	-- the coordinates of a point
	MyX		:	ShortReal from Standard;
	MyY		:	ShortReal from Standard;
	MyZ		:	ShortReal from Standard;

end Vertex;
