-- Created on: 1993-01-09
-- Created by: CKY / Contract Toubro-Larsen ( TCD )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class DrawingUnits from IGESGraph  inherits IGESEntity

        ---Purpose: defines IGESDrawingUnits, Type <406> Form <17>
        --          in package IGESGraph
        --
        --          Specifies the drawing space units as outlined
        --          in the Drawing entity

uses

        HAsciiString from TCollection

is

        Create returns mutable DrawingUnits;

        -- Specific Methods pertaining to the class

        Init (me      : mutable;
              nbProps : Integer;
              aFlag   : Integer;
              aUnit   : HAsciiString from TCollection);
        ---Purpose : This method is used to set the fields of the class
        --           DrawingUnits
        --      - nbProps : Number of property values (NP = 2)
        --      - aFlag   : DrawingUnits Flag
        --      - aUnit   : DrawingUnits Name

        NbPropertyValues  (me) returns Integer;
        ---Purpose : returns the number of property values in <me>

        Flag (me) returns Integer;
        ---Purpose : returns the drawing space units of <me>

        Unit (me) returns HAsciiString from TCollection;
        ---Purpose : returns the name of the drawing space units of <me>

    	    --  additionnal information, deducted from Flag

    	UnitValue (me) returns Real;
	---Purpose : Computes the value of the unit, in meters, according Flag
	--           (same values as for GlobalSection from IGESData)

fields

--
-- Class    : IGESGraph_DrawingUnits
--
-- Purpose  : Declaration of the variables specific to a Drawing Unit.
--
-- Reminder : A Drawing Unit is defined by :
--                  - Number of property values (NP = 2)
--                  - Units Flag
--                  - Units Name
--

        theNbPropertyValues : Integer;

        theFlag             : Integer;

        theUnit             : HAsciiString from TCollection;

end DrawingUnits;
