-- Created on: 1993-09-01
-- Created by: Laurent PAINNOT
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class Function from AppCont

    ---Purpose: deferred class describing a continous 3d function f(u)


uses Pnt from gp,
     Vec from gp

is

    Delete(me:out) is virtual;
    ---C++: alias "Standard_EXPORT virtual ~AppCont_Function(){Delete() ; }"
    

    FirstParameter(me) returns Real
    	---Purpose: returns the first parameter of the function.
    is deferred;

    LastParameter(me) returns Real
    	---Purpose: returns the last parameter of the function.
    is deferred;

    Value(me; U: Real) returns Pnt
    	---Purpose: returns the point at parameter <U>.
    is deferred;

    D1(me; U: Real; P: in out Pnt; V: in out Vec) returns Boolean
    	---Purpose: returns the point and the derivative values at
    	--          the parameter <U>.
    is deferred;
    
    
end Function;    
