-- Created on: 2012-12-06
-- Created by: Sergey KHROMOV
-- Copyright (c) 2004-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class POnSurfParams from Extrema inherits POnSurf from Extrema
    ---Purpose: Data container for point on surface parameters. These parameters
    --          are required to compute an initial approximation for extrema
    --          computation.
    
uses
    
    POnSurf     from Extrema,
    ElementType from Extrema,
    Pnt         from gp
    
is
    Create returns POnSurfParams;
	    ---Purpose: empty constructor
    	---C++: inline

    Create (theU, theV: Real from Standard; thePnt: Pnt from gp)
    	---Purpose: Creation of a point on surface with parameter 
    	--          values on the surface and a Pnt from gp.
    	---C++: inline
    returns POnSurfParams;

    SetSqrDistance(me: in out; theSqrDistance: Real from Standard);
	    ---Purpose: Sets the square distance from this point to another one
	    --          (e.g. to the point to be projected).
    	---C++: inline

    GetSqrDistance(me)
	    ---Purpose: Query the square distance from this point to another one.
    	---C++: inline
    returns Real from Standard;

    SetElementType(me: in out; theElementType: ElementType from Extrema);
	    ---Purpose: Sets the element type on which this point is situated.
    	---C++: inline

    GetElementType(me)
	    ---Purpose: Query the element type on which this point is situated.
    	---C++: inline
    returns ElementType from Extrema;
    
    SetIndices(me: in out; theIndexU: Integer from Standard;
                           theIndexV: Integer from Standard);
	    ---Purpose: Sets the U and V indices of an element that contains
	    --          this point.
    	---C++: inline

    GetIndices(me; theIndexU: out Integer from Standard;
                   theIndexV: out Integer from Standard);
	    ---Purpose: Query the U and V indices of an element that contains
	    --          this point.
    	---C++: inline

fields

    mySqrDistance : Real        from Standard;
    myElementType : ElementType from Extrema;
    myIndexU      : Integer     from Standard;
    myIndexV      : Integer     from Standard;
    
end POnSurfParams;
