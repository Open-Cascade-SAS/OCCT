-- Created on: 1992-10-14
-- Created by: Gilles DEBARBOUILLE
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Edge from MAT 

	---Purpose: 

inherits

    TShared from MMgt
    
uses

    Bisector from MAT,
    ListOfEdge from MAT

--raises

is

    Create returns mutable Edge from MAT;
    
    EdgeNumber(me : mutable ; anumber : Integer)

    is static;
    
    FirstBisector(me : mutable ; abisector : any Bisector from MAT)

    is static;
    
    SecondBisector(me : mutable ; abisector : any Bisector from MAT)

    is static;
    
    Distance(me : mutable ; adistance : Real)

    is static;
    
    IntersectionPoint(me : mutable ; apoint : Integer)

    is static;

    EdgeNumber(me) returns Integer

    is static;
    
    FirstBisector(me) returns any Bisector from MAT

    is static;
    
    SecondBisector(me) returns any Bisector from MAT

    is static;
    
    Distance(me) returns Real

    is static;
    
    IntersectionPoint(me) returns Integer

    is static;

    Dump(me ; ashift , alevel : Integer)
    
    is static;
    
fields

    theedgenumber        : Integer;
    thefirstbisector     : Bisector from MAT;
    thesecondbisector    : Bisector from MAT;
    thedistance          : Real;
    theintersectionpoint : Integer;

end Edge;
