-- Created on: 1999-11-26
-- Created by: Andrey BETENEV
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0

class CcDesignSecurityClassification from StepAP203
inherits SecurityClassificationAssignment from StepBasic

    ---Purpose: Representation of STEP entity CcDesignSecurityClassification

uses
    SecurityClassification from StepBasic,
    HArray1OfClassifiedItem from StepAP203

is
    Create returns CcDesignSecurityClassification from StepAP203;
	---Purpose: Empty constructor

    Init (me: mutable; aSecurityClassificationAssignment_AssignedSecurityClassification: SecurityClassification from StepBasic;
                       aItems: HArray1OfClassifiedItem from StepAP203);
	---Purpose: Initialize all fields (own and inherited)

    Items (me) returns HArray1OfClassifiedItem from StepAP203;
	---Purpose: Returns field Items
    SetItems (me: mutable; Items: HArray1OfClassifiedItem from StepAP203);
	---Purpose: Set field Items

fields
    theItems: HArray1OfClassifiedItem from StepAP203;

end CcDesignSecurityClassification;
