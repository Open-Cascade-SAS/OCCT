-- File:	Extrema_GenExtPS.cdl
-- Created:	Tue Jul 18 08:20:44 1995
-- Author:	Modelistation
--		<model@metrox>
---Copyright:	 Matra Datavision 1995


class   GenExtPS from Extrema 

    	---Purpose: It calculates all the extremum distances
    	--          between a point and a surface.
    	--          These distances can be minimum or maximum.

uses  	POnSurf       from Extrema,
    	Pnt           from gp,
	HArray2OfPnt  from TColgp,
	FuncExtPS     from Extrema,
	Surface       from Adaptor3d,
	SurfacePtr    from Adaptor3d

raises  NotDone      from StdFail,
    	OutOfRange   from Standard,
	TypeMismatch from Standard
	

is

    Create returns GenExtPS;
    
    Create (P: Pnt; S: Surface from Adaptor3d; NbU,NbV: Integer; TolU,TolV: Real)
    	returns GenExtPS;
      	---Purpose: It calculates all the distances.
        --          The function F(u,v)=distance(P,S(u,v)) has an 
        --          extremum when gradient(F)=0. The algorithm searchs
        --          all the zeros inside the definition ranges of the 
        --          surface.
      	--          NbU and NbV are used to locate the close points
      	--          to find the zeros. They must be great enough
      	--          such that if there is N extrema, there will
      	--          be N extrema between P and the grid.
      	--          TolU et TolV are used to determine the conditions 
      	--          to stop the iterations; at the iteration number n:
      	--           (Un - Un-1) < TolU and (Vn - Vn-1) < TolV .


    Create (P: Pnt; S: Surface from Adaptor3d; NbU,NbV: Integer; 
    	    Umin, Usup, Vmin, Vsup: Real; TolU,TolV: Real)
    	returns GenExtPS;
      	---Purpose: It calculates all the distances.
        --          The function F(u,v)=distance(P,S(u,v)) has an 
        --          extremum when gradient(F)=0. The algorithm searchs
        --          all the zeros inside the definition ranges of the 
        --          surface.
      	--          NbU and NbV are used to locate the close points
      	--          to find the zeros. They must be great enough
      	--          such that if there is N extrema, there will
      	--          be N extrema between P and the grid.
      	--          TolU et TolV are used to determine the conditions 
      	--          to stop the iterations; at the iteration number n:
      	--           (Un - Un-1) < TolU and (Vn - Vn-1) < TolV .

    
    Initialize(me: in out; S: Surface from Adaptor3d; NbU, NbV: Integer; TolU, TolV: Real)
    	---Pupose: sets the fields of the algorithm.
    is static;


    Initialize(me: in out; S: Surface from Adaptor3d; NbU, NbV: Integer; 
    	       Umin, Usup, Vmin, Vsup: Real; TolU, TolV: Real)
    	---Pupose: sets the fields of the algorithm.
    is static;
    

    Perform(me: in out; P: Pnt from gp)
        ---Purpose: the algorithm is done with the point P.
        --          An exception is raised if the fields have not
        --          been initialized.  
    raises TypeMismatch from Standard
    is static;


    IsDone (me) returns Boolean
    	---Purpose: Returns True if the distances are found.
    	is static;
    
    NbExt (me) returns Integer
    	---Purpose: Returns the number of extremum distances.
    	raises  NotDone from StdFail
	    	-- if IsDone(me)=False.
    	is static;

    SquareDistance (me; N: Integer) returns Real
    	---Purpose: Returns the value of the Nth resulting square distance.
    	raises  NotDone from StdFail,
    	    	-- if IsDone(me)=False.
    	        OutOfRange
		-- if N < 1 or N > NbPoints(me).
    	is static;

    Point (me; N: Integer) returns POnSurf
    	---Purpose: Returns the point of the Nth resulting distance.
    	raises  NotDone from StdFail,
    	    	-- if IsDone(me)=False.
    	        OutOfRange
		-- if N < 1 or N > NbPoints(me).
    	is static;

    Bidon(me) returns SurfacePtr from Adaptor3d
    is static private;

fields
    myDone    : Boolean;
    myInit    : Boolean;
    myumin    : Real;
    myusup    : Real;
    myvmin    : Real;
    myvsup    : Real;
    myusample : Integer;
    myvsample : Integer;
    mypoints  : HArray2OfPnt from TColgp;
    mytolu    : Real;
    mytolv    : Real;
    myF	      : FuncExtPS from Extrema;
    myS       : SurfacePtr from Adaptor3d;

end GenExtPS;
