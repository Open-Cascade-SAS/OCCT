-- Created on: 2000-03-01
-- Created by: Denis PASCAL
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Reference from TDF inherits Attribute from TDF

	---Purpose: 

uses Attribute       from TDF,
     Label           from TDF,
     GUID            from Standard,
     DataSet         from TDF,
     RelocationTable from TDF

is


    GetID (myclass)   
    	---C++: return const &  
    returns GUID from Standard;


    Set (myclass; I : Label from TDF; Origin : Label from TDF)
    returns Reference from TDF;
    

    Set (me : mutable; Origin : Label from TDF);
    
    Get (me)
    returns Label from TDF;

    	---Category: TDF_Attribute methods
    	--           =====================
    
    ID (me)
    	---C++: return const & 
    returns GUID from Standard;

    Restore (me: mutable; With : Attribute from TDF);

    NewEmpty (me)
    returns mutable Attribute from TDF;

    Paste (me; Into : mutable Attribute from TDF;
	       RT   : mutable RelocationTable from TDF);    


    References (me; DS : DataSet from TDF) is redefined;

    Dump(me; anOS : in out OStream from Standard)
        returns OStream from Standard
    	is redefined;
	---C++: return &

    Create
    returns mutable Reference from TDF;    


fields

    myOrigin : Label from TDF;

end Reference;
