-- Created on: 1997-08-07
-- Created by: Jean-Louis Frenkel
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package CDF


uses CDM, PCDM, TCollection, TColStd, Resource, Quantity, OSD

is
    class Directory;
    class DirectoryIterator;
    
    class Session;
    
    enumeration TypeOfActivation is TOA_New,TOA_Modified,TOA_Unchanged
    end TypeOfActivation from CDF;
    
    deferred class Application;

    private class StoreList;

---Category: API for Store and retrieve
--           
    
    class Store;

    
    enumeration TryStoreStatus is TS_OK,TS_NoCurrentDocument,TS_NoDriver,TS_NoSubComponentDriver
    end TryStoreStatus;

    enumeration SubComponentStatus is SCS_Consistent, SCS_Unconsistent,SCS_Stored,SCS_Modified
    end SubComponentStatus;
    
    enumeration StoreSetNameStatus  is  
    SSNS_OK, 
    SSNS_ReplacingAnExistentDocument, 
    SSNS_OpenDocument
    end StoreSetNameStatus;
    
    
    ---Category: MetaData management
    --           

    deferred class MetaDataDriver;

    class FWOSDriver;


    exception MetaDataDriverError inherits Failure from Standard;
    ---Purpose: this exception is used in the deferred methods.
    --          Programmer implementing such methods may use this
    --          exception or any exception inheriting MetaDataDriverError.


    deferred class MetaDataDriverFactory;


    private class Timer;
    
    GetLicense(anApplicationIdentifier: Integer from Standard);
    
    IsAvailable(anApplicationIdentifier: Integer from Standard)
    returns Boolean from Standard;

end CDF;
