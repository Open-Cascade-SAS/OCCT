-- Created on: 1992-09-23
-- Created by: Christian CAILLET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class ExternalSources  from IFGraph  inherits GraphContent

    	---Purpose : this class gives entities which are Source of entities of
    	--           a sub-part, but are not contained by this sub-part

uses Transient, EntityIterator, Graph

is

    Create (agraph : Graph) returns ExternalSources;
    ---Purpose : creates empty ExternalSources, ready to work

    GetFromEntity (me : in out; ent : any Transient);
    ---Purpose : adds an entity and its shared ones to the list

    GetFromIter (me : in out; iter : EntityIterator);
    ---Purpose : adds a list of entities (as an iterator) with shared ones

    ResetData (me : in out);
    ---Purpose : Allows to restart on a new data set

    	-- --   Results   -- --
    	--   More-Next-Value give External Source entities

    Evaluate (me : in out) is redefined;
    ---Purpose : Evaluates external sources of a set of entities

    IsEmpty(me : in out) returns Boolean;
    ---Purpose : Returns True if no External Source are found
    --           It means that we have a "root" set
    --           (performs an Evaluation as necessary)

fields

    thegraph : Graph;

end ExternalSources;
