-- Created on: 1995-12-04
-- Created by: Laurent BOURESCHE
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



deferred class TgtField from GeomFill inherits TShared from MMgt

	---Purpose: Root class defining the methods we need to make an
	--          algorithmic tangents field.

uses
    Vec from gp,
    BSpline from Law

is

    IsScalable(me) returns Boolean from Standard is virtual;
    Scale(me : mutable; Func : BSpline from Law) is virtual;

    Value(me; W : Real from Standard)
    returns Vec from gp
    ---Purpose: Computes  the value  of the    field of tangency    at
    --          parameter W.
    is deferred;

    D1(me; W : Real from Standard)
    returns Vec from gp
    ---Purpose: Computes the  derivative of  the field of  tangency at
    --          parameter W.
    is deferred;

    D1(me; W : Real from Standard; V, DV : out Vec from gp)
    ---Purpose: Computes the value and the  derivative of the field of
    --          tangency at parameter W.
    is deferred;

end TgtField;
