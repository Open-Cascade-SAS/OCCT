-- Created on: 1998-01-13
-- Created by: Christian CAILLET
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class SelectBypassSubfigure  from IGESSelect  inherits SelectExplore

    ---Purpose : Selects a list built as follows :
    --           Subfigures correspond to
    --           * Definition (basic : type 308, or Network : type 320)
    --           * Instance (Singular : type 408, or Network : 420, or
    --             patterns : 412,414)
    --           
    --           Entities which are not Subfigure are taken as such
    --           For Subfigures Instances, their definition is taken, then
    --           explored itself
    --           For Subfigures Definitions, the list of "Associated Entities"
    --           is explored
    --           Hence, level 0 (D) recursively explores a Subfigure if some of
    --           its Elements are Subfigures. level 1 explores just at first
    --           level (i.e. for an instance, returns its definition)

uses AsciiString from TCollection, Transient, EntityIterator, Graph

raises InterfaceError

is

    Create (level : Integer = 0) returns mutable SelectBypassSubfigure;
    ---Purpose : Creates a SelectBypassSubfigure, by default all level
    --           (level = 1 explores at first level)

    Explore (me; level : Integer; ent : Transient; G : Graph;
    	     explored : in out EntityIterator)
    	returns Boolean;
    ---Purpose : Explores an entity : for a Subfigure, gives its elements
    --           Else, takes the entity itself


    ExploreLabel (me) returns AsciiString from TCollection;
    ---Purpose : Returns a text defining the criterium : "Content of Subfigure"

end SelectBypassSubfigure;
