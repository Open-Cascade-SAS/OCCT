-- File:        CompositeCurveOnSurface.cdl
-- Created:     Mon Dec  4 12:02:24 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWCompositeCurveOnSurface from RWStepGeom

	---Purpose : Read & Write Module for CompositeCurveOnSurface

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     CompositeCurveOnSurface from StepGeom,
     EntityIterator from Interface

is

	Create returns RWCompositeCurveOnSurface;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable CompositeCurveOnSurface from StepGeom);

	WriteStep (me; SW : in out StepWriter; ent : CompositeCurveOnSurface from StepGeom);

	Share(me; ent : CompositeCurveOnSurface from StepGeom; iter : in out EntityIterator);

end RWCompositeCurveOnSurface;
