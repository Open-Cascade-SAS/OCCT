-- Created on: 1995-01-27
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class IntSS from GeomInt 

	---Purpose: 


uses Intersection    from IntPatch,
     LineConstructor from GeomInt,
     SequenceOfCurve from TColGeom,
     SequenceOfCurve from TColGeom2d,     
     Pnt             from gp,
     Pnt2d           from gp,
     Curve           from Geom,
     Curve           from Geom2d,     
     Surface         from Geom,
     HSurface        from GeomAdaptor,
     TopolTool       from Adaptor3d,
     Line            from IntPatch,
     RLine           from IntPatch,
     Box2d           from Bnd,
     VectorOfReal    from GeomInt
     

raises NotDone    from StdFail,
       OutOfRange from Standard

is

    Create
    	returns IntSS from GeomInt;
	---C++: inline

    Create(S1,S2: Surface from Geom; Tol: Real from Standard; 
           Approx    : Boolean  from  Standard  =  Standard_True;
           ApproxS1  : Boolean  from  Standard  =  Standard_False;
           ApproxS2  : Boolean  from  Standard  =  Standard_False)
    ---Purpose: performs general intersection of two surfaces just now
    	returns IntSS from GeomInt;
	---C++: inline
	
    Perform(me: in out;S1,S2  : Surface from Geom; Tol: Real from Standard;  
    	           Approx     : Boolean  from  Standard  =  Standard_True;
                   ApproxS1   : Boolean  from  Standard  =  Standard_False;
                   ApproxS2   : Boolean  from  Standard  =  Standard_False)
    ---Purpose: general intersection of two surfaces
    	is static;

    Perform(me: in out;HS1,HS2: HSurface from GeomAdaptor; Tol: Real from Standard;  
    	           Approx    : Boolean  from  Standard  =  Standard_True;
                   ApproxS1  : Boolean  from  Standard  =  Standard_False;
                   ApproxS2  : Boolean  from  Standard  =  Standard_False)
    ---Purpose: intersection of adapted surfaces
    	is static;
	---C++: inline

    Perform(me: in out;S1,S2: Surface from Geom; Tol: Real from Standard;  
                   U1,V1,U2,V2: Real from Standard;    	          
    	           Approx    : Boolean  from  Standard  =  Standard_True;
                   ApproxS1  : Boolean  from  Standard  =  Standard_False;
                   ApproxS2  : Boolean  from  Standard  =  Standard_False)
    ---Purpose: general intersection using a starting point
    	is static;

    Perform(me: in out;HS1,HS2: HSurface from GeomAdaptor; Tol: Real from Standard;  
                   U1,V1,U2,V2: Real from Standard;    	          
    	           Approx    : Boolean  from  Standard  =  Standard_True;
                   ApproxS1  : Boolean  from  Standard  =  Standard_False;
                   ApproxS2  : Boolean  from  Standard  =  Standard_False)
    ---Purpose: intersection of adapted surfaces using a starting point
    	is static;
	---C++: inline

    IsDone(me)
    	returns Boolean from Standard
	is static;
	---C++: inline

    TolReached3d(me) returns Real from Standard
    is static;
	---C++: inline

    TolReached2d(me) returns Real from Standard
    is static;
	---C++: inline

    NbLines(me)
    
    	returns Integer from Standard
	---C++: inline
	raises NotDone from StdFail
	is static;
	

    Line(me; Index: Integer from Standard)

    	returns any Curve from Geom
	---C++: return const&
	raises NotDone from StdFail,
	       OutOfRange from Standard

	is static;


    HasLineOnS1(me; Index: Integer from Standard)
    	returns Boolean from Standard;

    LineOnS1(me; Index: Integer from Standard)

    	returns any Curve from Geom2d
	---C++: return const&
	raises NotDone from StdFail,
	       OutOfRange from Standard

	is static;

    HasLineOnS2(me; Index: Integer from Standard)
    	returns Boolean from Standard;

    LineOnS2(me; Index: Integer from Standard)

    	returns any Curve from Geom2d
	---C++: return const&
	raises NotDone from StdFail,
	       OutOfRange from Standard

	is static;


    NbBoundaries(me)
    
    	returns Integer from Standard
	---C++: inline
	raises NotDone from StdFail
	is static;
	

    Boundary(me; Index: Integer from Standard)

    	returns any Curve from Geom
	---C++: return const&
	raises NotDone from StdFail,
	       OutOfRange from Standard

	is static;



    NbPoints(me)
    
    	returns Integer from Standard
	---C++: inline
	raises NotDone from StdFail
	is static;
	

    Point(me; Index: Integer from Standard)

    	returns Pnt from gp
	---C++: inline
	raises NotDone from StdFail,
	       OutOfRange from Standard

	is static;


    Pnt2d(me; Index: Integer from Standard;
              OnFirst: Boolean from Standard)
    
        returns Pnt2d from gp
	raises NotDone from StdFail,
	       OutOfRange from Standard
	is static;

    SetTolFixTangents(me:out;   
    	    aTolCheck:Real from Standard;
    	    aTolAngCheck:Real from Standard); 
	 
    TolFixTangents(me:out;   
    	    aTolCheck:out Real from Standard;
    	    aTolAngCheck:out Real from Standard);     

    TreatRLine(myclass; theRL: RLine from IntPatch;
                theHS1, theHS2: HSurface from GeomAdaptor;
                theC3d: out Curve from Geom;
                theC2d1, theC2d2: out Curve from Geom2d;
                theTolReached: out Real from Standard);
    ---Purpose: converts RLine to Geom(2d)_Curve.
            
    BuildPCurves(myclass; f, l : Real from Standard;
                  Tol: out Real from Standard;
                  S: Surface from Geom;
                  C: Curve from Geom;
                  C2d: out Curve from Geom2d);
    ---Purpose: creates 2D-curve on given surface from given 3D-curve
    
    TrimILineOnSurfBoundaries(myclass; theC2d1, theC2d2: Curve from Geom2d;
                              theBound1, theBound2: Box2d from Bnd;
                              theArrayOfParameters: out VectorOfReal from GeomInt);
    ---Purpose: puts into theArrayOfParameters the parameters of intersection
    --          points of given theC2d1 and theC2d2 curves with the boundaries
    --          of the source surface.

--- Private methods
--  
--   
    InternalPerform(me: in out; Tol: Real from Standard;
    	           Approx,ApproxS1,ApproxS2 : Boolean from Standard;
		   useStart : Boolean from Standard;
                   U1,V1,U2,V2: Real from Standard)
    	is static protected;
     
    MakeCurve(me: in out; Ind     : Integer from Standard;
    	                  D1,D2   : TopolTool from Adaptor3d;
			  Tol     : Real from Standard;
                          Approx  : Boolean from Standard;
                          Approx1 : Boolean from Standard;
                          Approx2 : Boolean from Standard)
    	is protected;

fields

    myIntersector  : Intersection    from IntPatch;
    myLConstruct   : LineConstructor from GeomInt;
    myHS1          : HSurface        from GeomAdaptor;
    myHS2          : HSurface        from GeomAdaptor;
    myNbrestr      : Integer         from Standard;
    sline          : SequenceOfCurve from TColGeom;
    slineS1        : SequenceOfCurve from TColGeom2d;
    slineS2        : SequenceOfCurve from TColGeom2d;
    myTolReached2d : Real            from Standard;
    myTolReached3d : Real            from Standard;     
    --
    myTolCheck     : Real            from Standard;  
    myTolAngCheck  : Real            from Standard;  
    --
end IntSS;
