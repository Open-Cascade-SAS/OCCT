-- Created on: 2001-04-24
-- Created by: Christian CAILLET
-- Copyright (c) 2001-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

--		ckyd@photox.paris1.matra-dtv.fr>

class ToleranceValue  from StepShape    inherits TShared

    ---Purpose : Added for Dimensional Tolerances

uses
    MeasureWithUnit from StepBasic

is

    Create returns mutable ToleranceValue;

    Init (me : mutable; lower_bound, upper_bound : MeasureWithUnit from StepBasic);

    LowerBound (me) returns MeasureWithUnit from StepBasic;
    SetLowerBound (me : mutable; lower_bound : MeasureWithUnit from StepBasic);

    UpperBound (me) returns MeasureWithUnit from StepBasic;
    SetUpperBound (me : mutable; upper_bound : MeasureWithUnit from StepBasic);

fields

    theLowerBound : MeasureWithUnit from StepBasic;
    theUpperBound : MeasureWithUnit from StepBasic;

end ToleranceValue;
