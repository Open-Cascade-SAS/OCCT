-- File:	BinMDataStd_NameDriver.cdl
-- Created:	Tue Nov 19 12:22:02 2002
-- Author:	Edward AGAPOV
--		<eap@strelox.nnov.matra-dtv.fr>
---Copyright:	 Matra Datavision 2002

class NameDriver from BinMDataStd  inherits ADriver from BinMDF

        ---Purpose: TDataStd_Name attribute Driver.

uses
    SRelocationTable from BinObjMgt,
    RRelocationTable from BinObjMgt,
    Persistent       from BinObjMgt,
    MessageDriver    from CDM,
    Attribute        from TDF

is
    Create (theMessageDriver:MessageDriver from CDM)
        returns mutable NameDriver from BinMDataStd;

    NewEmpty (me)  returns mutable Attribute from TDF;

    Paste(me; Source     : Persistent from BinObjMgt;
              Target     : mutable Attribute from TDF;
              RelocTable : out RRelocationTable from BinObjMgt)
        returns Boolean from Standard;
    ---Purpose: persistent -> transient (retrieve)

    Paste(me; Source     : Attribute from TDF;
              Target     : in out Persistent from BinObjMgt;
              RelocTable : out SRelocationTable from BinObjMgt);
    ---Purpose: transient -> persistent (store)

end NameDriver;
