-- Created on: 1994-06-16
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class GeneralModule from RWHeaderSection  inherits GeneralModule from StepData
	---Purpose : Defines General Services for HeaderSection Entities
	--           (Share,Check,Copy; Trace already inherited)
	--           Depends (for case numbers) of Protocol from HeaderSection

uses Transient,
     EntityIterator from Interface,
     ShareTool      from Interface,
     Check          from Interface,
     CopyTool       from Interface

is

	Create returns GeneralModule from RWHeaderSection;
	---Purpose : Creates a GeneralModule

	FillSharedCase (me; CN : Integer; ent : Transient;
	iter : in out EntityIterator);
	---Purpose : Specific filling of the list of Entities shared by an Entity
	--           <ent>, according to a Case Number <CN> (provided by HeaderSection
	--           Protocol).

	CheckCase (me; CN : Integer; ent : Transient; shares : ShareTool; ach : in out Check);
	---Purpose : Specific Checking of an Entity <ent>

	CopyCase (me; CN : Integer; entfrom : Transient; entto : Transient; TC : in out CopyTool);
	---Purpose : Specific Copy ("Deep") from <entfrom> to <entto> (same type)
	--           by using a CopyTool which provides its working Map.
	--           Use method Transferred from CopyTool to work


	NewVoid (me; CN : Integer; ent : out Transient) returns Boolean;

end GeneralModule;
