-- Created on: 1994-08-03
-- Created by: Christophe MARION
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class OutLiner from HLRTopoBRep inherits TShared from MMgt

uses
    Integer        from Standard,
    Shape          from TopoDS,
    Face           from TopoDS,
    Projector      from HLRAlgo,
    Data           from HLRTopoBRep,
    MapOfShapeTool from BRepTopAdaptor
is
    Create
    returns OutLiner from HLRTopoBRep;

    Create (OriSh : Shape from TopoDS)
    returns OutLiner from HLRTopoBRep;

    Create (OriS : Shape from TopoDS;
            OutS : Shape from TopoDS)
    returns OutLiner from HLRTopoBRep;

    OriginalShape(me : mutable; OriS : Shape from TopoDS)
    	---C++: inline
    is static;

    OriginalShape(me : mutable) returns Shape from TopoDS
    	---C++: inline
    	---C++: return &
    is static;

    OutLinedShape(me : mutable; OutS : Shape from TopoDS)
    	---C++: inline
    is static;

    OutLinedShape(me : mutable) returns Shape from TopoDS
    	---C++: inline
    	---C++: return &
    is static;

    DataStructure(me : mutable) returns Data from HLRTopoBRep
    	---C++: inline
    	---C++: return &
    is static;

    Fill(me : mutable;
         P     :        Projector      from HLRAlgo;
	 MST   :in out  MapOfShapeTool from BRepTopAdaptor;
         nbIso :        Integer        from Standard)
    is static;
    
    ProcessFace(me : mutable; F :        Face           from TopoDS;
                              S : in out Shape          from TopoDS;
                              M : in out MapOfShapeTool from BRepTopAdaptor)  
	---Purpose: Builds faces from F and add them to S.
    is static private;

    BuildShape(me : mutable; M : in out MapOfShapeTool from BRepTopAdaptor)
    is static private;
    
fields
    myOriginalShape : Shape from TopoDS;
    myOutLinedShape : Shape from TopoDS;
    myDS            : Data  from HLRTopoBRep;

end OutLiner;
