-- Created on: 1999-09-10
-- Created by: Andrey BETENEV
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Styles from STEPConstruct inherits Tool from STEPConstruct

    ---Purpose: Provides a mechanism for reading and writing shape styles
    --          (such as color) to and from the STEP file
    --          This tool maintains a list of styles, either taking them
    --          from STEP model (reading), or filling it by calls to 
    --          AddStyle or directly (writing).
    --          Some methods deal with general structures of styles and
    --          presentations in STEP, but there are methods which deal
    --          with particular implementation of colors (as described in RP)

uses
    WorkSession      from XSControl,
    InterfaceModel   from Interface,
    HGraph           from Interface,
    FinderProcess    from Transfer,
    TransientProcess from Transfer,
    Shape            from TopoDS,
    SequenceOfTransient from TColStd,
    HSequenceOfTransient from TColStd,
    MapOfShape       from TopTools,
    RepresentationItem from StepRepr,
    RepresentationContext from StepRepr,
    PresentationStyleAssignment from StepVisual,
    StyledItem       from StepVisual,
    Colour           from StepVisual,
    Color            from Quantity,
    IndexedDataMapOfTransientTransient from TColStd,
    MechanicalDesignGeometricPresentationRepresentation from StepVisual,
    ContextDependentShapeRepresentation from StepShape,
    ProductDefinitionShape from StepRepr,
    DataMapOfAsciiStringTransient from STEPConstruct,
    DataMapOfPointTransient from STEPConstruct
is

    Create returns Styles;
    	---Purpose: Creates an empty tool

    Create (WS: WorkSession from XSControl) returns Styles;
    	---Purpose: Creates a tool and initializes it
	
    Init (me: in out; WS: WorkSession from XSControl) returns Boolean;
    	---Purpose: Initializes tool; returns True if succeeded

    --Basic methods: general work with styles	

    NbStyles (me) returns Integer;
    	---Purpose: Returns number of defined styles

    Style (me; i: Integer) returns StyledItem from StepVisual;
    	---Purpose: Returns style with given index

    ClearStyles (me: in out);
    	---Purpose: Clears all defined styles and PSA sequence

    AddStyle (me: in out; style: StyledItem from StepVisual);
    	---Purpose: Adds a style to a sequence

    AddStyle (me: in out; item: RepresentationItem from StepRepr;
    	    	          PSA: PresentationStyleAssignment from StepVisual;
    	    	          Override: StyledItem from StepVisual)
    returns StyledItem from StepVisual;
    	---Purpose: Create a style linking giving PSA to the item, and add it to the
	--          sequence of stored styles. If Override is not Null, then 
	--          the resulting style will be of the subtype OverridingStyledItem.
	
    AddStyle (me: in out; Shape: Shape from TopoDS;
    	    	          PSA: PresentationStyleAssignment from StepVisual;
    	    	          Override: StyledItem from StepVisual)
    returns StyledItem from StepVisual;
    	---Purpose: Create a style linking giving PSA to the Shape, and add it to the
	--          sequence of stored styles. If Override is not Null, then 
	--          the resulting style will be of the subtype OverridingStyledItem.
	--          The Sape is used to find corresponding STEP entity by call to
	--          STEPConstruct::FindEntity(), then previous method is called.

    CreateMDGPR (me: in out; Context: RepresentationContext from StepRepr;
    	    	 MDGPR :in out MechanicalDesignGeometricPresentationRepresentation from StepVisual)
    returns Boolean;
    	---Purpose: Create MDGPR, fill it with all the styles previously defined,
	--          and add it to the model
	
    CreateNAUOSRD (me: in out; Context: RepresentationContext from StepRepr;
    	    	   CDSR : ContextDependentShapeRepresentation from StepShape;
    	    	   initPDS : ProductDefinitionShape from StepRepr)
    returns Boolean;
    	---Purpose: Create MDGPR, fill it with all the styles previously defined,
	--          and add it to the model
	--          IMPORTANT: <initPDS> must be null when use for NAUO colors
	--          <initPDS> initialised only for SHUO case.
	
    FindContext (me; Shape: Shape from TopoDS)
    returns RepresentationContext from StepRepr;
    	---Purpose: Searches the STEP model for the RepresentationContext in which
	--          given shape is defined. This context (if found) can be used
	--          then in call to CreateMDGPR()
	
    LoadStyles (me: in out) returns Boolean;
    	---Purpose: Searches the STEP model for the MDGPR or DM entities
	--          (which bring styles) and fills sequence of styles

    LoadInvisStyles (me; InvSyles : in out HSequenceOfTransient from TColStd)
    returns Boolean;
    	---Purpose: Searches the STEP model for the INISIBILITY enteties
	--          (which bring styles) and fills out sequence of styles

    --Specialized methods: work with colors	

    MakeColorPSA (me; item: RepresentationItem from StepRepr;
    	    	      SurfCol: Colour from StepVisual;
    	    	      CurveCol: Colour from StepVisual;
		      isForNAUO : Boolean from Standard = Standard_False)
    returns PresentationStyleAssignment from StepVisual;
    	---Purpose: Create a PresentationStyleAssignment entity which defines
	--          two colors (for filling surfaces and curves)
	--          if isForNAUO true then returns PresentationStyleByContext
	
    GetColorPSA (me: in out; item: RepresentationItem from StepRepr;
    	    	             Col: Colour from StepVisual)
    returns PresentationStyleAssignment from StepVisual;
    	---Purpose: Returns a PresentationStyleAssignment entity which defines 
	--          surface and curve colors as Col. This PSA is either created
	--          or taken from internal map where all PSAs created by this
	--          method are remembered.
	
    GetColors (me; style: StyledItem from StepVisual;
    	    	   SurfCol : out Colour from StepVisual;
    	    	   BoundCol: out Colour from StepVisual;
    	    	   CurveCol: out Colour from StepVisual;
    	    	   IsComponent: in out Boolean from Standard)
    returns Boolean;
    	---Purpose: Extract color definitions from the style entity
	--          For each type of color supported, result can be either
	--          NULL if it is not defined by that style, or last
	--          definition (if they are 1 or more)

    --Auxiliary methods: conversions between STEP and CASCADE color definitions

     EncodeColor (myclass; Col: Color from Quantity) returns Colour from StepVisual;
    	---Purpose: Create STEP color entity by given Quantity_Color
	--          The analysis is performed for whether the color corresponds to
	--          one of standard colors predefined in STEP. In that case, 
	--          PredefinedColour entity is created instead of RGBColour
    
    EncodeColor (myclass; Col: Color from Quantity;
    	    	    	  DPDCs : in out DataMapOfAsciiStringTransient from STEPConstruct;
    	    	    	  ColRGBs : in out DataMapOfPointTransient from STEPConstruct)
    returns Colour from StepVisual;
    	---Purpose: Create STEP color entity by given Quantity_Color
	--          The analysis is performed for whether the color corresponds to
	--          one of standard colors predefined in STEP. In that case, 
	--          PredefinedColour entity is created instead of RGBColour
    
    DecodeColor (myclass; Colour: Colour from StepVisual;
    	 	          Col : out Color from Quantity) 
    returns Boolean;
    	---Purpose: Decodes STEP color and fills the Quantity_Color. 
	--          Returns True if OK or False if color is not recognized
        
fields

    myMapOfStyles : IndexedDataMapOfTransientTransient from TColStd;
    myStyles      : SequenceOfTransient from TColStd;
    myPSA         : SequenceOfTransient from TColStd;

end Styles;
