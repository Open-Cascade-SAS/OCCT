-- Created on: 2005-10-14
-- Created by: Mikhail KLOKOV
-- Copyright (c) 2005-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class CurveRangeLocalizeData from IntTools
uses
    Box from Bnd,
    CurveRangeSample from IntTools,
    MapOfCurveSample from IntTools,
    ListOfCurveRangeSample from IntTools,
    DataMapOfCurveSampleBox from IntTools

is
    Create(theNbSample: Integer from Standard;
    	   theMinRange: Real from Standard)
    	returns CurveRangeLocalizeData from IntTools;

    GetNbSample(me)
    	returns Integer from Standard;
	---C++: inline

    GetMinRange(me)
    	returns Real from Standard;
	---C++: inline

    AddOutRange(me: in out; theRange: CurveRangeSample from IntTools);
    
    AddBox(me: in out; theRange: CurveRangeSample from IntTools;
    	    	       theBox: Box from Bnd);

    FindBox(me; theRange: CurveRangeSample from IntTools;
    	    	theBox: out Box from Bnd)
    	returns Boolean from Standard;

    IsRangeOut(me; theRange: CurveRangeSample from IntTools)
    	returns Boolean from Standard;

    ListRangeOut(me; theList: out ListOfCurveRangeSample from IntTools);

fields
    myNbSampleC: Integer from Standard;
    myMinRangeC: Real from Standard;
    myMapRangeOut: MapOfCurveSample from IntTools;
    myMapBox      : DataMapOfCurveSampleBox from IntTools;

end CurveRangeLocalizeData from IntTools;
