-- File:        HalfSpaceSolid.cdl
-- Created:     Mon Dec  4 12:02:27 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWHalfSpaceSolid from RWStepShape

	---Purpose : Read & Write Module for HalfSpaceSolid

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     HalfSpaceSolid from StepShape,
     EntityIterator from Interface

is

	Create returns RWHalfSpaceSolid;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable HalfSpaceSolid from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : HalfSpaceSolid from StepShape);

	Share(me; ent : HalfSpaceSolid from StepShape; iter : in out EntityIterator);

end RWHalfSpaceSolid;
