-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Axis1Placement from StepGeom 

inherits Placement from StepGeom 

uses

	Direction from StepGeom, 
	Boolean from Standard, 
	HAsciiString from TCollection, 
	CartesianPoint from StepGeom
is

	Create returns mutable Axis1Placement;
	---Purpose: Returns a Axis1Placement


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aLocation : mutable CartesianPoint from StepGeom) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aLocation : mutable CartesianPoint from StepGeom;
	      hasAaxis : Boolean from Standard;
	      aAxis : mutable Direction from StepGeom) is virtual;

	-- Specific Methods for Field Data Access --

	SetAxis(me : mutable; aAxis : mutable Direction);
	UnSetAxis (me:mutable);
	Axis (me) returns mutable Direction;
	HasAxis (me) returns Boolean;

fields

	axis : Direction from StepGeom;   -- OPTIONAL can be NULL
	hasAxis : Boolean from Standard;

end Axis1Placement;
