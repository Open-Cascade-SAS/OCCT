-- Created on: 1993-10-22
-- Created by: Laurent BOURESCHE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Map from ChFiDS 

	---Purpose: Encapsulation of IndexedDataMapOfShapeListOfShape.

uses

    Shape from TopoDS,
    ShapeEnum from TopAbs,
    ListOfShape from TopTools,
    IndexedDataMapOfShapeListOfShape from TopTools

is
    Create returns Map from ChFiDS;
    ---Purpose:  Create an empty Map

    Fill (me : in out; S : Shape from TopoDS; T1,T2 : ShapeEnum from TopAbs)
    ---Purpose: Fills the map with the subshapes of type T1 as keys
    --          and the list of ancestors  of type T2 as items.
    is static;

    Contains(me; S : Shape from TopoDS) 
    returns Boolean from Standard 
    is static;
    
    FindFromKey(me; S : Shape from TopoDS) 
    returns ListOfShape from TopTools 
    ---C++: alias operator()
    ---C++: return const &
    is static;
    
    FindFromIndex(me; I : Integer from Standard) 
    returns ListOfShape from TopTools
    ---C++: alias operator()
    ---C++: return const &
    is static;

fields

    myMap : IndexedDataMapOfShapeListOfShape from TopTools;

end Map;
