-- Created on: 1993-09-07
-- Created by: GG
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class TypeMap from Aspect inherits TShared from MMgt

	---Version: 0.0

	---Purpose: This class defines a TypeMap object.
	---Keywords:
	---Warning:
	---References:
uses
	LineStyle		from Aspect,
	TypeMapEntry 		from Aspect,
	SequenceOfTypeMapEntry 	from Aspect

raises
	BadAccess 	from Aspect

is
	Create returns mutable TypeMap from Aspect;

        AddEntry (me : mutable; AnEntry : TypeMapEntry from Aspect)
	---Level: Public
        ---Purpose: Adds an entry in the type map <me>.
        --  Warning: Raises BadAccess if TypeMap size is exceeded.
        raises BadAccess from Aspect;

        AddEntry (me : mutable; aStyle : LineStyle from Aspect)
                                        returns Integer from Standard;
        ---Level: Public
        ---Purpose: Search an identical type style entry in the type map <me>
        -- and returns the TypeMapEntry Index if exist.
        -- Or add a new entry and returns the computed TypeMapEntry index used.
 
        Size( me ) returns Integer from Standard is static;
        ---Level: Public
        ---Purpose: Returns the Allocated typemap Size
 
        Index( me ; aTypemapIndex : Integer ) returns Integer from Standard
        ---Level: Public
        ---Purpose: Returns the TypeMapEntry.Index of the TypeMap
        --          at rank <aTypemapIndex> .
        raises BadAccess from Aspect is static;
        ---Trigger: Raises BadAccess if the index less than 1 or
        --          greater than Size.
 
	Dump( me ) ;

	Entry ( me ;
		AnIndex : Integer from Standard )
	returns TypeMapEntry from Aspect
	---Level: Public
	---Purpose: Returns the Type map entry with the index <AnIndex>.
	--  Warning: Raises BadAccess if the index less than 1 or
	--	    greater than Size.
	raises BadAccess from Aspect is static;
	---C++: return const &

fields

	mydata	    : 	SequenceOfTypeMapEntry from Aspect is protected;

end TypeMap ;
