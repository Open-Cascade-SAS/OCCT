-- File:        Polyline.cdl
-- Created:     Fri Dec  1 11:11:25 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class Polyline from StepGeom 

inherits BoundedCurve from StepGeom 

uses

	HArray1OfCartesianPoint from StepGeom, 
	CartesianPoint from StepGeom, 
	HAsciiString from TCollection
is

	Create returns mutable Polyline;
	---Purpose: Returns a Polyline


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aPoints : mutable HArray1OfCartesianPoint from StepGeom) is virtual;

	-- Specific Methods for Field Data Access --

	SetPoints(me : mutable; aPoints : mutable HArray1OfCartesianPoint);
	Points (me) returns mutable HArray1OfCartesianPoint;
	PointsValue (me; num : Integer) returns mutable CartesianPoint;
	NbPoints (me) returns Integer;

fields

	points : HArray1OfCartesianPoint from StepGeom;

end Polyline;
