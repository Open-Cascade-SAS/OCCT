-- Created on: 1999-07-19
-- Created by: Denis PASCAL
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Logbook from TFunction

    ---Purpose: This class contains information which is written and
    --          read during the solving process. Information is divided
    --          in three groups.
    --          
    --          * Touched Labels  (modified by the end user), 
    --          * Impacted Labels (modified during execution of the function),
    --          * Valid Labels    (within the valid label scope).

        
uses Label      from TDF,
     LabelMap   from TDF, 
     Logbook    from TFunction

is
    ---Purpose: next methods are solving declaration
    --          ===================================

    Create returns Logbook from TFunction;

    Clear (me :  in  out);
    ---Purpose: Clears this logbook to its default, empty state.
    IsEmpty (me) 
    returns Boolean from Standard;

    SetTouched (me : in  out; L : Label from TDF);
    ---C++ : inline     
    ---Purpose: Sets the label L as a touched label in this logbook.
    -- In other words, L is understood to have been modified by the end user.

    SetImpacted (me : in  out; L : Label from TDF; 
    	    	    	       WithChildren : Boolean from Standard = Standard_False);
    ---Purpose: Sets the label L as an impacted label in this logbook.
    -- This method is called by execution of the function driver.
     
    SetValid (me : in  out; L : Label from TDF; 
    	    	    	    WithChildren : Boolean from Standard = Standard_False);
    ---Purpose: Sets the label L as a valid label in this logbook.

    ChangeValid (me : in  out)    
    ---C++: return &
    ---C++ : inline        
    returns LabelMap from TDF;

    IsModified (me; L : Label from TDF; 
    	    	    WithChildren : Boolean from Standard = Standard_False) 
    ---Purpose: Returns True if the label L is touched  or impacted. This method
    --          is called by <TFunction_FunctionDriver::MustExecute>. 
    --          If <WithChildren> is set to true, the method checks 
    --          all the sublabels of <L> too.
    returns Boolean from Standard; 


    ---Purpose: next method to consult solving result
    --          =====================================

    GetTouched (me)
    ---C++: return const &
    ---C++: inline     
    ---Purpose: 
    -- Returns the map of touched labels in this logbook.
    -- A touched label is the one modified by the end user.
    returns LabelMap from TDF;    

    GetImpacted (me)
    ---C++: return const &
    ---C++: inline     
    ---Purpose:
    -- Returns the map of impacted labels contained in this logbook.    
    returns LabelMap from TDF;

    GetValid (me)
    ---C++: return const &
    ---C++: inline    
    ---Purpose: Returns the map of valid labels in this logbook.
    returns LabelMap from TDF; 

    Done (me : in out; status : Boolean from Standard);
    ---Purpose: Sets if the execution failed
    ---C++: inline     

    IsDone (me)
    returns Boolean from Standard;
    ---C++: inline 

    Dump(me; stream : in out OStream from Standard) 
    ---C++: return &
    returns OStream from Standard;

fields
     
    myTouched        : LabelMap from TDF;  
    myImpacted       : LabelMap from TDF;
    myValid          : LabelMap from TDF;
    isDone           : Boolean  from Standard;

end Logbook;
