-- Created on: 1993-10-22
-- Created by: Laurent BOURESCHE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Map from ChFiDS 

	---Purpose: Encapsulation of IndexedDataMapOfShapeListOfShape.

uses

    Shape from TopoDS,
    ShapeEnum from TopAbs,
    ListOfShape from TopTools,
    IndexedDataMapOfShapeListOfShape from TopTools

is
    Create returns Map from ChFiDS;
    ---Purpose:  Create an empty Map

    Fill (me : in out; S : Shape from TopoDS; T1,T2 : ShapeEnum from TopAbs)
    ---Purpose: Fills the map with the subshapes of type T1 as keys
    --          and the list of ancestors  of type T2 as items.
    is static;

    Contains(me; S : Shape from TopoDS) 
    returns Boolean from Standard 
    is static;
    
    FindFromKey(me; S : Shape from TopoDS) 
    returns ListOfShape from TopTools 
    ---C++: alias operator()
    ---C++: return const &
    is static;
    
    FindFromIndex(me; I : Integer from Standard) 
    returns ListOfShape from TopTools
    ---C++: alias operator()
    ---C++: return const &
    is static;

fields

    myMap : IndexedDataMapOfShapeListOfShape from TopTools;

end Map;
