-- Created on: 1999-03-10
-- Created by: data exchange team
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class GroupItem from StepAP214 
inherits SelectType from StepData 

uses

    GeometricRepresentationItem from StepGeom


is
    	Create returns GroupItem;
	---Purpose : Returns a GroupItem SelectType
	
    	CaseNum (me; ent : Transient) returns Integer is virtual;
	---Purpose: Recognizes a GroupItem Kind Entity that is :
    	--        1 ->  GeometricRepresentationItem
	--        0 else
	 GeometricRepresentationItem(me) returns any  GeometricRepresentationItem is virtual ;
    	---Purpose : returns Value as a  GeometricRepresentationItem (Null if another type)
	
	
end GroupItem;
