-- Created on: 1992-08-28
-- Created by: Remi LEQUETTE
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package BRepTools 

        ---Level : Public. 
        --  All methods of all  classes will be public.

	---Purpose: The BRepTools package provides  utilities for BRep
	--          data structures.
	--          
	--          * WireExplorer : A tool to explore the topology of
	--          a wire in the order of the edges.
	--          
	--          * ShapeSet :  Tools used for  dumping, writing and
	--          reading.
	--          
	--          * UVBounds : Methods to compute the  limits of the
	--          boundary  of a  face,  a wire or   an edge in  the
	--          parametric space of a face.
	--          
	--          *  Update : Methods  to call when   a topology has
	--          been created to compute all missing data.
	--          
	--          * UpdateFaceUVPoints  :  Method to  update  the UV
	--          points stored   with  the edges   on a face.  This
	--          method ensure that connected  edges  have the same
	--          UV point on their common extremity.
	--          
	--          * Compare : Method to compare two vertices.
	--          
	--          * Compare : Method to compare two edges.
	--          
	--          * OuterWire : A method to find the outer wire of a
	--          face.
	--          
	--          * Map3DEdges : A method to map all the 3D Edges of
	--          a Shape.
	--          
	--          * Dump : A method to dump a BRep object.
	--          

uses
    BRep,
    TopExp,
    TopTools,
    TopoDS,
    TopAbs,
    TopLoc,
    GeomAbs,
    GeomTools,
    Geom,
    Geom2d,
    gp,
    Bnd,
    TColgp,
    TColStd,
    TCollection,
    MMgt,
    Message,
    Poly

is

    class WireExplorer;
    
    deferred class Modification;
    
    class Modifier;

    class TrsfModification;

    class NurbsConvertModification;

    class GTrsfModification;

    class Substitution;

    class Quilt;

    class ShapeSet;

    class ReShape;

    class MapOfVertexPnt2d instantiates DataMap from TCollection
    	(Shape from TopoDS,
    	 SequenceOfPnt2d from TColgp,
	 ShapeMapHasher  from TopTools);
	
    --
    --     Methods
    --     

    UVBounds(F : Face from TopoDS;
             UMin, UMax, VMin, VMax : out Real);
	---Purpose: Returns in UMin,  UMax, VMin,  VMax  the  bounding
	--          values in the parametric space of F.
    
    UVBounds(F : Face from TopoDS;
    	     W : Wire from TopoDS;
             UMin, UMax, VMin, VMax : out Real);
	---Purpose: Returns in UMin,  UMax, VMin,  VMax  the  bounding
	--          values of the wire in the parametric space of F.
    
    UVBounds(F : Face from TopoDS;
    	     E : Edge from TopoDS;
             UMin, UMax, VMin, VMax : out Real);
	---Purpose: Returns in UMin,  UMax, VMin,  VMax  the  bounding
	--          values of the edge in the parametric space of F.
        
    AddUVBounds(F : Face from TopoDS;
                B : in out Box2d from Bnd);
	---Purpose: Adds  to  the box <B>  the bounding values in  the
	--          parametric space of F.
    
    AddUVBounds(F : Face from TopoDS;
    	        W : Wire from TopoDS;
                B : in out Box2d from Bnd);
	---Purpose: Adds  to the box  <B>  the bounding  values of the
	--          wire in the parametric space of F.
    
    AddUVBounds(F : Face from TopoDS;
    	        E : Edge from TopoDS;
    	        B : in out Box2d from Bnd);
	---Purpose: Adds to  the box <B>  the  bounding values  of the
	--          edge in the parametric space of F.


    Update(V : Vertex from TopoDS);
	---Purpose: Update a vertex (nothing is done)

    Update(E : Edge from TopoDS);
	---Purpose: Update an edge, compute 2d bounding boxes.

    Update(W : Wire from TopoDS);
	---Purpose: Update a wire (nothing is done)

    Update(F : Face from TopoDS);
	---Purpose: Update a Face, update UV points.

    Update(S : Shell from TopoDS);
	---Purpose: Update a shell (nothing is done)

    Update(S : Solid from TopoDS);
	---Purpose: Update a solid (nothing is done)

    Update(C : CompSolid from TopoDS);
	---Purpose: Update a composite solid (nothing is done)

    Update(C : Compound from TopoDS);
	---Purpose: Update a compound (nothing is done)

    Update(S : Shape from TopoDS);
	---Purpose: Update a shape, call the corect update.



    UpdateFaceUVPoints(F : Face from TopoDS);
	---Purpose: For  all the edges  of the face  <F> reset  the UV
	--          points to  ensure that  connected  faces  have the
	--          same point at there common extremity.

    Clean(S: Shape from TopoDS);
    	---Purpose: Removes all the triangulations of the faces of <S>
    	--          and removes all polygons on triangulations of the
    	--          edges.

    RemoveUnusedPCurves(S: Shape from TopoDS);
    	---Purpose: Removes all the pcurves of the edges of <S> that
    	--          refer to surfaces not belonging to any face of <S>

    Triangulation(S: Shape from TopoDS; deflec: Real)
    returns Boolean from Standard;
    	---Purpose: verifies that each face from the shape <S> has got
    	--          a triangulation  with a  deflection <= deflec  and
    	--          the edges a discretisation on  this triangulation.


    Compare(V1,V2 : Vertex from TopoDS) returns Boolean;
	---Purpose: Returns  True if  the    distance between the  two
	--          vertices is lower than their tolerance.

    Compare(E1,E2 : Edge from TopoDS) returns Boolean;
	---Purpose: Returns  True if  the    distance between the  two
	--          edges is lower than their tolerance.

    OuterWire(F : Face from TopoDS) returns Wire from TopoDS;
	---Purpose: Returns the outer most wire of <F>. Returns a Null
	--          wire if <F> has no wires.
    
    Map3DEdges(S    : Shape from TopoDS;
    	       M    : in out IndexedMapOfShape from TopTools);
	  ---Purpose: Stores in the map  <M> all the 3D topology edges
	  --          of <S>. 

    IsReallyClosed(E: Edge from TopoDS; F: Face from TopoDS)
	---Purpose: Verifies that the edge  <E> is found two  times on
	--          the face <F> before calling BRep_Tool::IsClosed.
    	returns Boolean from Standard;


    Dump(Sh : Shape from TopoDS; S : in out OStream);
	  ---Purpose: Dumps the topological structure and the geometry 
	  --          of <Sh> on the stream <S>.

    Write(Sh : Shape from TopoDS; S : in out OStream;
          PR : ProgressIndicator from Message = NULL);
	  ---Purpose: Writes <Sh> on <S> in an ASCII format.

    Read(Sh : out Shape from TopoDS; S : in out IStream; 
    	 B  : Builder from  BRep; PR : ProgressIndicator from Message = NULL);
	  ---Purpose: Reads a Shape  from <S> in  returns it in  <Sh>.
	  --          <B> is used to build the shape.

    Write(Sh : Shape from TopoDS; File : CString;
          PR : ProgressIndicator from Message = NULL ) returns Boolean;
	  ---Purpose: Writes <Sh> in <File>.

    Read(Sh : out Shape from TopoDS; File : CString;
    	 B  : Builder from  BRep; PR : ProgressIndicator from Message = NULL)
          returns Boolean;
	  ---Purpose: Reads a Shape  from <File>,  returns it in  <Sh>.
	  --          <B> is used to build the shape.

end BRepTools;


