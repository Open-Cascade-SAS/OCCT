-- Created on: 1993-06-03
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred generic class IWFunction from IntWalk 
    (ThePSurface as any)
 
inherits FunctionSetWithDerivatives from math			 


	---Purpose: Template class for a function on a parametric surface.
	--          the form of the function is F(u,v) = 0 where u and v are
	--          the parameteric coordinates of a point on the surface.

uses Vector  from math,
     Matrix  from math,
     Pnt     from gp,
     Vec     from gp,
     Dir2d   from gp
       

raises UndefinedDerivative from StdFail

is

    Set(me: in out; PS: ThePSurface)
    
    	is static;


    NbVariables(me)

	---Purpose: This method has to return 2.
    	returns Integer from Standard;


    NbEquations(me)

	---Purpose: This method has to return 1.
    	returns Integer from Standard;


    Value(me : in out; X : Vector from math;
                       F : out Vector from math)

	---Purpose: The dimension of F is 1.

    	returns Boolean from Standard;


    Derivatives(me : in out; X : Vector from math;
                             D : out Matrix from math)

	---Purpose: The dimension of D is (1,2).

    	returns Boolean from Standard;


    Values(me : in out; X : Vector from math;
                        F : out Vector from math;
                        D : out Matrix from math)

    	returns Boolean from Standard;


    Root(me)

	---Purpose: Root is the value of the function at the solution.
	--          It is a vector of dimension 1, i-e a real.

    	returns Real from Standard
    	is static;


    Tolerance(me)
    
	---Purpose: Returns the value Tol so that if Abs(Func.Root())<Tol
	--          the function is considered null.
    
    	returns Real from Standard
	is static;


    Point(me)

	---Purpose: Returns the value of the solution point on the surface.

    	returns Pnt from gp
    	is static;
    

    IsTangent(me : in out)

    	returns Boolean from Standard 
    	is static;
    

    Direction3d(me: in out)

    	returns Vec from gp
    	raises UndefinedDerivative from StdFail
    	is static;
    

    Direction2d(me: in out)

    	returns Dir2d from gp
    	raises UndefinedDerivative from StdFail
    	is static;
    

end IWFunction;
