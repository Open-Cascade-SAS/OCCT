-- Created on: 1995-12-19
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Loop from TopOpeBRepBuild inherits TShared from MMgt

---Purpose: 
-- a Loop is an existing shape (Shell,Wire) or a set
-- of shapes (Faces,Edges) which are connex.
-- a set of connex shape is represented by a BlockIterator

uses

    Shape from TopoDS,
    BlockIterator from TopOpeBRepBuild,
    ShapeEnum from TopAbs

is

    Create(S : Shape from TopoDS) returns mutable Loop;
    Create(BI : BlockIterator) returns mutable Loop;
	
    IsShape(me) returns Boolean from Standard is virtual;

    Shape(me) returns Shape from TopoDS is virtual;
    ---C++: return const &
    -- only when IsShape() is true
    
    BlockIterator(me) returns BlockIterator is static;
    ---C++: return const &
    -- only when IsShape() is false

    Dump(me) is virtual;	

fields

    myIsShape       : Boolean from Standard is protected;
    myShape         : Shape from TopoDS     is protected;
    myBlockIterator : BlockIterator         is protected;

end Loop from TopOpeBRepBuild;
