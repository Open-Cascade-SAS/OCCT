-- Created on: 1995-06-12
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ShapeListOfShape from TopOpeBRepBuild

---Purpose: represent shape + a list of shape

uses
    
    ListOfShape from TopTools,
    Shape from TopoDS
    
is

    Create returns ShapeListOfShape from TopOpeBRepBuild;

    Create(S : Shape from TopoDS)
    returns ShapeListOfShape from TopOpeBRepBuild;

    Create(S : Shape from TopoDS;
     	   L : ListOfShape from TopTools)
    returns ShapeListOfShape from TopOpeBRepBuild;

    List(me)
    returns ListOfShape from TopTools is static;
    ---C++: return const &

    ChangeList(me : in out)
    returns ListOfShape from TopTools is static;
    ---C++: return &

    Shape(me) 
    returns Shape from TopoDS is static;
    ---C++: return const &

    ChangeShape(me : in out) 
    returns Shape from TopoDS is static;
    ---C++: return &

fields

    myList : ListOfShape from TopTools;
    myShape : Shape from TopoDS;

end ShapeListOfShape from TopOpeBRepBuild;
