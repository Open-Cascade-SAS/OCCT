-- File:	RWStepAP214_RWAppliedDocumentReference.cdl
-- Created:	Fri Mar 12 12:16:39 1999
-- Author:	data exchange team
--		<det@androx.nnov.matra-dtv.fr>
---Copyright:	 Matra Datavision 1999


class RWAppliedDocumentReference from RWStepAP214 

	---Purpose: Read & Write Module for AppliedDocumentReference

uses
     Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     AppliedDocumentReference from StepAP214,
     EntityIterator from Interface

is

    	Create returns RWAppliedDocumentReference;
    
    	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable AppliedDocumentReference from StepAP214);

	WriteStep (me; SW : in out StepWriter; ent : AppliedDocumentReference from StepAP214);

	Share(me; ent : AppliedDocumentReference from StepAP214; iter : in out EntityIterator);

end RWAppliedDocumentReference;
