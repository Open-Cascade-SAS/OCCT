-- Created on: 1992-10-21
-- Created by: Christian CAILLET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class SingleParentEntity  from IGESData  inherits IGESEntity

    ---Purpose : a SingleParentEntity is a kind of IGESEntity which can refer
    --           to a (Single) Parent, from Associativities list of an Entity
    --           a effective SingleParent definition entity must inherit it

uses Integer

raises OutOfRange

is

    SingleParent (me) returns IGESEntity  is deferred;
    ---Purpose : Returns the parent designated by the Entity, if only one !

    NbChildren (me) returns Integer  is deferred;
    ---Purpose : Returns the count of Entities designated as children

    Child (me; num : Integer) returns IGESEntity
    ---Purpose : Returns a Child given its rank
    	raises OutOfRange  is deferred;
    --           Error if <num> is below one or over <NbChildren>

end SingleParentEntity;
