-- Created on: 2003-08-21
-- Created by: Sergey KUUL
-- Copyright (c) 2003-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class ReprItemAndLengthMeasureWithUnit from StepRepr inherits RepresentationItem from StepRepr

uses
    LengthMeasureWithUnit from StepBasic,
    MeasureRepresentationItem from StepRepr,
    MeasureWithUnit from StepBasic

is

    Create returns mutable ReprItemAndLengthMeasureWithUnit;
    
    Init(me: mutable; aMWU: mutable MeasureWithUnit; aRI : RepresentationItem);

    SetLengthMeasureWithUnit(me: mutable; aLMWU: mutable LengthMeasureWithUnit);
    
    GetLengthMeasureWithUnit(me) returns mutable LengthMeasureWithUnit;

    GetMeasureRepresentationItem(me) returns mutable MeasureRepresentationItem;

    SetMeasureWithUnit(me: mutable; aMWU: mutable MeasureWithUnit);
    
    GetMeasureWithUnit(me) returns mutable MeasureWithUnit;

    GetRepresentationItem(me) returns mutable RepresentationItem;

fields

    myLengthMeasureWithUnit: LengthMeasureWithUnit from StepBasic;
    myMeasureRepresentationItem : MeasureRepresentationItem from StepRepr;
    myMeasureWithUnit: MeasureWithUnit from StepBasic;

end ReprItemAndLengthMeasureWithUnit;
