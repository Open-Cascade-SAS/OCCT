-- Created on: 2008-03-27
-- Created by: Sergey ZARITCHNY
-- Copyright (c) 2008-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class IntPackedMap_1 from PDataStd inherits Attribute from PDF

	---Purpose: Persistence

uses
    HArray1OfInteger  from  PColStd


is
    Create returns mutable  IntPackedMap_1 from  PDataStd;

    Init (me : mutable; theLow,  theUp:  Integer  from Standard);
    ---Purpose: Inits the internal container
    --  if  (upper  -  lower)  ==  0  and (upper  |  lower) == 0, the corresponding  
    --  array is empty (not requested)
     
    IsEmpty (me)
    ---Purpose: Returns true if the internal container is empty
    returns Boolean from Standard;  

    Upper  (me)
     ---Purpose: Returns an upper bound of the internal container
    returns Integer from Standard;   

    Lower  (me)
     ---Purpose: Returns a lower bound of the internal container
    returns Integer from Standard;   
    
    GetValue (me; theIndex : Integer from Standard)  
    returns Integer from Standard;
        
    SetValue (me : mutable; theIndex : Integer from Standard;  
    	    	    	    theValue : Integer from Standard);
     
    SetDelta(me : mutable; delta : Boolean from Standard); 
     
    GetDelta(me) returns Boolean from Standard;
    
fields 

    myIntValues      :  HArray1OfInteger from PColStd;       
    myDelta  : Boolean from Standard;

end IntPackedMap_1;


