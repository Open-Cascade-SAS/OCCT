-- File:	IGESDimen_ToolGeneralNote.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolGeneralNote  from IGESDimen

    ---Purpose : Tool to work on a GeneralNote. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses GeneralNote from IGESDimen,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolGeneralNote;
    ---Purpose : Returns a ToolGeneralNote, ready to work


    ReadOwnParams (me; ent : mutable GeneralNote;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : GeneralNote;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : GeneralNote;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a GeneralNote <ent>, from
    --           its specific (own) parameters

    DirChecker (me; ent : GeneralNote) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : GeneralNote;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : GeneralNote; entto : mutable GeneralNote;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : GeneralNote;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolGeneralNote;
