-- Created on: 2001-04-13
-- Created by: Peter KURNEV
-- Copyright (c) 2001-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class SFSCorrector from BOP 

	---Purpose: 
    	---  the algorithm is to change the Shell Faces Set (SFS)contents.      
    	---  The NewSFS will contain only shells   
    	---  instead of shells and faces.  
        --- 
	 
uses
 
    ShellFaceSet         from BOP,
    PShellFaceSet        from BOP,
    ListOfConnexityBlock from BOP 
    
is 
    Create   
    	returns SFSCorrector from BOP; 
    	---Purpose:  
    	--- Empty constructor; 
    	---
    SetSFS  (me:out; 
		aSFS: ShellFaceSet from BOP);  
    	---Purpose: 
    	--- Modifier 
    	---
    Do (me:out); 
    	---Purpose:
    	--- Performs the algorithm of  two  steps 
    	--- 1. Make conexity blocks (  DoConnexityBlocks()  )     
    	--- 2. Make corrections     (  DoCorrections()  )        
    	---
    DoConnexityBlocks(me:out) 
    	is  private; 
    	---Purpose: 
    	--- Internal Purpose  
    	---
    DoCorrections(me:out) 
    	is  private; 
    	---Purpose: 
    	--- Internal Purpose  
    	---
    IsDone(me)  
    	returns Boolean from Standard;   
    	---Purpose: 
    	--- Selector 
    	---
    ErrorStatus	(me)  
    	returns Integer from Standard; 
    	---Purpose: 
    	--- Selector  
    	--- - 1 - Nothing is done because only constructor has been called
    	---
    SFS     (me:out) 
    	returns ShellFaceSet from BOP; 
    	---C++:  return &  
    	---Purpose: 
    	--- Selector 
    	---
    NewSFS  (me:out) 
    	returns ShellFaceSet from BOP; 
    	---C++:  return &   
    	---Purpose: 
    	--- Selector 
    	--- Returns the resulting SFS
	---

fields 

    mySFS             : PShellFaceSet        from BOP; 
    myNewSFS          : ShellFaceSet         from BOP;  
    myConnexityBlocks : ListOfConnexityBlock from BOP;  
    myIsDone          : Boolean from Standard;  
    myErrorStatus     : Integer from Standard;  

end SFSCorrector;
