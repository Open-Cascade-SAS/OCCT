-- Created on: 1994-02-03
-- Created by: Gilles DEBARBOUILLE
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

generic class EnumerationParameter from Dynamic (Enum as any)

inherits

    Parameter from Dynamic     
    
    ---Purpose: This  generic class defines  a  parameter with a given
    --          enumeration.  For correct use an instanciation of this
    --          class,  the  Convert  method  must  be  defined.  This
    --          method is automaticaly called by the constructor which
    --          takes a  CString  as value for  the  enumeration.  The
    --          prototype  of the Convert method  must be described as
    --          follows :
    --          
    --          void Convert(const Standard_CString,Enum);
    --          
    --          The  prototype  and the body of  this   method, can be
    --          written  in   the  file   <mypackage.cxx>   where  the
    --          enumeration  is described.    No declaration  of   the
    --          Convert method in any .cdl file is necessary.


uses
    CString from Standard,
    OStream from Standard 

is

    Create(aparameter : CString from Standard)
    
    ---Level: Public 
    
    ---Purpose: Creates an  EnumerationParameter  of  <aparameter>  as
    --          name.

    returns mutable EnumerationParameter from Dynamic;

    Create(aparameter : CString from Standard; avalue : Enum)
    
    ---Level: Public 
    
    ---Purpose: Creates  an  EnumerationParameter  of  <aparameter> as
    --          name and <avalue> as value.

    returns mutable EnumerationParameter from Dynamic;
    
    Create(aparameter , avalue : CString from Standard) 

    ---Level: Public 
    
    ---Purpose: Creates an  EnumerationParameter  of  <aparameter>  as
    --          name  and <avalue> as value. The user has to define  a
    --          Convert method to translate  the string <avalue> in an
    --          enumeration term.

    returns mutable EnumerationParameter from Dynamic;
    
    Value(me) returns Enum
    
    ---Level: Public 
    
    ---Purpose: Returns the enumeration value <thevalue>.
    
    is static;
    
    Value (me : mutable ; avalue : Enum)
    
    ---Level: Public 
    
    ---Purpose: Sets the field <thevalue> with the enumeration value <avalue>

    is static;
    
    Dump(me ; astream : in out OStream from Standard)
    
    ---Level: Internal 
    
    ---Purpose: useful for debugging.
    
    is redefined;
    
fields

    thevalue : Enum;

end EnumerationParameter;
