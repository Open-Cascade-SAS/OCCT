-- Created on: 2002-04-01
-- Created by: Peter KURNEV
-- Copyright (c) 2002-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class CoupleOfInteger from BOPTools 

	---Purpose:  
	--  Auxiliary class providing structure to  
	--  store info about a couple of integers 
	 
--uses
--raises

is
    Create 
    	returns CoupleOfInteger from BOPTools; 
    	---Purpose: 
    	--- Empty Constructor
    	---
    Create(aFirst  : Integer from Standard; 
    	   aSecond : Integer from Standard) 
    	returns CoupleOfInteger from BOPTools; 
    	---Purpose: 
    	--- Constructor
    	---
    SetCouple(me:out; 
	   aFirst  : Integer from Standard; 
    	   aSecond : Integer from Standard); 
    	---Purpose: 
    	--- Modifier
    	---
    SetFirst(me:out; 
	   aFirst  : Integer from Standard); 
    	---Purpose: 
    	--- Modifier
    	---
    SetSecond(me:out; 
	   aSecond : Integer from Standard); 
    	---Purpose: 
    	--- Modifier
    	---
    Couple   (me; 
    	   aFirst  :out Integer from Standard; 
    	   aSecond :out Integer from Standard); 	   
    	---Purpose: 
    	--- Selector
    	---
    First(me) 
    	returns Integer from Standard;
    	---Purpose: 
    	--- Selector
    	---
    Second(me) 
    	returns Integer from Standard; 
    	---Purpose: 
    	--- Selector
    	---
  
    IsEqual(me; 
    	    aOther:like me) 
	returns Boolean from Standard;     

    HashCode(me; 
	    Upper : Integer  from Standard)  
    	returns Integer from Standard;  
	
fields 
    myFirst  : Integer from Standard; 
    mySecond : Integer from Standard;   

end CoupleOfInteger;
