-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class RepresentationMap from StepRepr 

inherits TShared from MMgt

uses

	RepresentationItem from StepRepr, 
	Representation from StepRepr
is

	Create returns RepresentationMap;
	---Purpose: Returns a RepresentationMap

	Init (me : mutable;
	      aMappingOrigin : RepresentationItem from StepRepr;
	      aMappedRepresentation : Representation from StepRepr) is virtual;

	-- Specific Methods for Field Data Access --

	SetMappingOrigin(me : mutable; aMappingOrigin : RepresentationItem);
	MappingOrigin (me) returns RepresentationItem;
	SetMappedRepresentation(me : mutable; aMappedRepresentation : Representation);
	MappedRepresentation (me) returns Representation;

fields

	mappingOrigin : RepresentationItem from StepRepr;
	mappedRepresentation : Representation from StepRepr;

end RepresentationMap;
