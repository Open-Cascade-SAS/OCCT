-- Created on: 1991-10-09
-- Created by: Michel CHAUVAT
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



generic class   ExtPSOfRev from Extrema (SurfaceOfRevolution as any;
    	    	    	    	    	 Tool                as any ; -- as ToolSurfaceOfRevolution(SurfaceOfRevolution)
					 Curve               as any;
					 ToolCurve           as any; -- as ToolCurve(Curve)
					 TheExtPC            as any
					)
    	---Purpose: It calculates all the extremum distances
    	--          between a point and a surface.
    	--          These distances can be minimum or maximum.

uses   	POnSurf           from Extrema,
    	SequenceOfPOnSurf from Extrema,
    	Pnt               from gp,
    	SequenceOfReal    from TColStd
	
raises  NotDone    from StdFail,
    	OutOfRange from Standard

is
    Create (P: Pnt; S: SurfaceOfRevolution; Tol: Real; NbV: Integer;
    	    TolV: Real) returns ExtPSOfRev;
      	---Purpose: It calculates all the distances between a point 
      	--          and a surface of revolution.
      	--          Tol is used to test if the point is on the axis.
      	--          NbV and TolV are used to compute the extrema on a 
      	--          meridian (see ExtPC.cdl).

    IsDone (me) returns Boolean
    	---Purpose: Returns True if the distances are found.
    	is static;
    
    NbExt (me) returns Integer
    	---Purpose: Returns the number of extremum distances.
    	raises  NotDone from StdFail
	    	-- if IsDone(me)=False.
    	is static;

    SquareDistance (me; N: Integer) returns Real
    	---Purpose: Returns the value of the Nth resulting square distance.
    	raises  NotDone from StdFail,
    	    	-- if IsDone(me)=False.
    	        OutOfRange
		-- if N < 1 or N > NbPoints(me).
    	is static;

    Point (me; N: Integer) returns POnSurf
    	---Purpose: Returns the point of the Nth resulting distance.
    	raises  NotDone from StdFail,
    	    	-- if IsDone(me)=False.
    	        OutOfRange
		-- if N < 1 or N > NbPoints(me).
    	is static;

fields
    myDone : Boolean;
    mySqDist: SequenceOfReal from TColStd;
    myPoint: SequenceOfPOnSurf from Extrema;

end ExtPSOfRev;
