-- Created on: 1994-03-03
-- Created by: Jean Louis FRENKEL
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



package TColQuantity 

---Purpose: the  classes of this package should be used
--          when exporting arrays of real representing lengths, 
--          for having benefit of the unit conversion.
uses

    TCollection,
    Quantity
    
is
    class Array1OfLength instantiates Array1 from TCollection (Length from Quantity);
    class Array2OfLength instantiates Array2 from TCollection (Length from Quantity);
    class HArray1OfLength        instantiates 
    	HArray1 from TCollection  (Length from Quantity, Array1OfLength from TColQuantity); 
    class HArray2OfLength        instantiates 
    	HArray2 from TCollection  (Length from Quantity, Array2OfLength from TColQuantity); 
end TColQuantity;
