-- Created on: 1997-04-24
-- Created by: Yves FRICAUD
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SameShapeIterator from TNaming 

	---Purpose:  To iterate on   all  the label which contained  a
	--          given shape.

uses
    Shape       from TopoDS,
    UsedShapes  from TNaming,
    Iterator    from TNaming,
    Label       from TDF,
    PtrNode     from TNaming 	

raises
     NoMoreObject from Standard,
     NoSuchObject from Standard 

is

    Create(aShape      : Shape     from TopoDS; 
    	   Shapes      : UsedShapes from TNaming)
    returns SameShapeIterator from TNaming 
    is private;    

    Create(aShape      : Shape     from TopoDS; 
    	   access      : Label from TDF)
    returns SameShapeIterator from TNaming;
    
    More(me) returns Boolean;
    	---C++: inline
    
    Next(me : in out)
    raises
       NoMoreObject from Standard;
       
    Label(me) returns Label from TDF
    raises
	NoSuchObject from Standard;
	
fields
    myNode  : PtrNode from TNaming;	
    myIsNew   : Boolean from Standard;

friends

    class Tool from TNaming
    
end SameShapeIterator;
