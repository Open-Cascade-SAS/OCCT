-- Created on: 2002-12-12
-- Created by: data exchange team
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package RWStepFEA

uses

	StepData, Interface, TCollection, TColStd, StepFEA

is

    class RWAlignedCurve3dElementCoordinateSystem;
    class RWArbitraryVolume3dElementCoordinateSystem;
    class RWCurve3dElementProperty;
    class RWCurve3dElementRepresentation;
    class RWCurveElementEndOffset;
    class RWCurveElementEndRelease;
    class RWCurveElementInterval;
    class RWCurveElementIntervalConstant;
    class RWCurveElementLocation;
    class RWDummyNode;
    class RWElementGeometricRelationship;
    class RWElementGroup;
    class RWElementRepresentation;
    class RWFeaAreaDensity;
    class RWFeaAxis2Placement3d;
    class RWFeaGroup;
    class RWFeaLinearElasticity;
    class RWFeaMassDensity;
    class RWFeaMaterialPropertyRepresentation;
    class RWFeaMaterialPropertyRepresentationItem;
    class RWFeaModel;
    class RWFeaModel3d;
    class RWFeaMoistureAbsorption;
    class RWFeaParametricPoint;
    class RWFeaRepresentationItem;
    class RWFeaSecantCoefficientOfLinearThermalExpansion;
    class RWFeaShellBendingStiffness;
    class RWFeaShellMembraneBendingCouplingStiffness;
    class RWFeaShellMembraneStiffness;
    class RWFeaShellShearStiffness;
    class RWFeaTangentialCoefficientOfLinearThermalExpansion;
    class RWGeometricNode;
    class RWNode;
    class RWNodeGroup;
    class RWNodeRepresentation;
    class RWNodeSet;
    class RWNodeWithSolutionCoordinateSystem;
    class RWNodeWithVector;
    class RWParametricCurve3dElementCoordinateDirection;
    class RWParametricCurve3dElementCoordinateSystem;
    class RWParametricSurface3dElementCoordinateSystem;
    class RWSurface3dElementRepresentation;
    class RWVolume3dElementRepresentation;
    class RWFeaModelDefinition;
    class RWFreedomAndCoefficient;
    class RWFreedomsList;
    class RWNodeDefinition;
    class RWAlignedSurface3dElementCoordinateSystem;
    class RWConstantSurface3dElementCoordinateSystem;
    class RWCurveElementIntervalLinearlyVarying;    -- added 23.01.2003
    class RWFeaCurveSectionGeometricRelationship;   -- added 23.01.2003
    class RWFeaSurfaceSectionGeometricRelationship; -- added 23.01.2003

end;
