-- Created on: 1997-02-06
-- Created by: Denis PASCAL
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Real from TDataStd inherits Attribute  from TDF

    ---Purpose: The basis to define a real number attribute.

uses Attribute       from TDF,
     Label           from TDF,
     GUID            from Standard,
     Real            from Standard,
     RelocationTable from TDF,
     RealEnum        from TDataStd

is

    ---Purpose: class methods
    --          =============

    GetID (myclass)    
    	---C++: return const & 
    	---Purpose:  Returns the GUID for real numbers.   
    returns GUID from Standard;

    Set (myclass ; label : Label from TDF; value : Real from Standard)
    ---Purpose: Finds, or creates, an Real attribute and sets <value> the
    --          Real attribute  is  returned. the  Real  dimension is
    --          Scalar by default. use SetDimension to overwrite.
    returns Real from TDataStd;
    
    ---Purpose: Real methods
    --          ============

    Create
    returns mutable Real from TDataStd; 
    
    SetDimension (me : mutable; DIM : RealEnum from TDataStd);

    
    GetDimension (me)
    returns RealEnum from TDataStd;

    
    Set (me : mutable; V : Real from Standard);
    	---Purpose:
    	-- Finds or creates the real number V.  

    Get (me)
    returns Real from Standard;
    	---Purpose:
    	-- Returns the real number value contained in the attribute.
    IsCaptured(me) returns Boolean;
	---Purpose: Returns True if there is a reference on the same label
    
    ---Category: TDF_Attribute methods
    --           =====================
    
    ID (me) 
    ---C++: return const &  
    returns GUID from Standard;

    Restore (me: mutable; With : Attribute from TDF);

    NewEmpty(me)
    returns mutable Attribute from TDF;

    Paste (me; Into : mutable Attribute from TDF;
	       RT   : mutable RelocationTable from TDF);    

    
    Dump(me; anOS : in out OStream from Standard)
    returns OStream from Standard
    is redefined;
    ---C++: return &

fields

    myValue     : Real     from Standard;
    myDimension : RealEnum from TDataStd;

end Real;
