-- Created on: 1992-04-29
-- Created by: Remi LEQUETTE
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Axis3D from Draw inherits Drawable3D from Draw

	---Purpose: 

uses Pnt from gp,
    Ax3 from gp,
    Color from Draw,
    Display from Draw

is

    Create(col : Color; Size : Integer = 5)
    returns Axis3D;

    Create(p : Pnt; col : Color; Size : Integer = 5)
    returns Axis3D;
    
    Create(A : Ax3 from gp; col : Color; Size : Integer = 5)
    returns Axis3D;
    
    DrawOn(me; dis : in out Display);

fields

    myAxes : Ax3 from gp;
    myColor : Color;
    mySize : Integer;
    
end Axis3D;
