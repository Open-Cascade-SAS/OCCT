-- Created on: 1999-03-25
-- Created by: data exchange team
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SelectAssembly from STEPSelections inherits SelectExplore from IFSelect

	---Purpose: 

uses
    AsciiString from TCollection,
    Transient,
    EntityIterator,
    Graph
is
    Create returns mutable SelectAssembly from STEPSelections;
    
    Explore (me; level : Integer; ent : Transient; G : Graph;
    	     explored : in out EntityIterator)
    returns Boolean;
    ---Purpose : Explores an entity, to take its faces
    --           Works recursively
    
    ExploreLabel (me) returns AsciiString from TCollection;
    ---Purpose : Returns a text defining the criterium : "Assembly structures"

end SelectAssembly;
