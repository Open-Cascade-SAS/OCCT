-- Created on: 1993-10-21
-- Created by: Jean-Louis FRENKEL
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Modified by rob Aug 20 98 : 
--               new Methods : Is3D() , AddToImmediateList (Prs)
--                            BeginDraw redefined		
--                            new field : myStrList
--               => allows users to store independant Graphic Structures
--                  which will be displayed in immediate mode when EndDraw 
--                  is applied


class PresentationManager3d from PrsMgr inherits PresentationManager from PrsMgr

    ---Purpose: A framework to manage 3D displays, graphic entities
    -- and their updates.
    -- Used in the AIS package (Application Interactive
    -- Services), to enable the advanced user to define the
    -- default display mode of a new interactive object which
    -- extends the list of signatures and types.
    -- Definition of new display types is handled by calling
    -- the presentation algorithms provided by the StdPrs package.
    
uses
    ListOfTransient      from TColStd,
    StructureManager     from Graphic3d,
    PresentableObject    from PrsMgr,
    Length,NameOfColor   from Quantity,
    Transformation       from Geom,
    NameOfMaterial     from Graphic3d,
    --NameOfMaterialPhysic from Graphic3d,
    --NameOfPhysicalMaterial  from Graphic3d,
    Presentation         from PrsMgr,
    Presentation3d       from PrsMgr,
    View                 from V3d,
    ShadingAspect        from Prs3d,
    Presentation         from Prs3d
is

    Create(aStructureManager: StructureManager from Graphic3d)
    returns mutable PresentationManager3d  from  PrsMgr;
    ---Purpose:
    -- Creates a framework to manage displays and graphic
    -- entities with the 3D view aStructureManager.
        
    Is3D(me) returns Boolean from Standard is redefined;

    Color(me: mutable; 
            aPresentableObject: mutable PresentableObject from PrsMgr;
            aColor: NameOfColor from Quantity = Quantity_NOC_YELLOW;
            aMode: Integer from Standard = 0)
    ---Purpose: Highlights the graphic object aPresentableObject in
    -- the color aColor.
    -- aPresentableObject has the display mode aMode;
    -- this has the default value of 0, that is, the wireframe display mode.
    is static;

    
    BoundBox(me: mutable; aPresentableObject: mutable PresentableObject from PrsMgr;
    	                  aMode: Integer from Standard = 0)
    ---Purpose: highlights the boundbox of the presentation 

    is static;
    
---Category: Immediate display methods.
--           

    BeginDraw(me:mutable) is redefined static;

    AddToImmediateList(me:mutable;aPrs:Presentation from Prs3d);
    ---Purpose: stores <aPrs> in a list of structure to be displayed
    --          in immediate mode. will be taken in account in EndDraw Method.
    
    EndDraw(me: mutable; theView: View from V3d; DoubleBuffer: Boolean from Standard = Standard_False)
    is redefined static;

    	    
---Category: references to other presentation.

    Connect(me: mutable; 
                aPresentableObject: PresentableObject from PrsMgr;
                anOtherObject: mutable PresentableObject from PrsMgr;
		aMode: Integer from Standard = 0;
                anOtherMode: Integer from Standard = 0)
    is static;
    
---Category: Transformation methods.

    Transform (me: mutable;  
                   aPresentableObject: PresentableObject from PrsMgr;
		   aTransformation: Transformation from Geom;
                   aMode: Integer from Standard = 0)
    ---Purpose:
    -- Sets the transformation aTransformation for the
    -- presentable object aPresentableObject.
    -- aPresentableObject has the display mode aMode;
    -- this has the default value of 0, that is, the wireframe
    -- display mode.
    is static;
        
    Place (me: mutable; aPresentableObject: PresentableObject from PrsMgr;
                        X,Y,Z: Length from Quantity;
			aMode: Integer from Standard = 0)
    ---Purpose:
    -- Sets a position to move the presentable object
    -- aPresentableObject to. This position is defined by the
    -- lengths along the x, y and z axes: X, Y and Z respectively.
    -- aPresentableObject has the display mode aMode;
    -- this has the default value of 0, that is, the wireframe display mode.
    is static;
        
    Multiply  (me: mutable;  
                   aPresentableObject: PresentableObject from PrsMgr;
		   aTransformation: Transformation from Geom;
                   aMode: Integer from Standard = 0)
    ---Purpose:
    -- Defines the transformation aTransformation for the
    -- presentable object aPresentableObject.
    -- aPresentableObject has the display mode aMode;
    -- this has the default value of 0, that is, the wireframe
    -- display mode.
    is static;
        
    Move (me: mutable; aPresentableObject: PresentableObject from PrsMgr;
                        X,Y,Z: Length from Quantity;
			aMode: Integer from Standard = 0)
    ---Purpose:
    -- Sets a position to move the presentable object
    -- aPresentableObject to. This position is defined by the
    -- lengths along the x, y and z axes: X, Y and Z respectively.
    -- aPresentableObject has the display mode aMode;
    -- this has the default value of 0, that is, the wireframe
    -- display mode.
    is static;
    
    StructureManager(me) returns mutable StructureManager from Graphic3d
    is static;
    ---C++: inline
    ---C++: return const&
    ---Purpose: Returns the structure manager.

    SetShadingAspect(me: mutable;  
                       aPresentableObject: PresentableObject from PrsMgr;
		       aColor: NameOfColor from Quantity;
		       aMaterial: NameOfMaterial from Graphic3d;
		       --aMaterial: NameOfPhysicalMaterial from Graphic3d;
		       aMode: Integer from Standard = 0)
    ---Purpose: this method will change the color and the aspect
    --          of the presentations containg shaded structures.
    is static;


    SetShadingAspect(me: mutable;  
                       aPresentableObject: PresentableObject from PrsMgr;
		       aShadingAspect: ShadingAspect from Prs3d;
		       aMode: Integer from Standard = 0)
    ---Purpose: this method will change the color and the aspect
    --          of the presentations containg shaded structures.
    is static;


    CastPresentation(me; aPresentableObject: PresentableObject from PrsMgr;
    	                 aMode: Integer from Standard = 0)
    returns  mutable Presentation3d from PrsMgr
    is static ;
    
    newPresentation(me: mutable; aPresentableObject: PresentableObject from PrsMgr) 
    returns mutable Presentation from PrsMgr
    ---Level: Internal 
    ---Purpose: Creates a new presentation in the presentation manager.
    is redefined static private;

fields

    myStructureManager : StructureManager from Graphic3d;
    myStrList          : ListOfTransient  from TColStd;
    
end PresentationManager3d from PrsMgr;
