-- Created on: 1995-01-05
-- Created by: Frederic MAUPAS
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class GeometricTool from StepToTopoDS

  ---Purpose: This class contains some algorithmic services 
  --          specific to the mapping STEP to CAS.CADE              

uses

    Tool         from StepToTopoDS,
    SurfaceCurve from StepGeom,
    Surface      from StepGeom,
    Pcurve       from StepGeom,
    EdgeLoop     from StepShape,    
    Edge         from StepShape,    
    Curve        from Geom2d,
    Line         from Geom2d,
    Curve        from Geom,
    Surface      from Geom,
    Pnt2d        from gp,
    Pnt          from gp,
    Face         from TopoDS,
    Wire         from TopoDS,
    Edge         from TopoDS,
    Vertex       from TopoDS
    
is

    PCurve(myclass;
 	      SC : SurfaceCurve from StepGeom;
    	      S  : Surface      from StepGeom;
	      PC : out Pcurve   from StepGeom;
	      last : Integer = 0)
    	returns Integer;

    IsSeamCurve(myclass;
    	    	SC : SurfaceCurve from StepGeom;
    	      	S  : Surface      from StepGeom;
		E  : Edge         from StepShape;
    	    	EL : EdgeLoop     from StepShape)
    	returns Boolean;

		
    IsLikeSeam(myclass;
    	       SC : SurfaceCurve from StepGeom;
       	       S  : Surface      from StepGeom;
	       E  : Edge         from StepShape;
    	       EL : EdgeLoop     from StepShape)
    	returns Boolean;


    UpdateParam3d(myclass; C  : Curve from Geom;
    	    	  w1, w2 : in out Real from Standard;
		  preci  : Real)
    	returns Boolean;
			 
end GeometricTool from StepToTopoDS;
