-- Created on: 1997-09-11
-- Created by: Philippe MANGIN
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class SmoothCriterion from AppDef
inherits  TShared  from MMgt

	---Purpose: defined criterion to smooth  points in  curve
                             

uses
   Vector  from  math, 
   Matrix  from  math, 
   Curve   from  FEmTool, 
   HAssemblyTable    from  FEmTool,  
   HArray2OfInteger  from TColStd, 
   HArray1OfReal    from TColStd,
   Array1OfReal    from TColStd 
    
raises 
  NotImplemented,   
  DomainError 
   
 

is 
    SetParameters(me  :  mutable;  Parameters  : HArray1OfReal) 
    is  deferred; 

    SetCurve(me  :  mutable;  C  :Curve from FEmTool) 
    is  deferred; 
     
    GetCurve(me;  C  :  out  Curve  from FEmTool) 
    is  deferred; 
     
    SetEstimation(me  :  mutable;  E1,  E2,  E3  :  Real)   
    is  deferred; 
     
    EstLength(me  :  mutable)   
    ---C++: return &
    returns  Real  is  deferred;     
     
    GetEstimation(me;  E1,  E2,  E3  : out Real)   
    is  deferred; 
     
    AssemblyTable(me)  
    returns HAssemblyTable  from  FEmTool   
    is  deferred; 
     
    DependenceTable(me)  
    returns  HArray2OfInteger  from TColStd   
    is  deferred;  
    
    QualityValues  (me : mutable; J1min,  J2min,  J3min  :  Real; 
    	    	    	    	  J1,  J2,  J3  :  out  Real)
    returns  Integer  is  deferred;
     
    ErrorValues(me  :  mutable;   
                MaxError,  QuadraticError,  AverageError  :  out  Real) 
    is  deferred;
     
    Hessian(me  :  mutable ;  
            Element    :  Integer; 
	    Dimension1  :  Integer; 
	    Dimension2  :  Integer;
            H  :  out  Matrix  from  math)  
     raises  DomainError -- If DependenceTable(Dimension1,Dimension2) is False 
     is  deferred;  
   
    
    Gradient(me  :  mutable;  
             Element  :  Integer; 
	     Dimension  :  Integer;
             G  :  out  Vector  from  math) 
    is  deferred; 
    
    InputVector(me  :  mutable;  X : Vector from math;   
                                 AssTable  :  HAssemblyTable  from  FEmTool)  
    ---Purpose: Convert the assembly Vector in an Curve;
    --          
    raises  DomainError  is  deferred; 
     
    SetWeight(me:  mutable;  
              QuadraticWeight,  QualityWeight  :  Real; 
	      percentJ1,  percentJ2,  percentJ3  :  Real) 
    is  deferred;  
     
    GetWeight(me;  QuadraticWeight,  QualityWeight  :  out  Real)  
    is  deferred;  
     
    SetWeight(me:  mutable;  
              Weight  :  Array1OfReal)
    is  deferred;
          
end SmoothCriterion;


