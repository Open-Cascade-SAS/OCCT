-- Created on: 1995-07-18
-- Created by: Modelistation
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class   GenLocateExtPS from Extrema
					 
    	---Purpose: With a close point, it calculates the distance 
    	--          between a point and a surface.
    	--          This distance can be a minimum or a maximum.

uses    POnSurf from Extrema,
        Pnt     from gp,
	Surface from Adaptor3d
 
raises  DomainError from Standard,
    	NotDone     from StdFail


is
    Create returns GenLocateExtPS;

    Create (P: Pnt; S: Surface from Adaptor3d; U0,V0: Real; TolU,TolV: Real)
    	returns GenLocateExtPS
    	---Purpose: Calculates the distance with a close point.
    	--          The close point is defined by the parameter values
    	--          U0 and V0.
    	--          The function F(u,v)=distance(S(u,v),p) has an
    	--          extremun when gradient(F)=0. The algorithm searchs
    	--          a zero near the close point.
    	raises  DomainError;
	    	-- if U0,V0 are outside the definition ranges of the 
	    	-- surface.
    
    IsDone (me) returns Boolean
    	---Purpose: Returns True if the distance is found.
    	is static;

    SquareDistance (me) returns Real
    	---Purpose: Returns the value of the extremum square distance.
    	raises  NotDone from StdFail
	    	-- if IsDone(me)=False.
    	is static;

    Point (me) returns POnSurf
        ---C++: return const &
    	---Purpose: Returns the point of the extremum distance.
    	raises  NotDone from StdFail
	    	-- if IsDone(me)=False.
    	is static;

fields
    myDone : Boolean;
    mySqDist: Real;
    myPoint: POnSurf from Extrema;

end GenLocateExtPS;
