-- Created on: 1992-08-20
-- Created by: Christophe MARION
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Coincidence from HLRAlgo

	---Purpose: The Coincidence class is used in an Inteference to
	--          store informations on the "hiding" edge.
	--          
	--          2D  Data : The  tangent  and the  curvature of the
	--          projection of the edge  at the intersection point.
	--          This is necesserary  when the intersection  is  at
	--          the extremity of the edge.
	--          
	--          3D   Data  :  The   state of  the   edge  near the
	--          intersection   with  the face (before  and after).
	--          This is necessary  when the  intersection is  "ON"
	--          the face.

uses
    Integer from Standard,
    Real    from Standard,
    State   from TopAbs

is
    Create returns Coincidence from HLRAlgo;
    
    Set2D(me : in out; FE    : Integer from Standard;
                       Param : Real    from Standard)
    	---C++: inline
    is static;
    
    SetState3D(me : in out; stbef,staft : State from TopAbs)
    	---C++: inline
    is static;

    Value2D(me; FE    : out Integer from Standard;
                Param : out Real    from Standard)
    	---C++: inline
    is static;
    
    State3D(me; stbef,staft : out State from TopAbs)
    	---C++: inline
    is static;
	    
fields
    myFE    : Integer from Standard;
    myParam : Real    from Standard;
    myStBef : State from TopAbs;
    myStAft : State from TopAbs;

end Coincidence;
