-- Created on: 1995-05-29
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class PntFace from LocOpe

	---Purpose: 

uses Pnt         from gp,
     Face        from TopoDS,
     Orientation from TopAbs
     

is

    Create
	---Purpose: Empty constructor. Useful only for the list.
    	returns PntFace from LocOpe;


    Create (P: Pnt from gp; F: Face from TopoDS;
            Or: Orientation from TopAbs; Param,UPar,VPar: Real from Standard) 
	    
    	returns PntFace from LocOpe;
	---C++: inline

    Pnt(me)
    
    	returns Pnt from gp
	---C++: return const&
	---C++: inline
	is static;


    Face(me)
    
    	returns Face from TopoDS
	---C++: return const&
	---C++: inline
	is static;

    Orientation(me)
    
    	returns Orientation from TopAbs
	---C++: inline
	is static;


    ChangeOrientation(me: in out)
    
    	returns Orientation from TopAbs
	---C++: return &
	---C++: inline
	is static;


    Parameter(me)
    
    	returns Real from Standard
	---C++: inline
	is static;


    UParameter(me)
    
    	returns Real from Standard
	---C++: inline
	is static;


    VParameter(me)
    
    	returns Real from Standard
	---C++: inline
	is static;


fields

    myPnt  : Pnt         from gp;
    myFace : Face        from TopoDS;
    myOri  : Orientation from TopAbs;
    myPar  : Real        from Standard;
    myUPar : Real        from Standard;
    myVPar : Real        from Standard;

end PntFace;
