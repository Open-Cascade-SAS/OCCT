-- Created on: 1998-09-23
-- Created by: Philippe MANGIN
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



private  class LogSample from GeomLib inherits FunctionSample  from  math

	---Purpose: 
raises 
   OutOfRange  from  Standard
is 
 
  Create(A,B: Real; N: Integer)
  returns LogSample from GeomLib; 
   
  GetParameter(me; Index: Integer)
    
	---Purpose: Returns the value of parameter of the point of 
	--          range Index : A + ((Index-1)/(NbPoints-1))*B.
	--          An exception is raised if Index<=0 or Index>NbPoints.

    returns Real
    raises OutOfRange
    is redefined;

fields 
  myF    :  Real; 
  myexp  :  Real;

end LogSample;
