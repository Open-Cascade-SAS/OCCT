-- Created on: 2000-05-10
-- Created by: Andrey BETENEV
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1

class RoleSelect from StepBasic
inherits SelectType from StepData

    ---Purpose: Representation of STEP SELECT type RoleSelect

uses
    ActionAssignment from StepBasic,
    ActionRequestAssignment from StepBasic,
    ApprovalAssignment from StepBasic,
    ApprovalDateTime from StepBasic,
    CertificationAssignment from StepBasic,
    ContractAssignment from StepBasic,
    DocumentReference from StepBasic,
    EffectivityAssignment from StepBasic,
    GroupAssignment from StepBasic,
    NameAssignment from StepBasic,
    SecurityClassificationAssignment from StepBasic

is
    Create returns RoleSelect from StepBasic;
	---Purpose: Empty constructor

    CaseNum (me; ent: Transient) returns Integer;
	---Purpose: Recognizes a kind of RoleSelect select type
	--          1 -> ActionAssignment from StepBasic
	--          2 -> ActionRequestAssignment from StepBasic
	--          3 -> ApprovalAssignment from StepBasic
	--          4 -> ApprovalDateTime from StepBasic
	--          5 -> CertificationAssignment from StepBasic
	--          6 -> ContractAssignment from StepBasic
	--          7 -> DocumentReference from StepBasic
	--          8 -> EffectivityAssignment from StepBasic
	--          9 -> GroupAssignment from StepBasic
	--          10 -> NameAssignment from StepBasic
	--          11 -> SecurityClassificationAssignment from StepBasic
	--          0 else

    ActionAssignment (me) returns ActionAssignment from StepBasic;
	---Purpose: Returns Value as ActionAssignment (or Null if another type)

    ActionRequestAssignment (me) returns ActionRequestAssignment from StepBasic;
	---Purpose: Returns Value as ActionRequestAssignment (or Null if another type)

    ApprovalAssignment (me) returns ApprovalAssignment from StepBasic;
	---Purpose: Returns Value as ApprovalAssignment (or Null if another type)

    ApprovalDateTime (me) returns ApprovalDateTime from StepBasic;
	---Purpose: Returns Value as ApprovalDateTime (or Null if another type)

    CertificationAssignment (me) returns CertificationAssignment from StepBasic;
	---Purpose: Returns Value as CertificationAssignment (or Null if another type)

    ContractAssignment (me) returns ContractAssignment from StepBasic;
	---Purpose: Returns Value as ContractAssignment (or Null if another type)

    DocumentReference (me) returns DocumentReference from StepBasic;
	---Purpose: Returns Value as DocumentReference (or Null if another type)

    EffectivityAssignment (me) returns EffectivityAssignment from StepBasic;
	---Purpose: Returns Value as EffectivityAssignment (or Null if another type)

    GroupAssignment (me) returns GroupAssignment from StepBasic;
	---Purpose: Returns Value as GroupAssignment (or Null if another type)

    NameAssignment (me) returns NameAssignment from StepBasic;
	---Purpose: Returns Value as NameAssignment (or Null if another type)

    SecurityClassificationAssignment (me) returns SecurityClassificationAssignment from StepBasic;
	---Purpose: Returns Value as SecurityClassificationAssignment (or Null if another type)

end RoleSelect;
