-- Created on: 1996-04-09
-- Created by: Joelle CHAUVET
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Node from AdvApp2Var


uses
    XY,Pnt           from gp,
    HArray2OfPnt     from TColgp,
    HArray2OfReal    from TColStd
    
	 
is
    Create returns Node;    
    Create(iu,iv : Integer) returns Node;   
    Create(UV : XY from gp; iu,iv : Integer) returns Node;    
    Create(Other : Node) returns Node is private;    
    Coord(me) returns XY from gp;    
    SetCoord(me : in out; x1,x2 : Real);    
    UOrder(me) returns Integer;
    VOrder(me) returns Integer;
    SetPoint(me : in out; iu,iv : Integer; Cte : Pnt from gp);    
    Point(me; iu,iv : Integer) returns Pnt from gp;    
    SetError(me : in out; iu,iv : Integer; error : Real);    
    Error(me; iu,iv : Integer) returns Real;     
    
    
fields

    myCoord            : XY               from gp;
    myOrdInU, myOrdInV : Integer;
    myTruePoints       : HArray2OfPnt     from TColgp;
    myErrors           : HArray2OfReal    from TColStd;
    
end Node;







