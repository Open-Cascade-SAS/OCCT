-- Created on: 1992-10-20
-- Created by: Remi GILET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Circ2dTanOnRad from Geom2dGcc

	---Purpose: This class implements the algorithms used to 
	--          create a 2d circle tangent to a 2d entity, 
	--          centered on a 2d entity and with a given radius.
	--          More than one argument must be a curve.
	--          The arguments of all construction methods are :
	--             - The qualified element for the tangency constrains 
	--             (QualifiedCirc, QualifiedLin, QualifiedCurvPoints).
	--             - The Center element (circle, line, curve).
	--             - A real Tolerance.
	--          Tolerance is only used in the limits cases.
    	--          For example : 
    	--          We want to create a circle tangent to an OutsideCurv Cu1
    	--          centered on a line OnLine with a radius Radius and with
    	--          a tolerance Tolerance.
    	--          If we did not used Tolerance it is impossible to 
    	--          find a solution in the the following case : OnLine is 
    	--          outside Cu1. There is no intersection point between Cu1
    	--          and OnLine. The distance between the line and the 
    	--          circle is greater than Radius.
    	--          With Tolerance we will give a solution if the 
    	--          distance between Cu1 and OnLine is lower than or 
    	--          equal Tolerance.

-- inherits Entity from Standard

uses Lin2d            from gp, 
     Circ2d           from gp,  
     Pnt2d            from gp,
     Point            from Geom2d,
     Array1OfCirc2d   from TColgp,
     Array1OfPnt2d    from TColgp,
     Curve            from Geom2dAdaptor,
     QualifiedCurve   from Geom2dGcc,
     Array1OfReal     from TColStd,
     Array1OfInteger  from TColStd,
     Circ2dTanOnRad   from GccAna,
     MyCirc2dTanOnRad from Geom2dGcc,
     Position         from GccEnt,
     Array1OfPosition from GccEnt
     
raises NegativeValue from Standard,
       OutOfRange    from Standard,
       BadQualifier  from GccEnt,
       NotDone       from StdFail

is

Create(Qualified1 :  QualifiedCurve from Geom2dGcc    ;
       OnCurv     :  Curve          from Geom2dAdaptor;
       Radius     :  Real           from Standard     ;
       Tolerance  :  Real           from Standard     )
returns Circ2dTanOnRad from Geom2dGcc
raises NegativeValue,BadQualifier;
    	---Purpose: Constructs one or more 2D circles of radius Radius,
    	-- centered on the 2D curve OnCurv and:
    	-- -   tangential to the curve Qualified1
        
Create(Point1     :  Point  from Geom2d       ;
       OnCurv     :  Curve  from Geom2dAdaptor;
       Radius     :  Real   from Standard     ;
       Tolerance  :  Real   from Standard     ) 
returns Circ2dTanOnRad from Geom2dGcc
raises NegativeValue;
    	---Purpose: Constructs one or more 2D circles of radius Radius,
    	-- centered on the 2D curve OnCurv and:
    	-- passing through the point Point1.
    	--  OnCurv is an adapted curve, i.e. an object which is an
    	-- interface between:
    	-- -   the services provided by a 2D curve from the package Geom2d,
    	-- -   and those required on the curve by the construction algorithm.
    	-- Similarly, the qualified curve Qualified1 is created from
    	-- an adapted curve.
    	-- Adapted curves are created in the following way:
    	-- Handle(Geom2d_Curve) myCurveOn = ... ;
    	-- Geom2dAdaptor_Curve OnCurv ( myCurveOn ) ;
    	-- The algorithm is then constructed with this object:
    	-- Handle(Geom2d_Curve) myCurve1 = ...
    	-- ;
    	-- Geom2dAdaptor_Curve Adapted1 ( myCurve1 ) ;
	-- Geom2dGcc_QualifiedCurve
    	--           Qualified1 = Geom2dGcc::Outside(Adapted1);
    	-- Standard_Real Radius = ... , Tolerance = ... ;
    	-- Geom2dGcc_Circ2dTanOnRad
    	--             myAlgo ( Qualified1 , OnCurv , Radius , Tolerance ) ;
    	-- if ( myAlgo.IsDone() )
    	--     { Standard_Integer Nbr = myAlgo.NbSolutions() ;
    	--     gp_Circ2d Circ ;
    	--     for ( Standard_Integer i = 1 ;
    	-- i <= nbr ; i++ )
    	--        { Circ = myAlgo.ThisSolution (i) ;
    	--           ...
    	--        }
    	--     }

Results(me   : in out                         ;
    	Circ :        Circ2dTanOnRad from GccAna)
is static;

Results(me   : in out                              ;
    	Circ :        MyCirc2dTanOnRad from Geom2dGcc)
is static;

IsDone(me) returns Boolean from Standard
is static;
    	---Purpose: Returns true if the construction algorithm does not fail
    	-- (even if it finds no solution).
    	-- Note: IsDone protects against a failure arising from a
    	-- more internal intersection algorithm which has reached
    	-- its numeric limits.
NbSolutions(me) returns Integer from Standard
raises NotDone
is static;
    	---Purpose: Returns the number of circles, representing solutions
    	-- computed by this algorithm.
    	-- Exceptions: StdFail_NotDone if the construction fails.
    
ThisSolution(me ; Index : Integer from Standard) returns Circ2d from gp 
raises OutOfRange, NotDone
is static;
	---Purpose: Returns the solution number Index and raises OutOfRange 
    	-- exception if Index is greater than the number of solutions.
    	-- Be carefull: the Index is only a way to get all the 
    	-- solutions, but is not associated to theses outside the context
    	-- of the algorithm-object.
    	-- Exceptions
    	-- Standard_OutOfRange if Index is less than zero or
    	-- greater than the number of solutions computed by this algorithm.
    	-- StdFail_NotDone if the construction fails.
        
WhichQualifier(me                                  ;
    	       Index   :     Integer  from Standard;
	       Qualif1 : out Position from GccEnt  )
raises OutOfRange, NotDone
is static;
    	--- Purpose: Returns the qualifier Qualif1 of the tangency argument
    	-- for the solution of index Index computed by this algorithm.
    	-- The returned qualifier is:
    	-- -   that specified at the start of construction when the
    	--   solutions are defined as enclosed, enclosing or
    	--   outside with respect to the arguments, or
    	-- -   that computed during construction (i.e. enclosed,
    	--   enclosing or outside) when the solutions are defined
    	--   as unqualified with respect to the arguments, or
    	-- -   GccEnt_noqualifier if the tangency argument is a point.
    	--  Exceptions
    	-- Standard_OutOfRange if Index is less than zero or
    	-- greater than the number of solutions computed by this algorithm.
    	-- StdFail_NotDone if the construction fails.

Tangency1(me                                     ;
          Index         : Integer   from Standard;
          ParSol,ParArg : out Real  from Standard;
          PntSol        : out Pnt2d from gp      )
raises OutOfRange, NotDone
is static;
    	---Purpose: Returns informations about the tangency point between the 
    	-- result number Index and the first argument.
	-- ParSol is the intrinsic parameter of the point on the solution curv.
	-- ParArg is the intrinsic parameter of the point on the argument curv.
    	-- PntSol is the tangency point on the solution curv.
    	-- PntArg is the tangency point on the argument curv.
    	-- Exceptions
    	-- Standard_OutOfRange if Index is less than zero or
    	-- greater than the number of solutions computed by this algorithm.
    	-- StdFail_NotDone if the construction fails.
        
CenterOn3 (me                                     ;
           Index         : Integer   from Standard;
           ParArg        : out Real  from Standard;
           PntSol        : out Pnt2d from gp      )
raises OutOfRange, NotDone
is static;
    	---Purpose: Returns the center PntSol on the second argument (i.e.
    	-- line or circle) of the solution of index Index computed by
    	-- this algorithm.
    	-- ParArg is the intrinsic parameter of the point on the argument curv.
    	-- PntSol is the center point of the solution curv.
    	-- PntArg is the projection of PntSol on the argument curv.
    	-- Exceptions:
    	-- Standard_OutOfRange if Index is less than zero or
    	-- greater than the number of solutions computed by this algorithm.
    	-- StdFail_NotDone if the construction fails.
        
IsTheSame1(me                            ;
           Index : Integer  from Standard) returns Boolean from Standard
raises OutOfRange, NotDone
is static;
    	---Purpose: Returns true if the solution of index Index and the first
    	-- argument of this algorithm are the same (i.e. there are 2
    	-- identical circles).
    	-- If Rarg is the radius of the first argument, Rsol is the
    	-- radius of the solution and dist is the distance between
    	-- the two centers, we consider the two circles to be
    	-- identical if |Rarg - Rsol| and dist are less than
    	-- or equal to the tolerance criterion given at the time of
    	-- construction of this algorithm.
    	-- OutOfRange is raised if Index is greater than the number of solutions.
    	-- notDone is raised if the construction algorithm did not succeed.

fields

    WellDone : Boolean from Standard;
    -- True if the algorithm succeeded.

    NbrSol   : Integer from Standard;
    -- The number of possible solutions. We have to decide about the
    -- status of the multiple solutions...

    cirsol   : Array1OfCirc2d from TColgp;
    ---Purpose : The solutions.

    qualifier1 : Array1OfPosition from GccEnt;
    -- The qualifiers of the first argument.

    TheSame1 : Array1OfInteger from TColStd;

    pnttg1sol   : Array1OfPnt2d from TColgp;
    -- The tangency point between the solution and the first argument on 
    -- the solution.

    par1sol   : Array1OfReal from TColStd;
    -- The parameter of the tangency point between the solution and the 
    -- first argument on the solution.

    pararg1   : Array1OfReal from TColStd;
    -- The parameter of the tangency point between the solution and the first 
    -- argument on the first argument.

    pntcen3   : Array1OfPnt2d from TColgp;
    -- The center point of the solution on the first argument.

    parcen3   : Array1OfReal from TColStd;
    -- The parameter of the center point of the solution on the second 
    -- argument.

end Circ2dTanOnRad;


