-- Created on: 1998-06-03
-- Created by: data exchange team
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class EdgeProjAux from ShapeFix inherits TShared from MMgt

    ---Purpose: Project 3D point (vertex) on pcurves to find Vertex Parameter
    --          on parametric representation of an edge

uses

    Curve   from Geom2d,
    Face    from TopoDS,
    Edge    from TopoDS,
    Surface from Geom
    
is

    Create returns mutable EdgeProjAux from ShapeFix;

    Create (F: Face from TopoDS; E: Edge from TopoDS)
    returns mutable EdgeProjAux from ShapeFix;
    
    Init (me: mutable; F: Face from TopoDS; E: Edge from TopoDS);

    Compute (me: mutable; preci: Real);

    IsFirstDone (me) returns Boolean from Standard;

    IsLastDone (me) returns Boolean from Standard;

    FirstParam (me) returns Real from Standard;

    LastParam (me) returns Real from Standard;

    IsIso (me: mutable; C: Curve from Geom2d) returns Boolean;

    Init2d (me: mutable; preci: Real) is protected;

    Init3d (me: mutable; preci: Real) is protected;

    UpdateParam2d (me: mutable; C: Curve from Geom2d) is protected;

fields

    myFace: Face from TopoDS is protected;
    myEdge: Edge from TopoDS is protected;
    myFirstParam: Real is protected;
    myLastParam: Real is protected;
    myFirstDone: Boolean is protected;
    myLastDone: Boolean is protected;
    
end EdgeProjAux;
