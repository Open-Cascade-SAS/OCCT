-- File:	RWStepBasic_RWNameAssignment.cdl
-- Created:	Wed May 10 15:09:08 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class RWNameAssignment from RWStepBasic

    ---Purpose: Read & Write tool for NameAssignment

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    NameAssignment from StepBasic

is
    Create returns RWNameAssignment from RWStepBasic;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : NameAssignment from StepBasic);
	---Purpose: Reads NameAssignment

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: NameAssignment from StepBasic);
	---Purpose: Writes NameAssignment

    Share (me; ent : NameAssignment from StepBasic;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWNameAssignment;
