-- File:        Path.cdl
-- Created:     Fri Dec  1 11:11:23 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class Path from StepShape 

inherits TopologicalRepresentationItem from StepShape 

uses

	HArray1OfOrientedEdge from StepShape, 
	OrientedEdge from StepShape, 
	HAsciiString from TCollection
is

	Create returns mutable Path;
	---Purpose: Returns a Path


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aEdgeList : mutable HArray1OfOrientedEdge from StepShape) is virtual;

	-- Specific Methods for Field Data Access --

	SetEdgeList(me : mutable; aEdgeList : mutable HArray1OfOrientedEdge)
    	is virtual;
	EdgeList (me) returns mutable HArray1OfOrientedEdge
    	is virtual;
	EdgeListValue (me; num : Integer) returns mutable OrientedEdge
    	is virtual;
	NbEdgeList (me) returns Integer
    	is virtual;

fields

	edgeList : HArray1OfOrientedEdge from StepShape;

end Path;
