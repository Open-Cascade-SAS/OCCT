-- File:	TopoDSToStep_MakeFacetedBrepAndBrepWithVoids.cdl
-- Created:	Fri Jul 23 15:09:44 1993
-- Author:	Martine LANGLOIS
--		<mla@mastox>
---Copyright:	 Matra Datavision 1993

class MakeFacetedBrepAndBrepWithVoids from TopoDSToStep inherits
    Root from TopoDSToStep

    ---Purpose: This class implements the mapping between classes 
    --          Solid from TopoDS and FacetedBrepAndBrepWithVoids from
    --          StepShape. All the topology and geometry comprised 
    --          into the shell or the solid are taken into account and
    --          translated.
  
uses Solid from TopoDS,
     FacetedBrepAndBrepWithVoids from StepShape,
     FinderProcess from Transfer
          
raises NotDone from StdFail
     
is 

Create ( S  : Solid from TopoDS;
         FP : mutable FinderProcess from Transfer)
        returns MakeFacetedBrepAndBrepWithVoids;

Value (me) returns FacetedBrepAndBrepWithVoids from StepShape
    raises NotDone
    is static;
    ---C++: return const&

fields

    theFacetedBrepAndBrepWithVoids : FacetedBrepAndBrepWithVoids from StepShape;

    	-- The solution from StepShape
    	
end MakeFacetedBrepAndBrepWithVoids;


