-- File:	Prs3d_WFDeflectionRestrictedFace.cdl
-- Created:	Mon Jan 18 18:27:19 1993
-- Author:	Jean Louis FRENKEL
--		<jlf@mastox>
---Copyright:	 Matra Datavision 1993

generic class WFDeflectionRestrictedFace from Prs3d 
          (DrawFaceIso     as any;
    	   RestrictionTool as any)
	  
inherits Root from Prs3d
	 

	---Purpose: 

uses
    HSurface             from BRepAdaptor,
    Presentation         from Prs3d,
    Drawer               from Prs3d,
    Length               from Quantity, 
    NListOfSequenceOfPnt from Prs3d

    
is
    Add(myclass; aPresentation: Presentation from Prs3d; 
        	 aFace        : HSurface     from BRepAdaptor;
    	    	 aDrawer      : Drawer       from Prs3d);
		 
    AddUIso(myclass; aPresentation: Presentation from Prs3d; 
        	     aFace        : HSurface     from BRepAdaptor;
    	    	     aDrawer      : Drawer       from Prs3d);
		 
    AddVIso(myclass; aPresentation: Presentation from Prs3d; 
        	     aFace        : HSurface     from BRepAdaptor;
    	    	     aDrawer      : Drawer       from Prs3d);
		 
    Add(myclass;  aPresentation: Presentation from Prs3d; 
    	          aFace        : HSurface     from BRepAdaptor;
		  DrawUIso, DrawVIso: Boolean from Standard;
		  Deflection   : Length       from Quantity;
		  NBUiso,NBViso: Integer      from Standard;
		  aDrawer      : Drawer       from Prs3d; 
    	    	  Curves       : out NListOfSequenceOfPnt from Prs3d);

		   
    Match(myclass; X,Y,Z    : Length   from Quantity;
                   aDistance: Length   from Quantity;
        	   aFace    : HSurface from BRepAdaptor;
    	    	   aDrawer  : Drawer   from Prs3d)
    returns Boolean from Standard;
		 
    MatchUIso(myclass; X,Y,Z    : Length   from Quantity;
                       aDistance: Length   from Quantity;
        	       aFace    : HSurface from BRepAdaptor;
    	    	       aDrawer  : Drawer   from Prs3d)
    returns Boolean from Standard;
		 
    MatchVIso(myclass; X,Y,Z    : Length   from Quantity;
                       aDistance: Length   from Quantity;
         	       aFace    : HSurface from BRepAdaptor;
    	    	       aDrawer  : Drawer   from Prs3d)
    returns Boolean from Standard;
		 

    Match(myclass;X,Y,Z        : Length       from Quantity;
                  aDistance    : Length       from Quantity;
    	          aFace        : HSurface     from BRepAdaptor; 
    	    	  aDrawer      : Drawer       from Prs3d;
		  DrawUIso, DrawVIso: Boolean from Standard;
		  aDeflection  : Length       from Quantity;
		  NBUiso,NBViso: Integer      from Standard)

    returns Boolean from Standard;	  
		   
end WFDeflectionRestrictedFace;

