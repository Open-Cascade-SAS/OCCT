-- Created on: 2005-10-14
-- Created by: Mikhail KLOKOV
-- Copyright (c) 2005-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class CurveRangeLocalizeData from IntTools
uses
    Box from Bnd,
    CurveRangeSample from IntTools,
    MapOfCurveSample from IntTools,
    ListOfCurveRangeSample from IntTools,
    DataMapOfCurveSampleBox from IntTools

is
    Create(theNbSample: Integer from Standard;
    	   theMinRange: Real from Standard)
    	returns CurveRangeLocalizeData from IntTools;

    GetNbSample(me)
    	returns Integer from Standard;
	---C++: inline

    GetMinRange(me)
    	returns Real from Standard;
	---C++: inline

    AddOutRange(me: in out; theRange: CurveRangeSample from IntTools);
    
    AddBox(me: in out; theRange: CurveRangeSample from IntTools;
    	    	       theBox: Box from Bnd);

    FindBox(me; theRange: CurveRangeSample from IntTools;
    	    	theBox: out Box from Bnd)
    	returns Boolean from Standard;

    IsRangeOut(me; theRange: CurveRangeSample from IntTools)
    	returns Boolean from Standard;

    ListRangeOut(me; theList: out ListOfCurveRangeSample from IntTools);

fields
    myNbSampleC: Integer from Standard;
    myMinRangeC: Real from Standard;
    myMapRangeOut: MapOfCurveSample from IntTools;
    myMapBox      : DataMapOfCurveSampleBox from IntTools;

end CurveRangeLocalizeData from IntTools;
