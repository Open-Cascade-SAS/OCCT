-- Created on: 1993-10-08
-- Created by: Gilles DEBARBOUILLE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

private class UnitsLexicon from Units 

inherits

    Lexicon from Units
	---Purpose: This class defines a lexicon useful to analyse and
	--          recognize the different key  words  included  in a
	--          sentence. The  lexicon is stored  in a sequence of
	--          tokens.

uses

    HAsciiString from TCollection,
    AsciiString  from TCollection


is

    Create returns UnitsLexicon from Units;
    
    ---Level: Internal 
    
    ---Purpose: Returns an empty instance of UnitsLexicon
    
    Creates(me : mutable ; afilename1 , afilename2 : CString ;
                 amode : Boolean = Standard_True)
    
    ---Level: Internal 
    
    ---Purpose: Reads  the files  <afilename1>  and  <afilename2>   to
    --          create     a   sequence     of    tokens   stored   in
    --          <thesequenceoftokens>.
    
    is static;
    
    FileName2(me) returns AsciiString from TCollection
    
    ---Level: Internal 
    
    ---Purpose: Returns in a AsciiString from TCollection the name of the file.
    
    is static;
    
    UpToDate(me) returns Boolean
    
    ---Level: Internal 
    
    ---Purpose: Returns true if  the  file has not  changed  since the
    --          creation   of   the  Lexicon   object.   Returns false
    --          otherwise.
    
    is redefined;
    
    Dump(me)
    
    ---Level: Internal 
    
    ---C++: inline
    ---Purpose: Useful for debugging.
    
    is redefined;

fields

    thefilename     : HAsciiString from TCollection;
    thetime         : Time from Standard;

end UnitsLexicon;
