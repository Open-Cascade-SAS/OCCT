-- Created on: 1998-03-24
-- Created by: # Andre LIEUTIER
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class LinearXYZConstraint from Plate
---Purpose : define on or several constraints as linear combination of
--         PinPointConstraint unlike the LinearScalarConstraint, usage
--         of this kind of constraint preserve the X,Y and Z uncoupling.

uses 
   XY from gp, 
   XYZ from gp, 
   PinpointConstraint  from  Plate,
   Array1OfPinpointConstraint  from  Plate,
   HArray1OfPinpointConstraint  from  Plate,
   Array1OfReal from TColStd,
   Array2OfReal from TColStd,
   HArray2OfReal from TColStd
         
raises
    DimensionMismatch from Standard,
    OutOfRange from Standard
   
is
    Create returns LinearXYZConstraint; 
    
    Create  (PPC  :  Array1OfPinpointConstraint; coeff  :  Array1OfReal )
           returns LinearXYZConstraint 
	   raises DimensionMismatch from Standard;
    --  the length of PPC  have to be the  Row lentgth of  coeff
    --  
    Create  (PPC  :  Array1OfPinpointConstraint; coeff  :  Array2OfReal )
           returns LinearXYZConstraint 
	   raises DimensionMismatch from Standard;
    --  the length of PPC  have to be the  Row lentgth of  coeff

    Create  (ColLen,RowLen  :  Integer ) 
    -- initialize with 0 valued PPC and Coeffs
           returns LinearXYZConstraint;

     -- Accessors :
    GetPPC(me) returns Array1OfPinpointConstraint;
    ---C++: inline 
    ---C++: return  const &

    Coeff(me) returns Array2OfReal;
    ---C++: inline 
    ---C++: return  const &

    SetPPC (me : in out;  
    	Index: Integer from Standard;  
    	Value: PinpointConstraint) 
    	---Purpose:  Sets   the PinPointConstraint of   index Index to
    	--          Value raise if Index is greater than the length of
    	--          PPC or the Row length of coeff or lower  than 1
    	raises OutOfRange from Standard;

    SetCoeff (me : in out;  
    	Row, Col: Integer from Standard;  
    	Value: Real) 
    	---Purpose:  Sets the coeff  of index (Row,Col)  to Value 
    	--           raise if  Row (respectively Col)  is greater than the
    	--          Row (respectively Column) length of coeff
    	raises OutOfRange from Standard;

fields
    
    myPPC  :  HArray1OfPinpointConstraint;
    myCoef :  HArray2OfReal;

end;
