-- Created on: 1992-01-21
-- Created by: GG
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Update: 	FDA Oct 15 1994, 
--		ZOV - Mars 30 1998


class AmbientLight from V3d

    	---Purpose: Creation of an ambient light source in a viewer.


inherits Light from V3d

uses 

	Viewer from V3d,
        TypeOfRepresentation from V3d,
	NameOfColor from Quantity,
	View from V3d,
	Coordinate from V3d,
	Structure from Graphic3d,
	Vertex from Graphic3d,
	Group from Graphic3d

is

    	Create ( VM : mutable Viewer ;
		 Color : NameOfColor = Quantity_NOC_WHITE ) 
				returns mutable AmbientLight;
	---Purpose: Constructs an ambient light source in the viewer VM.
    	-- The default Color of this light source is WHITE.

end AmbientLight;
