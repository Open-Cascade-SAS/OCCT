-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Strips from Graphic3d

uses

	Array1OfInteger from TColStd,
	SequenceOfInteger from TColStd

is

	STRIPT_INIT (myclass; NBVERTICES: Integer; TABTRIANGLES: Array1OfInteger from TColStd);
	STRIPT_GET_STRIP(myclass; NBTRIANGLES, V1, V2: out Integer);
	STRIPT_GET_VERTEX(myclass; VERTEX, TRIANGLE: out Integer);
	STRIPQ_INIT(myclass; NBVERTICES, NBQUADRANG: Integer; TABQUADRANGLES: SequenceOfInteger from TColStd);
	STRIPQ_GET_STRIP(myclass; NBQUAD, V1, V2: out Integer);
	STRIPQ_GET_NEXT(myclass; VERTEX1, VERTEX2, QUADRANGLE: out Integer);

end Strips;
