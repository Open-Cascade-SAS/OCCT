-- Created on: 1991-06-27
-- Created by: Remi LEQUETTE
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package BRep 

	---Purpose: This package describes  a Boundary  Representation
	--          Data   Structure   inherited  from   the  abstract
	--          Topology   defined  in the   TopoDS  package.  The
	--          geometric data are provided by the Geom and Geom2d
	--          packages.
	--          
	--          The TVertex,  TEdge,  and TFace  are  redefined in
	--          this package to add geometric information.

        ---Level : Public  
        --  All methods of all  classes will be public.

uses
    MMgt,        -- Memory management
    TCollection, -- Basic data structures
    TColStd,     -- HArray1OfInteger
    gp,          -- Elementary geometry
    Bnd,         -- Bounding boxes
    TopLoc,      -- Local coordinate systems
    TopAbs,      -- Enumerations : Orientation, ShapeType
    TopoDS,      -- Abstract topological data structure
    GeomAbs,     -- Enumerations : Shape
    Geom,        -- 3D geometry : curves and surfaces
    Geom2d,      -- 2D geometry : curves in parametric space
    Poly         -- Triangulations and Polygons

is

    --
    --  Face
    --  

    class TFace;

    --
    --  Edge
    --
    --  An Edge is  defined by a list  of curve representations  which
    --  are either :
    --  
    --  Geometric representations :
    --  
    --  * A 3d curve (at most one)
    --  
    --  * A curve on surface, curve in parametric space.
    --  
    --  * A curve on closed surface, two curves in parametric space.
    --  
    --  Polygonal representations :
    --  
    --  * A 3d polygon (at most one).
    --  
    --  * A Polygon on triangulation (array of node indices)
    --  
    --  * A Polygon on closed triangulation (2 arrays of node indices)
    --  
    --  * A polygon on surface (array of 2d points in parametric space)
    --  
    --  Curve on 2 surfaces :
    --  
    --  * This is used for storing shape continuity.
    --  

    deferred class CurveRepresentation;

    class ListOfCurveRepresentation instantiates
    List from TCollection (CurveRepresentation from BRep);
    
    deferred class GCurve;

    class Curve3D;

    class CurveOnSurface;

    class CurveOnClosedSurface;

    class Polygon3D;

    class PolygonOnTriangulation;

    class PolygonOnClosedTriangulation;

    class PolygonOnSurface;

    class PolygonOnClosedSurface;

    class CurveOn2Surfaces;

    class TEdge;

    --
    --  Vertex
    --

    deferred class PointRepresentation;

    class ListOfPointRepresentation instantiates
    List from TCollection (PointRepresentation from BRep);
    
    class PointOnCurve;

    deferred class PointsOnSurface;

    class PointOnCurveOnSurface;

    class PointOnSurface;

    class TVertex;

    class Builder;

    class Tool;


end BRep;
