-- File:        SecurityClassification.cdl
-- Created:     Mon Dec  4 12:02:31 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWSecurityClassification from RWStepBasic

	---Purpose : Read & Write Module for SecurityClassification

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     SecurityClassification from StepBasic,
     EntityIterator from Interface

is

	Create returns RWSecurityClassification;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable SecurityClassification from StepBasic);

	WriteStep (me; SW : in out StepWriter; ent : SecurityClassification from StepBasic);

	Share(me; ent : SecurityClassification from StepBasic; iter : in out EntityIterator);

end RWSecurityClassification;
