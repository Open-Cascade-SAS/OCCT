-- Created on: 1997-02-11
-- Created by: Alexander BRIVIN
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Texture2Transform from Vrml 

	---Purpose: defines a Texture2Transform node of VRML specifying properties of geometry
	---          and its appearance.
    	--  This  node  defines  a 2D  transformation  applied  to  texture  coordinates.   
	--  This  affect  the  way  textures  are  applied  to  the  surfaces  of  subsequent 
    	--  shapes. 
    	--  Transformation  consisits  of(in  order)  a  non-uniform  scale  about  an   
    	--  arbitrary  center  point,  a  rotation  about  that  same  point,  and 
	--  a  translation.  This  allows  a  user  to  change  the  size  and  position  of 
	--  the  textures  on  the  shape.
    	--  By  default  : 
	--    myTranslation (0 0)
	--    myRotation (0)
	--    myScaleFactor (1 1)
	--    myCenter (0 0) 
 
uses
 
   Vec2d from gp 

is
 
    Create  returns  Texture2Transform from Vrml;
 
    Create  ( aTranslation  :  Vec2d   from  gp;
    	      aRotation     :  Real    from  Standard; 
    	      aScaleFactor  :  Vec2d   from  gp;
    	      aCenter       :  Vec2d   from  gp ) 
        returns  Texture2Transform from Vrml;

    SetTranslation ( me : in out; aTranslation : Vec2d  from  gp );
    Translation ( me  )  returns  Vec2d  from  gp;

    SetRotation ( me : in out; aRotation : Real from Standard );
    Rotation ( me )  returns  Real from Standard;

    SetScaleFactor( me : in out; aScaleFactor : Vec2d  from  gp );
    ScaleFactor( me )  returns  Vec2d  from  gp;

    SetCenter ( me : in out; aCenter : Vec2d  from  gp );
    Center ( me )  returns  Vec2d  from  gp;

    Print  ( me;  anOStream: in out OStream from Standard) returns OStream from Standard;
    ---C++:  return  & 

fields
 
    myTranslation  :  Vec2d  from  gp;       -- Translation vector
    myRotation     :  Real   from  Standard; -- Rotation
    myScaleFactor  :  Vec2d  from  gp;       -- Scale factors
    myCenter       :  Vec2d  from  gp;       -- Center point for scale and rotate
    
end Texture2Transform;

