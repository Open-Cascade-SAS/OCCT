-- Created on: 2000-05-11
-- Created by: data exchange team
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1

class CharacterizedDefinition from StepRepr
inherits SelectType from StepData

    ---Purpose: Representation of STEP SELECT type CharacterizedDefinition

uses
    CharacterizedObject from StepBasic,
    ProductDefinition from StepBasic,
    ProductDefinitionRelationship from StepBasic,
    ProductDefinitionShape from StepRepr,
    ShapeAspect from StepRepr,
    ShapeAspectRelationship from StepRepr,
    DocumentFile from StepBasic

is
    Create returns CharacterizedDefinition from StepRepr;
	---Purpose: Empty constructor

    CaseNum (me; ent: Transient) returns Integer;
	---Purpose: Recognizes a kind of CharacterizedDefinition select type
	--          1 -> CharacterizedObject from StepBasic
	--          2 -> ProductDefinition from StepBasic
	--          3 -> ProductDefinitionRelationship from StepBasic
	--          4 -> ProductDefinitionShape from StepRepr
	--          5 -> ShapeAspect from StepRepr
	--          6 -> ShapeAspectRelationship from StepRepr
	--          7 -> DocumentFile from StepBasic
	--          0 else

    CharacterizedObject (me) returns CharacterizedObject from StepBasic;
	---Purpose: Returns Value as CharacterizedObject (or Null if another type)

    ProductDefinition (me) returns ProductDefinition from StepBasic;
	---Purpose: Returns Value as ProductDefinition (or Null if another type)

    ProductDefinitionRelationship (me) returns ProductDefinitionRelationship from StepBasic;
	---Purpose: Returns Value as ProductDefinitionRelationship (or Null if another type)

    ProductDefinitionShape (me) returns ProductDefinitionShape from StepRepr;
	---Purpose: Returns Value as ProductDefinitionShape (or Null if another type)
 
    ShapeAspect (me) returns ShapeAspect from StepRepr;
	---Purpose: Returns Value as ShapeAspect (or Null if another type)

    ShapeAspectRelationship (me) returns ShapeAspectRelationship from StepRepr;
	---Purpose: Returns Value as ShapeAspectRelationship (or Null if another type)

    DocumentFile (me) returns DocumentFile from StepBasic;
	---Purpose: Returns Value as DocumentFile (or Null if another type)

end CharacterizedDefinition;
