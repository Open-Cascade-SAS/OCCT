-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class ProductDefinition from StepBasic 

inherits TShared from MMgt

uses

	HAsciiString from TCollection, 
	ProductDefinitionFormation from StepBasic, 
	ProductDefinitionContext from StepBasic
is

	Create returns mutable ProductDefinition;
	---Purpose: Returns a ProductDefinition

	Init (me : mutable;
	      aId : mutable HAsciiString from TCollection;
	      aDescription : mutable HAsciiString from TCollection;
	      aFormation : mutable ProductDefinitionFormation from StepBasic;
	      aFrameOfReference : mutable ProductDefinitionContext from StepBasic) is virtual;

	-- Specific Methods for Field Data Access --

	SetId(me : mutable; aId : mutable HAsciiString);
	Id (me) returns mutable HAsciiString;
	SetDescription(me : mutable; aDescription : mutable HAsciiString);
	Description (me) returns mutable HAsciiString;
	SetFormation(me : mutable; aFormation : mutable ProductDefinitionFormation);
	Formation (me) returns mutable ProductDefinitionFormation;
	SetFrameOfReference(me : mutable; aFrameOfReference : mutable ProductDefinitionContext);
	FrameOfReference (me) returns mutable ProductDefinitionContext;

fields

	id : HAsciiString from TCollection;
	description : HAsciiString from TCollection;
	formation : ProductDefinitionFormation from StepBasic;
	frameOfReference : ProductDefinitionContext from StepBasic;

end ProductDefinition;
