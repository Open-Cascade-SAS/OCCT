-- Created on: 1995-03-06
-- Created by: Laurent PAINNOT
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Triangulation from DrawTrSurf inherits Drawable3D from Draw

	---Purpose: Used to display a triangulation.
	--          
	--          Display internal edges in blue
	--          Display boundary edges in red
	--          Optional display of triangles and nodes indices.

uses
    HArray1OfInteger from TColStd,
    Triangulation from Poly,
    Display       from Draw,
    Interpretor   from Draw,
    OStream

is

    Create(T : Triangulation from Poly)
    returns mutable Triangulation from DrawTrSurf;
    
    Triangulation(me)
    returns Triangulation from Poly;
    
    ShowNodes(me : mutable; B : Boolean);

    ShowNodes(me) returns Boolean;

    ShowTriangles(me : mutable; B : Boolean);

    ShowTriangles(me) returns Boolean;

    DrawOn(me; dis : in out Display);
    
    Copy(me) returns mutable Drawable3D from Draw
    is redefined;
	---Purpose: For variable copy.
	
    Dump(me; S : in out OStream)
    is redefined;
	---Purpose: For variable dump.

    Whatis(me; I : in out Interpretor from Draw)
    is redefined;
	---Purpose: For variable whatis command. Set  as a result  the
	--          type of the variable.

fields

    myTriangulation : Triangulation from Poly;
    myInternals     : HArray1OfInteger from TColStd;
    myFree          : HArray1OfInteger from TColStd;
    myNodes         : Boolean;
    myTriangles     : Boolean;

end Triangulation;
