-- Created on: 2001-04-24
-- Created by: Christian CAILLET
-- Copyright (c) 2001-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PlusMinusTolerance  from StepShape    inherits TShared

    ---Purpose : Added for Dimensional Tolerances

uses
    ToleranceMethodDefinition from StepShape,
    DimensionalCharacteristic from StepShape

is

    Create returns mutable PlusMinusTolerance;

    Init (me : mutable;
    	    range : ToleranceMethodDefinition from StepShape;
	    toleranced_dimension : DimensionalCharacteristic from StepShape);

    Range (me) returns ToleranceMethodDefinition from StepShape;
    SetRange (me : mutable; range : ToleranceMethodDefinition from StepShape);

    TolerancedDimension (me) returns DimensionalCharacteristic from StepShape;
    SetTolerancedDimension (me : mutable; toleranced_dimension : DimensionalCharacteristic from StepShape);

fields

    theRange : ToleranceMethodDefinition from StepShape;
    theTolerancedDimension : DimensionalCharacteristic from StepShape;

end PlusMinusTolerance;
