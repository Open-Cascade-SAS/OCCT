-- File:	Extrema_GenLocateExtCC.cdl
-- Created:	Tue Jul 18 17:43:18 1995
-- Author:	Modelistation
--		<model@metrox>
---Copyright:	 Matra Datavision 1995

generic class  GenLocateExtCC from Extrema 
(Curve1    as any;
 Tool1     as any;  -- as ToolCurve(Curve1);
 Curve2    as any;
 Tool2     as any;  -- as ToolCurve(Curve2);
 POnC      as any;
 Pnt       as any;
 Vec       as any)
					
    	---Purpose: It calculates the distance between two curves with
    	--          a close point; these distances can be maximum or 
    	--          minimum.


raises  DomainError  from Standard,
    	NotDone      from StdFail

private class CCLocF instantiates FuncExtCC (Curve1, Tool1,  
    	    	    	    	    	     Curve2, Tool2,  
    	    	    	    	    	     POnC, Pnt, Vec);

is
    Create (C1: Curve1; C2: Curve2; U0,V0: Real; TolU,TolV: Real)
    	returns GenLocateExtCC
    	---Purpose: Calculates the distance with a close point. The
    	--          close point is defined by a parameter value on each 
    	--          curve.
    	--          The function F(u,v)=distance(C1(u),C2(v)) has an 
    	--          extremun when gradient(f)=0. The algorithm searchs
    	--          the zero near the close point.
    	raises  DomainError;
    	    	-- if U0 and V0 are outside the definition ranges of the 
    	    	-- curves.
    
    IsDone (me) returns Boolean
    	---Purpose: Returns True if the distance is found.
    	is static;

    SquareDistance (me) returns Real
    	---Purpose: Returns the value of the extremum square distance.
	raises  NotDone from StdFail
	    	-- if IsDone(me)=False.
    	is static;

    Point (me; P1, P2: out POnC)
    	---Purpose: Returns the points of the extremum distance. 
    	--          P1 is on the first curve, P2 on the second one.
    	raises  NotDone from StdFail
    	    	-- if IsDone(me)=False.
    	is static;


fields
    myDone  : Boolean;
    mySqDist: Real;
    myPoint1: POnC;
    myPoint2: POnC;

end GenLocateExtCC;
