-- Created on: 1997-12-16
-- Created by: Denis PASCAL
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Expression from TDataStd inherits Attribute from TDF
    
    ---Purpose: Expression attribute. 
    --          ====================
    --
    --            * Data Structure  of the Expression   is stored in a
    --           string and references to variables used by the string
    --
    --  Warning:  To be consistent,  each  Variable  referenced by  the
    --          expression must have its equivalent in the string


uses Attribute         from TDF,
     Label             from TDF,
     GUID              from Standard,
     Real              from Standard,
     DataSet           from TDF,
     RelocationTable   from TDF,
     ExtendedString    from TCollection,
     AttributeList     from TDF
     

is

    ---Purpose: class methods
    --          =============

    GetID (myclass)    
    	---C++: return const & 
    returns GUID from Standard;
    

    Set (myclass ; label : Label from TDF)
    ---Purpose: Find, or create, an Expression attribute.
    returns Expression from TDataStd;
    
    ---Purpose: Expressionmethods
    --          ============

    Create
    returns mutable Expression from TDataStd;
    
    Name (me)
    ---Purpose: build and return the expression name
    returns ExtendedString from TCollection;
    
    SetExpression (me : mutable; E : ExtendedString from TCollection);
    
    GetExpression (me)
    returns ExtendedString from TCollection;    
    ---C++: return const &  

    GetVariables (me : mutable)
    ---C++: return &
    returns AttributeList from TDF;    

    ---Category: TDF_Attribute methods
    --           =====================
    
    ID (me) 
    ---C++: return const &  
    returns GUID from Standard;

    Restore (me: mutable; With : Attribute from TDF);

    NewEmpty(me)
    returns mutable Attribute from TDF;

    Paste (me; Into : mutable Attribute from TDF;
	       RT   : mutable RelocationTable from TDF);    

    Dump(me; anOS : in out OStream from Standard)
    returns OStream from Standard
    is redefined;
    ---C++: return &

fields

    myExpression : ExtendedString from TCollection;
    myVariables  : AttributeList from TDF;   
    
end Expression;
