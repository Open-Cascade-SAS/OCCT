-- Created on: 1993-06-02
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



deferred generic class SIFunction from IntStart 
    (ThePSurface as any)

inherits FunctionSetWithDerivatives from math 
    
	---Purpose: Template class for a function on a parametric surface.
	--          the form of the function is F(u,v) = 0 where u and v are
	--          the parameteric coordinates of a point on the surface.
       

uses Vector  from math,
     Matrix  from math,
     Pnt     from gp,
     Vec     from gp,
     Dir2d   from gp


raises UndefinedDerivative from StdFail

is

    Set(me: in out; PS: ThePSurface)
    
    	is static;


    NbVariables(me)

	---Purpose: This method has to return 2.
    	returns Integer from Standard;


    NbEquations(me)

	---Purpose: This method has to return 1.
    	returns Integer from Standard;


    Value(me : in out; X : Vector from math;
                       F : out Vector from math)

	---Purpose: The dimension of F is 1.

    	returns Boolean from Standard;


    Derivatives(me : in out; X : Vector from math;
                             D : out Matrix from math)

	---Purpose: The dimension of D is (1,2).

    	returns Boolean from Standard;


    Values(me : in out; X : Vector from math;
                        F : out Vector from math;
                        D : out Matrix from math)

    	returns Boolean from Standard;


    Root(me)

	---Purpose: Root is the value of the function at the solution.
	--          It is a vector of dimension 1, i-e a real.

    	returns Real from Standard
    	is static;


    Tolerance(me)
    
	---Purpose: Returns the value Tol so that if Abs(Func.Root())<Tol
	--          the function is considered null.
    
    	returns Real from Standard
	is static;


    Point(me)

	---Purpose: Returns the value of the solution point on the surface.

    	returns Pnt from gp
    	is static;
    

    IsTangent(me : in out)

    	returns Boolean from Standard 
    	is static;
    

    Direction3d(me: in out)

    	returns Vec from gp
    	raises UndefinedDerivative from StdFail
    	is static;
    

    Direction2d(me: in out)

    	returns Dir2d from gp
    	raises UndefinedDerivative from StdFail
    	is static;
    

end SIFunction;
