-- File:	MeshDS_Element2d.cdl
-- Created:	Tue Mar 16 15:28:35 1993
-- Author:	Didier PIFFAULT
--		<dpf@phylox>
---Copyright:	 Matra Datavision 1993


deferred generic class Element2d from MeshDS (dummyarg as any)

	---Purpose: Describes the necessary  services of an  Element2d
	--          for a mesh data structure.


uses    Integer from Standard,
    	Boolean from Standard,
	DegreeOfFreedom from MeshDS


is      Edges         (me; e1, e2, e3 : out Integer from Standard;
    	    	    	   o1, o2, o3 : out Boolean from Standard);
	   ---Purpose: Gives the   indices  of  the   edges    and the
	   --          orientation of each one.


    	Movability    (me)
	    	returns DegreeOfFreedom from MeshDS;
    	    ---Purpose: The movability of the triangle.


	SetMovability     (me      : in out;
    	    	    	   canMove : DegreeOfFreedom from MeshDS);


---Purpose: For maping the Elements.
--          Same Element -> Same HashCode
--          Different Elements -> Not IsEqual but can have same HashCode 

    	HashCode      (me;
    	    	       Upper : Integer from Standard)
	---C++: function call
    	        returns Integer from Standard;


    	IsEqual       (me; Other: Element2d from MeshDS)
	    ---C++: alias operator ==
    	    	returns Boolean from Standard;


end Element2d;
