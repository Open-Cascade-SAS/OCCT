-- Created on: 1992-03-25
-- Created by: Isabelle GRIGNON
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Couple from IntSurf

	---Purpose: creation d 'un couple de 2 entiers

is

     Create
     	returns Couple from IntSurf;
     	---C++: inline

     Create(Index1, Index2 : Integer from Standard)
    	---C++: inline
    	returns Couple from IntSurf;
	
     
     First(me) returns Integer from Standard
     ---Purpose: returns the first element 
     ---C++: inline
     is static;


     Second (me) returns Integer from Standard
     ---Purpose: returns the Second element 
     ---C++: inline
     is static;


fields

    firstInteger  : Integer from Standard;
    secondInteger : Integer from Standard;

end Couple;


