-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ProductDefinitionFormationWithSpecifiedSource from StepBasic 

inherits ProductDefinitionFormation from StepBasic 

uses

	Source from StepBasic, 
	HAsciiString from TCollection, 
	Product from StepBasic
is

	Create returns mutable ProductDefinitionFormationWithSpecifiedSource;
	---Purpose: Returns a ProductDefinitionFormationWithSpecifiedSource


	Init (me : mutable;
	      aId : mutable HAsciiString from TCollection;
	      aDescription : mutable HAsciiString from TCollection;
	      aOfProduct : mutable Product from StepBasic) is redefined;

	Init (me : mutable;
	      aId : mutable HAsciiString from TCollection;
	      aDescription : mutable HAsciiString from TCollection;
	      aOfProduct : mutable Product from StepBasic;
	      aMakeOrBuy : Source from StepBasic) is virtual;

	-- Specific Methods for Field Data Access --

	SetMakeOrBuy(me : mutable; aMakeOrBuy : Source);
	MakeOrBuy (me) returns Source;

fields

	makeOrBuy : Source from StepBasic; -- an Enumeration

end ProductDefinitionFormationWithSpecifiedSource;
