-- Created on: 1998-01-26
-- Created by: Sergey ZARITCHNY
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class EllipseRadiusPresentation from DsgPrs 

	---Purpose: 

uses
    Presentation from Prs3d,
    Pnt          from gp,
    Elips        from gp, 
    OffsetCurve  from Geom,
    Drawer       from Prs3d,
    ArrowSide    from DsgPrs,
    ExtendedString from TCollection

is
      Add( myclass; aPresentation   : Presentation   from Prs3d;
    	    	    aDrawer         : Drawer         from Prs3d; 
		    theval          : Real           from Standard;
		    aText           : ExtendedString from TCollection; 
                    AttachmentPoint : Pnt            from gp;
    	    	    anEndOfArrow    : Pnt            from gp; 
		    aCenter         : Pnt            from gp; 
		    IsMaxRadius     : Boolean        from  Standard;
		    ArrowSide: ArrowSide             from DsgPrs);
		   ---Purpose: draws a  Radius  (Major  or  Minor)   
    	    	   -- representation for whole ellipse  case
		   
    Add( myclass; aPresentation   : Presentation   from Prs3d;
    	    	  aDrawer         : Drawer         from Prs3d; 
		  theval          : Real           from Standard;
		  aText           : ExtendedString from TCollection; 
		  anEllipse       : Elips          from gp;  
                  AttachmentPoint : Pnt            from gp; 
		  anEndOfArrow    : Pnt            from gp; 
		  aCenter         : Pnt            from gp;
		  uFirst          : Real           from Standard;  
		  IsInDomain      : Boolean        from Standard; 
		  IsMaxRadius     : Boolean        from Standard;
	          ArrowSide       : ArrowSide      from DsgPrs);
		   ---Purpose: draws a  Radius  (Major  or  Minor) representation     
    	    	   --  for arc of an ellipse  case 

		   
    Add( myclass; aPresentation   : Presentation   from Prs3d;
    	    	  aDrawer         : Drawer         from Prs3d; 
		  theval          : Real           from Standard;
		  aText           : ExtendedString from TCollection; 
    	    	  aCurve          : OffsetCurve    from Geom;
                  AttachmentPoint : Pnt            from gp; 
		  anEndOfArrow    : Pnt            from gp; 
		  aCenter         : Pnt            from gp;
		  uFirst          : Real           from Standard;  
		  IsInDomain      : Boolean        from Standard; 
		  IsMaxRadius     : Boolean        from Standard;
	          ArrowSide       : ArrowSide      from DsgPrs);
		   ---Purpose: draws a  Radius  (Major  or  Minor) representation     
    	    	   --  for arc of an offset  curve  from  ellipse

end EllipseRadiusPresentation;
