-- Created on: 1994-12-21
-- Created by: Christian CAILLET
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class DispPerSignature  from IFSelect  inherits Dispatch

    ---Purpose : A DispPerSignature sorts input Entities according to a
    --           Signature : it works with a SignCounter to do this.

uses AsciiString from TCollection, Graph, SubPartsIterator, SignCounter

raises InterfaceError

is

    Create returns mutable DispPerSignature;
    ---Purpose : Creates a DispPerSignature with no SignCounter (by default,
    --           produces only one packet)

    SignCounter (me) returns mutable SignCounter;
    ---Purpose : Returns the SignCounter used for splitting

    SetSignCounter (me : mutable; sign : mutable SignCounter);
    ---Purpose : Sets a SignCounter for sort
    --           Remark : it is set to record lists of entities, not only counts

    SignName (me) returns CString;
    ---Purpose : Returns the name of the SignCounter, which caracterises the
    --           sorting criterium for this Dispatch

    Label (me) returns AsciiString from TCollection;
    ---Purpose : Returns as Label, "One File per Signature <name>"

    	--  --    Evaluation    --  --

    LimitedMax (me; nbent : Integer; max : out Integer) returns Boolean
    	is redefined;
    ---Purpose : Returns True, maximum count is given as <nbent>

--    PacketsCount (me; G : Graph; count : out Integer) returns Boolean
--    	is not redefined : Packets must be first determined before counting

    Packets (me; G : Graph; packs : in out SubPartsIterator)
    	raises InterfaceError;
    ---Purpose : Computes the list of produced Packets. It defines Packets from
    --           the SignCounter, which sirts the input Entities per Signature
    --           (specific of the SignCounter).

fields

    thesign : SignCounter;

end DispPerSignature;
