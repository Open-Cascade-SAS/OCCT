-- Created on: 1993-10-18
-- Created by: Christophe MARION
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class EdgeFaceTool from HLRBRep

	---Purpose: The EdgeFaceTool computes the  UV coordinates at a
	--          given parameter on a Curve and a Surface.  It also
	--          compute the signed  curvature value in a direction
	--          at a given u,v point on a surface.

uses
    Address  from Standard,
    Boolean  from Standard,
    Real     from Standard,
    Dir      from gp

is
    CurvatureValue(myclass;
                   F  : Address from Standard; -- as Surface from HLRBRep
                   U  : Real    from Standard;
                   V  : Real    from Standard;
                   Tg : Dir     from gp)       -- as tangent of the  edge
    returns Real from Standard;                -- at U,V point.
    
    UVPoint(myclass;
            Par :     Real    from Standard;
            E   :     Address from Standard; -- as Curve   from HLRBRep
            F   :     Address from Standard; -- as Surface from HLRBRep
	    U,V : out Real    from Standard)
    	---Purpose: return True if U and V are found.
    returns Boolean from Standard;
    
end EdgeFaceTool;
