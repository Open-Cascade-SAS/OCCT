-- Created on: 1998-06-03
-- Created by: data exchange team
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package ShapeFix 

  ---Purpose:  This package provides algorithms for fixing
  -- problematic (violating Open CASCADE requirements) shapes.
  -- Tools from package ShapeAnalysis are used for detecting the problems. The
  -- detecting and fixing is done taking in account various
  -- criteria implemented in BRepCheck package. 
  -- Each class of package ShapeFix deals with one
	-- certain type of shapes or with some family of problems.

uses

    gp,
    Geom,
    Geom2d,
    Geom2dAPI,
    GeomAbs,
    Adaptor3d,
    TCollection,
    TColStd,
    TopAbs,
    TopLoc,
    TopoDS, 
    TopTools,
    Message,
    ShapeExtend,
    ShapeAnalysis,
    ShapeConstruct,
    ShapeBuild,
    Bnd

is

    -- classes
    class Root;    

    class EdgeProjAux;

    class Edge;

    class Wire;

    class Face;

    class FixSmallFace;

    class FixSmallSolid;

    class WireVertex;

    class Wireframe;

    class FreeBounds;

    class FaceConnect;

    class Shell;

    class Solid;

    class ShapeTolerance;

    class Shape;

    class EdgeConnect;

    class ComposeShell;

    class SplitCommonVertex;

    class WireSegment;

    class IntersectionTool;

    class SplitTool;

    imported SequenceOfWireSegment;
    
    imported DataMapOfShapeBox2d;
    
    imported DataMapIteratorOfDataMapOfShapeBox2d;


    SameParameter (shape       : Shape from TopoDS;
                   enforce     : Boolean;
                   preci       : Real = 0.0;
                   theProgress : ProgressIndicator from Message = 0;
                   theMsgReg   : BasicMsgRegistrator from ShapeExtend = 0)
    returns Boolean;
    	---Purpose : Runs SameParameter from BRepLib with these adaptations :
    	--           <enforce> forces computations, else they are made only on
    	--             Edges with flag SameParameter false
    	--           <preci>, if not precised, is taken for each EDge as its own
    	--           Tolerance
    	--           Returns True when done, False if an exception has been raised
    	--           In case of exception anyway, as many edges as possible have
    	--           been processed. The passed progress indicator allows user
    	--           to consult the current progress stage and abort algorithm
    	--           if needed.

    EncodeRegularity (shape: Shape from TopoDS; tolang: Real = 1.0e-10);
    	---Purpose : Runs EncodeRegularity from BRepLib taking into account
      --           shared components of assemblies, so that each component
      --           is processed only once

    RemoveSmallEdges (shape: in out Shape from TopoDS; Tolerance: Real; context: in out ReShape from ShapeBuild) 
    	returns Shape from TopoDS;
      ---Purpose: Removes edges which are less than given tolerance from shape
      --          with help of ShapeFix_Wire::FixSmall()

    FixVertexPosition(theshape: in out Shape from TopoDS;
		      theTolerance: Real; 
    	    	      thecontext: ReShape from ShapeBuild) returns Boolean;
      ---Purpose: Fix position of the vertices having tolerance more tnan specified one.;       
    	 
    LeastEdgeSize(theshape: in out Shape from TopoDS) returns Real;
      ---Purpose: Calculate size of least edge;       
    	 

end ShapeFix;
