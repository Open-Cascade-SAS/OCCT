-- Created on: 2002-01-04
-- Created by: data exchange team
-- Copyright (c) 2002-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1

class Subedge from StepShape
inherits Edge from StepShape

    ---Purpose: Representation of STEP entity Subedge

uses
    HAsciiString from TCollection,
    Vertex from StepShape,
    Edge from StepShape

is
    Create returns Subedge from StepShape;
	---Purpose: Empty constructor

    Init (me: mutable; aRepresentationItem_Name: HAsciiString from TCollection;
                       aEdge_EdgeStart: Vertex from StepShape;
                       aEdge_EdgeEnd: Vertex from StepShape;
                       aParentEdge: Edge from StepShape);
	---Purpose: Initialize all fields (own and inherited)

    ParentEdge (me) returns Edge from StepShape;
	---Purpose: Returns field ParentEdge
    SetParentEdge (me: mutable; ParentEdge: Edge from StepShape);
	---Purpose: Set field ParentEdge

fields
    theParentEdge: Edge from StepShape;

end Subedge;
