-- Created on: 2004-07-14
-- Created by: Sergey KUUL
-- Copyright (c) 2004-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class SplitTool from ShapeFix

	---Purpose: Tool for splitting and cutting edges; includes methods
	--          used in OverlappingTool and IntersectionTool

uses

    Face from TopoDS,
    Edge from TopoDS,
    Vertex from TopoDS,
    ReShape from ShapeBuild,
    SequenceOfShape from TopTools

is
    Create returns SplitTool from ShapeFix;
    	---Purpose: Empty constructor
	
    SplitEdge(me; edge: Edge from TopoDS;
    	    	  param: Real from Standard;
    	          vert: Vertex from TopoDS;
    	    	  face: Face from TopoDS;
	          newE1: in out Edge from TopoDS;
    	    	  newE2: in out Edge from TopoDS;
    	          tol3d, tol2d : Real from Standard)
    returns Boolean from Standard;
    	---Purpose: Split edge on two new edges using new vertex "vert"
	--          and "param" - parameter for splitting
	--          The "face" is necessary for pcurves and using TransferParameterProj

    SplitEdge (me; edge: Edge from TopoDS;
    	       	   param1: Real from Standard;
    	       	   param2: Real from Standard;
    	       	   vert: Vertex from TopoDS;
	       	   face: Face from TopoDS;
	           newE1: in out Edge from TopoDS;
    	    	   newE2: in out Edge from TopoDS;
               	   tol3d, tol2d : Real from Standard)
    returns Boolean from Standard;
    	---Purpose: Split edge on two new edges using new vertex "vert"
	--          and "param1" and "param2" - parameter for splitting and cutting
	--          The "face" is necessary for pcurves and using TransferParameterProj

    CutEdge(me; edge: Edge from TopoDS; pend: Real from Standard;
    	        cut: Real from Standard; face: Face from TopoDS;
	        iscutline: in out Boolean from Standard)
    returns Boolean from Standard;
    	---Purpose: Cut edge by parameters pend and cut

    SplitEdge(me; edge: Edge from TopoDS; fp: Real from Standard;
    	          V1: Vertex from TopoDS; lp: Real from Standard;
    	          V2: Vertex from TopoDS; face: Face from TopoDS;
	          SeqE: in out SequenceOfShape from TopTools;
		  aNum: in out Integer from Standard;
		  context: ReShape from ShapeBuild;
   	          tol3d, tol2d : Real from Standard)
    returns Boolean from Standard;
    	---Purpose: Split edge on two new edges using two new vertex V1 and V2
	--          and two parameters for splitting - fp and lp correspondingly
	--          The "face" is necessary for pcurves and using TransferParameterProj
	--          aNum - number of edge in SeqE which corresponding to [fp,lp]



end SplitTool;
