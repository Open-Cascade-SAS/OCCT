-- File:        AutoDesignNominalDateAndTimeAssignment.cdl
-- Created:     Mon Dec  4 12:02:23 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWAutoDesignNominalDateAndTimeAssignment from RWStepAP214

	---Purpose : Read & Write Module for AutoDesignNominalDateAndTimeAssignment

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     AutoDesignNominalDateAndTimeAssignment from StepAP214,
     EntityIterator from Interface

is

	Create returns RWAutoDesignNominalDateAndTimeAssignment;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable AutoDesignNominalDateAndTimeAssignment from StepAP214);

	WriteStep (me; SW : in out StepWriter; ent : AutoDesignNominalDateAndTimeAssignment from StepAP214);

	Share(me; ent : AutoDesignNominalDateAndTimeAssignment from StepAP214; iter : in out EntityIterator);

end RWAutoDesignNominalDateAndTimeAssignment;
