-- Created on: 1992-09-01
-- Created by: Remi GILET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class MakeMirror

from gce

    ---Purpose: This class mplements elementary construction algorithms for a
    -- symmetrical transformation in 3D space about a point,
    -- axis or plane. The result is a gp_Trsf transformation.
    -- A MakeMirror object provides a framework for:
    -- -   defining the construction of the transformation,
    -- -   implementing the construction algorithm, and
    -- -   consulting the result.
 

uses Pnt  from gp,
     Ax1  from gp,
     Ax2  from gp,
     Dir  from gp,
     Pln  from gp,
     Lin  from gp,
     Trsf from gp,
     Real from Standard
     
is

Create(Point : Pnt from gp) returns MakeMirror;
    ---Puprose: Makes a symmetry transformation of center <Point>.

Create(Axis : Ax1 from gp) returns MakeMirror;
    ---Puprose: Makes a symmetry transformation of axis <Axis>.

Create(Line : Lin from gp) returns MakeMirror;
    ---Puprose: Makes a symmetry transformation of axis <Line>.

Create(Point : Pnt from gp;
       Direc : Dir from gp) returns MakeMirror;
    ---Purpose: Makes a symmetry transformation af axis defined by 
    --          <Point> and <Direc>.

Create(Plane : Pln from gp) returns MakeMirror;
    ---Purpose: Makes a symmetry transformation of plane <Plane>.

Create(Plane : Ax2 from gp) returns MakeMirror;
    ---Purpose: Makes a symmetry transformation of plane <Plane>.

Value(me) returns Trsf from gp
    is static;
    ---C++: return const&
    ---Purpose: Returns the constructed transformation.
    
Operator(me) returns Trsf from gp
    is static;
    ---C++: return const&
    ---C++: alias "Standard_EXPORT operator gp_Trsf() const;"

fields

    TheMirror : Trsf from gp;

end MakeMirror;

