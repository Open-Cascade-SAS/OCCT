-- Created on: 1992-09-28
-- Created by: Remi GILET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MakeArcOfCircle from GCE2d inherits Root from GCE2d
    	---Purpose: Implements construction algorithms for an arc of
    	-- circle in the plane. The result is a Geom2d_TrimmedCurve curve.
    	-- A MakeArcOfCircle object provides a framework for:
    	-- -   defining the construction of the arc of circle,
    	-- -   implementing the construction algorithm, and
    	-- -   consulting the results. In particular, the Value
    	--   function returns the constructed arc of circle.
        
uses Pnt2d        from gp,
     Circ2d       from gp,
     Vec2d       from gp,
     Real         from Standard,
     Boolean      from Standard,
     TrimmedCurve from Geom2d

raises NotDone from StdFail

is

Create(Circ           : Circ2d  from gp                      ;
       Alpha1, Alpha2 : Real    from Standard                ;
       Sense          : Boolean from Standard = Standard_True) 
    returns MakeArcOfCircle;
    	---Purpose: Makes an arc of circle (TrimmedCurve from Geom2d) from 
    	--          a circle between two parameters Alpha1 and Alpha2.
    	--          The two parameters are angles. The parameters are 
    	--          in radians.

Create(Circ  : Circ2d  from gp                      ;
       P     : Pnt2d   from gp                      ;
       Alpha : Real    from Standard                ;
       Sense : Boolean from Standard = Standard_True) 
    returns MakeArcOfCircle;
    	---Purpose: Makes an arc of circle (TrimmedCurve from Geom2d) from 
    	--          a circle between point <P> and the parameter
        --          Alpha. Alpha is given in radians.

Create(Circ  : Circ2d  from gp                      ;
       P1    : Pnt2d   from gp                      ;
       P2    : Pnt2d   from gp                      ;
       Sense : Boolean from Standard = Standard_True) 
    returns MakeArcOfCircle;
    	---Purpose: Makes an arc of circle (TrimmedCurve from Geom2d) from 
    	--          a circle between two points P1 and P2.

Create(P1    : Pnt2d   from gp       ;
       P2    : Pnt2d   from gp       ;
       P3    : Pnt2d   from gp       ) 
    returns MakeArcOfCircle;
    	---Purpose: Makes an arc of circle (TrimmedCurve from Geom2d) from 
    	--          three points P1,P2,P3 between two points P1 and P3,
    	--          and passing through the point P2.

Create(P1    : Pnt2d   from gp       ;
       V     : Vec2d   from gp       ;
       P2    : Pnt2d   from gp       )
    returns MakeArcOfCircle;
    	---Purpose: Makes an arc of circle (TrimmedCurve from Geom2d) from 
    	--          two points P1,P2 and the tangente to the solution at 
    	--          the point P1.

Value(me) returns TrimmedCurve from Geom2d
    raises NotDone
    is static;
    	---C++: return const&
    	---Purpose: Returns the constructed arc of circle.
    	-- Exceptions StdFail_NotDone if no arc of circle is constructed.

Operator(me) returns TrimmedCurve from Geom2d
    is static;
    	---C++: return const&
    	---C++: alias "Standard_EXPORT operator Handle_Geom2d_TrimmedCurve() const;"

fields

    TheArc : TrimmedCurve from Geom2d;
    --The solution from Geom2d.
    
end MakeArcOfCircle;
