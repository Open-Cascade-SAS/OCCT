-- Created on: 1995-03-15
-- Created by: Laurent PAINNOT
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PolygonOnTriangulation from BRep inherits CurveRepresentation from  BRep


    	---Purpose: A representation by an array of nodes on a 
    	--          triangulation.


uses Location               from TopLoc,
     PolygonOnTriangulation from Poly,
     Triangulation          from Poly


is

    Create(P: PolygonOnTriangulation from Poly;
    	   T: Triangulation          from Poly;
	   L: Location               from TopLoc)
    returns mutable PolygonOnTriangulation from BRep;


    IsPolygonOnTriangulation(me) returns Boolean
    	---Purpose: returns True.
    is redefined;

    IsPolygonOnTriangulation(me; T : Triangulation from Poly;
                            	 L : Location from TopLoc)    returns Boolean
	---Purpose: Is it a polygon in the definition of <T> with
	--          location <L>.
    is redefined;

    PolygonOnTriangulation(me: mutable; P: PolygonOnTriangulation from Poly)
    	---Purpose: returns True.
    is redefined;

    Triangulation(me) returns any Triangulation from Poly
    	---C++: return const&
    is redefined;
    
    PolygonOnTriangulation(me) returns any PolygonOnTriangulation from Poly
    	---C++: return const&
    is redefined;

    
    Copy(me) returns mutable CurveRepresentation from BRep is virtual;
	---Purpose: Return a copy of this representation.


fields

myPolygon       : PolygonOnTriangulation    from Poly;
myTriangulation : Triangulation             from Poly;

end PolygonOnTriangulation;
