-- Created on: 1999-02-26
-- Created by: Christian CAILLET
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class SelectPCurves  from IGESSelect    inherits SelectExplore

    ---Purpose : This Selection returns the pcurves which lie on a face
    --           In two modes : global (i.e. a CompositeCurve is not explored)
    --           or basic (all the basic curves are listed)

uses AsciiString from TCollection, Transient, EntityIterator, Graph

is

    Create (basic : Boolean) returns mutable SelectPCurves;
    ---Purpose : Creates a SelectPCurves
    --           basic True  : lists all the components of pcurves
    --           basic False : lists the uppest level definitions
    --             (i.e. stops at CompositeCurve)

    Explore (me; level : Integer; ent : Transient; G : Graph;
    	     explored : in out EntityIterator)
    	returns Boolean;
    ---Purpose : Explores an entity, to take its contained PCurves
    --           An independant curve is IGNORED : only faces are explored

    ExploreLabel (me) returns AsciiString from TCollection;
    ---Purpose : Returns a text defining the criterium : "Basic PCurves" or
    --           "Global PCurves"

fields

    thebasic : Boolean;

end SelectPCurves;
