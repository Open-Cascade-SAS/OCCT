-- Created on: 1993-07-06
-- Created by: Yves FRICAUD
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package MAT2d 

	---Purpose : Package of computation of Bisector locus on a
        --           Set of geometrys from Geom2d.

uses
    GeomAbs,
    MMgt,
    gp,
    Geom2d,
    TColStd,
    TCollection,
    TColgp,
    TColGeom2d,
    MAT,
    Bisector

is

    deferred class SketchExplorer;

    class Tool2d;

    class Mat2d;

    class Connexion;

    class MiniPath;

    class Circuit;

    class CutCurve;   

    imported SequenceOfConnexion; 

    imported DataMapOfIntegerSequenceOfConnexion;

    imported DataMapIteratorOfDataMapOfIntegerSequenceOfConnexion;
                                         
    imported Array2OfConnexion; 
               

    imported DataMapOfIntegerBisec;
               

    imported DataMapIteratorOfDataMapOfIntegerBisec; 
					    
    imported DataMapOfIntegerPnt2d;
					    
    imported DataMapIteratorOfDataMapOfIntegerPnt2d;  
	    
    imported DataMapOfIntegerVec2d;
	    
    imported DataMapIteratorOfDataMapOfIntegerVec2d; 

    imported SequenceOfSequenceOfCurve; 
					    
    imported SequenceOfSequenceOfGeometry; 

    imported DataMapOfIntegerConnexion;

    imported DataMapIteratorOfDataMapOfIntegerConnexion;

    class BiInt;
	
    class MapBiIntHasher;
    
    imported DataMapOfBiIntSequenceOfInteger;
    
    imported DataMapIteratorOfDataMapOfBiIntSequenceOfInteger;
        
    imported DataMapOfBiIntInteger;
        
    imported DataMapIteratorOfDataMapOfBiIntInteger;
end MAT2d;



