-- Created on: 1995-02-01
-- Created by: Marie Jose MARTZ
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Geom2dPoint from Geom2dToIGES inherits Geom2dEntity from Geom2dToIGES

    ---Purpose: This class implements the transfer of the Point Entity from Geom2d
    --          to IGES . These are :
    --          . 2dPoint
    --              * 2dCartesianPoint 

  
uses

    Point          from Geom2d,
    CartesianPoint from Geom2d,
    Point          from IGESGeom,
    Geom2dEntity   from Geom2dToIGES
     
is 
    
    Create returns Geom2dPoint from Geom2dToIGES;


    Create(G2dE : Geom2dEntity from Geom2dToIGES)  
    	 returns Geom2dPoint from Geom2dToIGES;
    ---Purpose : Creates a tool Geom2dPoint ready to run and sets its
    --         fields as G2dE's.

    Transfer2dPoint            (me    : in out;
                                start : Point from Geom2d)
    	 returns Point from IGESGeom;
    ---Purpose :  Transfert  a  Point from Geom to IGES. If this
    --            Entity could not be converted, this member returns a NullEntity.

    Transfer2dPoint            (me    : in out;
                                start : CartesianPoint from Geom2d)
    	 returns Point from IGESGeom;
    ---Purpose :  Transfert  a  CartesianPoint from Geom to IGES. If this
    --            Entity could not be converted, this member returns a NullEntity.


end Geom2dPoint;


