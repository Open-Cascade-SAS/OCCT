-- Created on: 1995-12-21
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class EdgeBuilder from TopOpeBRepBuild 
    inherits Area1dBuilder from TopOpeBRepBuild 

uses
    
    Shape from TopoDS,
    PaveSet from TopOpeBRepBuild,
    PaveClassifier from TopOpeBRepBuild,
    LoopSet from TopOpeBRepBuild,
    LoopClassifier from TopOpeBRepBuild
    
is

    Create returns EdgeBuilder;

    Create(LS : in out PaveSet; LC : in out PaveClassifier;
    	   ForceClass : Boolean = Standard_False) returns EdgeBuilder;
    ---Purpose: Creates a EdgeBuilder to find the areas of
    -- the shapes described by <LS> using the classifier <LC>.
    
    InitEdgeBuilder(me : in out;
    	    	    LS : in out LoopSet; LC : in out LoopClassifier;
    	    	    ForceClass : Boolean = Standard_False) is static;

    -- Output methods 
    InitEdge(me : in out) is static;
    MoreEdge(me) returns Boolean from Standard is static;
    NextEdge(me : in out) is static;
    
    -- Exploration of the vertex of current edge
    InitVertex(me : in out) is static;
    MoreVertex(me) returns Boolean from Standard is static;
    NextVertex(me : in out) is static;
    Vertex(me) returns Shape from TopoDS is static;
    ---C++: return const &
    Parameter(me) returns Real is static;
    
end EdgeBuilder from TopOpeBRepBuild;
