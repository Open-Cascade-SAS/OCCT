-- Created on: 1996-12-16
-- Created by: Christian CAILLET
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SelectReal  from StepData    inherits SelectMember

    ---Purpose : A SelectReal is a SelectMember specialised for a basic real
    --           type in a select which also accepts entities : this one has
    --           NO NAME
    --           For a named select, see SelectNamed

uses CString, Logical

is

    Create returns mutable SelectReal;

    Kind (me) returns Integer  is redefined;
    --  fixed kind : Real

    Real  (me) returns Real  is redefined;

    SetReal (me : mutable; val : Real)  is redefined;

fields

    theval  : Real;

end SelectReal;
