-- Created on: 1993-07-21
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class MakeShape from BRepBuilderAPI inherits Command from BRepBuilderAPI

	---Purpose: This    is  the  root     class for     all  shape
	--          constructions.  It stores the result.
	--          
	--          It  provides deferred methods to trace the history
	--          of sub-shapes.

uses
    Shape             from TopoDS,
    Face              from TopoDS,
    Edge              from TopoDS,
    Vertex            from TopoDS,
    ShapeModification from BRepBuilderAPI,
    ListOfShape       from TopTools
    
    
raises
    NotDone           from StdFail

is
    Delete(me:out) is redefined;
    ---C++: alias "Standard_EXPORT virtual ~BRepBuilderAPI_MakeShape(){Delete() ; }"
    
    Initialize;
    
    Build(me : in out)
	---Purpose: This is  called by  Shape().  It does  nothing but
	--          may be redefined.
	---Level: Public
    is virtual;
	
    Shape(me) returns Shape from TopoDS
    	---Purpose: Returns a shape built by the shape construction algorithm.
    	-- Raises exception StdFail_NotDone if the shape was not built.
	---C++: return const &
	---C++: alias "Standard_EXPORT operator TopoDS_Shape() const;"
	---Level: Public
	    raises
    	NotDone from StdFail
    is static;


    ------------------------------------------------------------------
    --- The following methods are not implemented at this level.
    --  An empty list is returned.
    --- They are optional and must be redefined. 
    ------------------------------------------------------------------

    Generated (me: in out; S : Shape from TopoDS)
    	---Purpose: Returns the  list   of shapes generated   from the
    	--          shape <S>. 
        ---C++: return const & 
        ---Level: Public
    returns ListOfShape from TopTools
    is virtual;
    

    Modified (me: in out; S : Shape from TopoDS)
    	---Purpose: Returns the list  of shapes modified from the shape
    	--          <S>. 
        ---C++: return const & 
        ---Level: Public
    returns ListOfShape from TopTools
    is virtual;


    IsDeleted (me: in out; S : Shape from TopoDS)
    returns Boolean
    is virtual;
    	---Purpose: Returns true if the shape S has been deleted.

    
fields
 
    myShape      : Shape       from TopoDS   is protected;
    myGenerated  : ListOfShape from TopTools is protected;
    
end MakeShape;
