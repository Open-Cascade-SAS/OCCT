-- File:	RWStepAP203_RWStartRequest.cdl
-- Created:	Fri Nov 26 16:26:40 1999 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0
-- Copyright:	Matra Datavision 1999

class RWStartRequest from RWStepAP203

    ---Purpose: Read & Write tool for StartRequest

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    StartRequest from StepAP203

is
    Create returns RWStartRequest from RWStepAP203;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : StartRequest from StepAP203);
	---Purpose: Reads StartRequest

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: StartRequest from StepAP203);
	---Purpose: Writes StartRequest

    Share (me; ent : StartRequest from StepAP203;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWStartRequest;
