-- Created on: 1999-01-05
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Explorer from TopOpeBRepDS

uses

    Shape from TopoDS,
    Edge from TopoDS,
    Face from TopoDS,
    Vertex from TopoDS,
    ShapeEnum from TopAbs,
    HDataStructure from TopOpeBRepDS

raises

    NoMoreObject from Standard,
    NoSuchObject from Standard

is

    Create returns Explorer;

    Create(HDS:HDataStructure;T:ShapeEnum = TopAbs_SHAPE;findkeep : Boolean = Standard_True) returns Explorer;
    
    Init(me:in out;HDS:HDataStructure;T:ShapeEnum = TopAbs_SHAPE;findkeep : Boolean = Standard_True);

    Type(me) returns ShapeEnum from TopAbs;

    More(me) returns Boolean;

    Next(me : in out) raises NoMoreObject; -- when More returned False

    Current(me) returns Shape raises NoSuchObject from Standard; -- when More returns False;
    ---C++: return const &

    Index(me) returns Integer raises NoSuchObject from Standard; -- when More returns False;

    Face(me) returns Face raises NoSuchObject from Standard; -- when More returns False;
    ---C++: return const &

    Edge(me) returns Edge raises NoSuchObject from Standard; -- when More returns False;
    ---C++: return const &

    Vertex(me) returns Vertex raises NoSuchObject from Standard; -- when More returns False;
    ---C++: return const &        


    Find(me:in out) is private;
    
fields

    myHDS : HDataStructure from TopOpeBRepDS;
    myT : ShapeEnum from TopAbs;
    myI,myN : Integer;
    myB : Boolean;
    myFK : Boolean;

end Explorer from TopOpeBRepDS;
