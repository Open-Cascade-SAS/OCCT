-- Created on: 1993-03-03
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class LoopClassifier from TopOpeBRepBuild 

---Purpose: classify loops in order to build Areas

uses

    ShapeEnum from TopAbs,
    State from TopAbs,
    Loop from TopOpeBRepBuild
    
is

    Delete(me:out) is virtual;
    ---C++: alias "Standard_EXPORT virtual ~TopOpeBRepBuild_LoopClassifier(){Delete() ; }"
    
    Compare(me : in out; L1,L2 : Loop from TopOpeBRepBuild) 
    returns State from TopAbs is deferred;
    ---Purpose: Returns the state of loop <L1> compared with loop <L2>.

end LoopClassifier from TopOpeBRepBuild;
