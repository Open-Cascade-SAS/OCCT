-- Created on: 2002-01-16
-- Created by: Michael PONIKAROV
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ExtStringArray from PDataStd inherits Attribute from PDF

	---Purpose: 

uses HExtendedString          from PCollection,
     HArray1OfExtendedString from PColStd
     
     
is

    Create returns mutable ExtStringArray from PDataStd;

    Init(me : mutable; lower, upper : Integer from Standard);

    SetValue(me: mutable; Index : Integer from Standard; Value : HExtendedString from PCollection);
    
    Value(me;  Index : Integer from Standard) returns HExtendedString from PCollection;
   
    Lower (me) returns Integer from Standard;      

    Upper (me) returns Integer from Standard;   
     
fields
    myValue     :  HArray1OfExtendedString from PColStd;
end ExtStringArray;
