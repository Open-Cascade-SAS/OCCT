-- Created on: 1992-08-26
-- Created by: Remi GILET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class MakeTranslation

from gce

    ---Purpose: This class implements elementary construction algorithms for a
    -- translation in 3D space. The result is a gp_Trsf transformation.
    -- A MakeTranslation object provides a framework for:
    -- -   defining the construction of the transformation,
    -- -   implementing the construction algorithm, and
    -- -   consulting the result.

uses Pnt  from gp,
     Trsf from gp,
     Vec  from gp,
     Real from Standard
     
is

Create(Vect : Vec from gp) returns MakeTranslation;
    --- Purpose: Constructs a translation along the vector " Vect"
    
Create(Point1 : Pnt from gp;
       Point2 : Pnt from gp) returns MakeTranslation;
    ---Purpose: Constructs a translation along the vector
    --   (Point1,Point2) defined from the point Point1 to the point Point2.
        
Value(me) returns Trsf from gp
    is static;
    ---C++: return const&
    ---Purpose:
    -- Returns the constructed transformation.

Operator(me) returns Trsf from gp
    is static;
    ---C++: return const&
    ---C++: alias "Standard_EXPORT operator gp_Trsf() const;"

fields

    TheTranslation : Trsf from gp;

end MakeTranslation;

