-- Created on: 2005-12-21
-- Created by: Sergey KHROMOV
-- Copyright (c) 2005-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class UFunction from BRepGProp inherits Function from math

    ---Purpose: This class represents the integrand function for 
    --          computation of an inner integral. The returned value 
    --          depends on the value type and the flag IsByPoint. 
    --  
    --          The type of returned value is the one of the following 
    --          values: 
    --            -  GProp_Mass - volume computation. 
    --            -  GProp_CenterMassX, GProp_CenterMassY, 
    --               GProp_CenterMassZ - X, Y and Z coordinates of center 
    --                                   of mass computation. 
    --            -  GProp_InertiaXX, GProp_InertiaYY, GProp_InertiaZZ, 
    --               GProp_InertiaXY, GProp_InertiaXZ, GProp_InertiaYZ 
    --                                 - moments of inertia computation. 
    --  
    --          If the flag IsByPoint is set to Standard_True, the value is 
    --          returned for the region of space that is delimited by a 
    --          surface and a point. Otherwise all computations are 
    --          performed for the region of space delimited by a surface 
    --          and a plane.
 
uses
    Pnt       from gp,
    XYZ       from gp,
    Address   from Standard,
    Boolean   from Standard,
    Real      from Standard,
    ValueType from GProp,
    Face      from BRepGProp

is

    Create(theSurface: Face from BRepGProp; 
           theVertex : Pnt     from gp; 
           IsByPoint : Boolean from Standard; 
           theCoeffs : Address from Standard) 
    ---Purpose: Constructor. Initializes the function with the face, the 
    --          location point, the flag IsByPoint and the coefficients 
    --          theCoeff that have different meaning depending on the value 
    --          of IsByPoint. 
    --          If IsByPoint is equal to Standard_True, the number of the 
    --          coefficients is equal to 3 and they represent X, Y and Z 
    --          coordinates (theCoeff[0], theCoeff[1] and theCoeff[2] 
    --          correspondingly) of the shift, if the inertia is computed 
    --          with respect to the point different then the location. 
    --          If IsByPoint is equal to Standard_False, the number of the 
    --          coefficients is 4 and they represent the combination of 
    --          plane parameters and shift values.
    returns UFunction from BRepGProp;  
 
    SetValueType(me: in out; theType: ValueType from GProp); 
    ---Purpose: Setting the type of the value to be returned. 
    ---C++: inline 
 
    SetVParam(me: in out; theVParam: Real from Standard);
    ---Purpose: Setting the V parameter that is constant during the 
    --          integral computation.
    ---C++: inline 
 
    Value(me: in out; X:     Real from Standard; 
                      F: out Real from Standard) 
    ---Purpose: Returns a value of the function.
    returns Boolean from Standard 
    is redefined; 
 
    -----------------------
    --  Private methods  --
    -----------------------

    VolumeValue(me: in out; X      :     Real from Standard; 
                            thePMP0: out XYZ  from gp; 
                            theS   : out Real from Standard; 
                            theD1  : out Real from Standard) 
    ---Purpose: Private method. Returns the value for volume computation. 
    --          Other returned values are: 
    --            -  thePMP0 - PSurf(X,Y) minus Location. 
    --            -  theS and theD1 coeffitients that are computed and used 
    --               for computation of center of mass and inertia values 
    --               by plane.
    returns Real from Standard
    is private;
 
    CenterMassValue(me: in out; X:     Real from Standard;
                                F: out Real from Standard)
    ---Purpose: Private method. Returns a value for the center of mass
    --          computation. If the value type other then GProp_CenterMassX,
    --          GProp_CenterMassY or GProp_CenterMassZ this method returns
    --          Standard_False. Returns Standard_True in case of successful
    --          computation of a value.
    returns Boolean from Standard
    is private;
 
    InertiaValue(me: in out; X:     Real from Standard;
                             F: out Real from Standard)
    ---Purpose: Private method. Computes the value of intertia. The type of
    --          a value returned is defined by the value type. If it is
    --          other then GProp_InertiaXX, GProp_InertiaYY,
    --          GProp_InertiaZZ, GProp_InertiaXY, GProp_InertiaXZ or
    --          GProp_InertiaYZ, the method returns Standard_False. Returns
    --          Standard_True in case of successful computation of a value
    returns Boolean from Standard
    is private;

fields

    mySurface  : Face      from BRepGProp;
    myVertex   : Pnt       from gp;
    myCoeffs   : Address   from Standard;
    myVParam   : Real      from Standard;
    myValueType: ValueType from GProp;
    myIsByPoint: Boolean   from Standard;

end UFunction;
