-- Created on: 1992-11-10
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PathPoint from IntSurf 

	---Purpose: 

uses Pnt           from gp,
     Vec           from gp,
     Dir2d         from gp,
     HSequenceOfXY from TColgp

raises UndefinedDerivative from StdFail,
       OutOfRange          from Standard

is

    Create
    
    	returns PathPoint from IntSurf;


    Create (P: Pnt from gp; U,V: Real from Standard)
    
    	returns PathPoint from IntSurf;


    SetValue (me: in out; P: Pnt from gp; U,V: Real from Standard)
    
    	is static;


    AddUV(me: in out; U,V : Real from Standard)
    
	---C++: inline

    	is static;
	

    SetDirections(me: in out; V: Vec from gp; D: Dir2d from gp)
    
	---C++: inline

    	is static;
	

    SetTangency(me: in out; Tang: Boolean from Standard)
    
	---C++: inline

    	is static;



    SetPassing(me: in out; Pass: Boolean from Standard)
    
	---C++: inline

    	is static;


    Value(me)
    
    	returns Pnt from gp
	---C++: return const &
	---C++: inline

	is static;


    Value2d(me; U,V: out Real from Standard)
    
	---C++: inline
    	is static;


    IsPassingPnt(me)
    
    	returns Boolean from Standard
	---C++: inline

	is static;


    IsTangent(me)
    
    	returns Boolean from Standard
	---C++: inline

	is static;


    Direction3d(me)
    
    	returns Vec from gp
	---C++: return const &
	---C++: inline

	raises UndefinedDerivative from StdFail
	is static;


    Direction2d(me)
    
    	returns Dir2d from gp
	---C++: return const &
	---C++: inline

	raises UndefinedDerivative from StdFail
	is static;


    Multiplicity(me)
    
    	returns Integer from Standard
	---C++: inline

	is static;


    Parameters(me; Index: Integer from Standard;
                   U,V: out Real from Standard)

	---C++: inline

    	raises OutOfRange from Standard
    	is static;


fields

    pt     : Pnt           from gp;
    ispass : Boolean       from Standard;
    istgt  : Boolean       from Standard;
    vectg  : Vec           from gp;
    dirtg  : Dir2d         from gp;
    sequv  : HSequenceOfXY from TColgp;

end PathPoint;
