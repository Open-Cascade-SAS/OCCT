-- File:	Law_Interpol.cdl
-- Created:	Fri Feb  3 12:59:33 1995
-- Author:	Laurent BOURESCHE
--		<lbo@phylox>
---Copyright:	 Matra Datavision 1995


class Interpol from Law inherits BSpFunc from Law

	---Purpose: Provides an evolution law that interpolates a set
	--          of parameter and value pairs (wi, radi)

uses
    Array1OfPnt2d from TColgp

is

    Create returns mutable Interpol from Law;
    	---Purpose: Constructs an empty interpolative evolution law.
    	-- The function Set is used to define the law.
    Set(me        : mutable; 
    	ParAndRad : Array1OfPnt2d from TColgp;
    	Periodic  : Boolean from Standard = Standard_False);
    	---Purpose:
    	--    Defines this evolution law by interpolating the set of 2D
    	-- points ParAndRad. The Y coordinate of a point of
    	-- ParAndRad is the value of the function at the parameter
    	-- point given by its X coordinate.
    	-- If Periodic is true, this function is assumed to be periodic.
    	-- Warning
    	-- -   The X coordinates of points in the table ParAndRad
    	--   must be given in ascendant order.
    	-- -   If Periodic is true, the first and last Y coordinates of
    	--   points in the table ParAndRad are assumed to be
    	--   equal. In addition, with the second syntax, Dd and Df
    	--   are also assumed to be equal. If this is not the case,
    	--   Set uses the first value(s) as last value(s).
         
    SetInRelative(me        : mutable; 
    	          ParAndRad : Array1OfPnt2d from TColgp;
    	          Ud,Uf     : Real from Standard;
    	    	  Periodic  : Boolean from Standard = Standard_False);

    Set(me        : mutable; 
    	ParAndRad : Array1OfPnt2d from TColgp;
    	Dd,Df     : Real from Standard;
    	Periodic  : Boolean from Standard = Standard_False);
    	---Purpose:
    	--    Defines this evolution law by interpolating the set of 2D
    	-- points ParAndRad. The Y coordinate of a point of
    	-- ParAndRad is the value of the function at the parameter
    	-- point given by its X coordinate.
    	-- If Periodic is true, this function is assumed to be periodic.
    	-- In the second syntax, Dd and Df define the values of
    	-- the first derivative of the function at its first and last points.
    	-- Warning
    	-- -   The X coordinates of points in the table ParAndRad
    	--   must be given in ascendant order.
    	-- -   If Periodic is true, the first and last Y coordinates of
    	--   points in the table ParAndRad are assumed to be
    	--   equal. In addition, with the second syntax, Dd and Df
    	--   are also assumed to be equal. If this is not the case,
    	--   Set uses the first value(s) as last value(s).
    SetInRelative(me        : mutable; 
    	          ParAndRad : Array1OfPnt2d from TColgp;
    	          Ud,Uf     : Real from Standard;
    	          Dd,Df     : Real from Standard;
                  Periodic  : Boolean from Standard = Standard_False);

end Interpol;
