-- Created on: 1994-06-01
-- Created by: Christian CAILLET
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SelectSingleViewFrom  from IGESSelect  inherits SelectDeduct

    ---Purpose : This selection gets the Single Views attached to its input
    --           IGES entities. Single Views themselves or Drawings as passed
    --           as such (Drawings, for their Annotations)


uses AsciiString from TCollection, EntityIterator, Graph

raises InterfaceError

is

    Create returns SelectSingleViewFrom;
    ---Purpose : Creates a SelectSingleViewFrom

    HasUniqueResult (me) returns Boolean  is redefined protected;
    ---Purpose : Returns True, because selection works with a ViewSorter which
    --           gives a unique result

    RootResult (me; G : Graph) returns EntityIterator  raises InterfaceError;
    ---Purpose : Selects the Single Views attached (in Directory Part) to
    --           input entities

    Label (me) returns AsciiString from TCollection;
    ---Purpose : Returns the label, with is "Single Views attached"

end SelectSingleViewFrom;
