-- File:        ToroidalSurface.cdl
-- Created:     Mon Dec  4 12:02:32 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWToroidalSurface from RWStepGeom

	---Purpose : Read & Write Module for ToroidalSurface
	--           Check added by CKY , 7-OCT-1996

uses Check from Interface, ShareTool from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     ToroidalSurface from StepGeom,
     EntityIterator from Interface

is

	Create returns RWToroidalSurface;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable ToroidalSurface from StepGeom);

	WriteStep (me; SW : in out StepWriter; ent : ToroidalSurface from StepGeom);

	Share(me; ent : ToroidalSurface from StepGeom; iter : in out EntityIterator);

	Check(me; ent : ToroidalSurface from StepGeom; shares : ShareTool; ach : in out Check);

end RWToroidalSurface;
