-- File:	BOP_AreaBuilder.cdl
-- Created:	Thu Dec 21 17:07:40 1995
-- Author:	Jean Yves LEBEY
--		<jyl@meteox>
---Copyright:	 Matra Datavision 1995

class AreaBuilder from BOP

    ---Purpose:  
     
    --  The Root class for the algorithms that are used  to   
     
    --      Reconstruct complex  topological  
    --  objects as  Faces or Solids.
    --      Loop is  the  composite topological object of
    --  the boundary. Wire for a Face. Shell for a Solid.
    --      LoopSet is a  tool describing the object  to
    --  build.  It gives an iteration  on Loops.  For each
    --  Loop it tells if it is on the boundary or if it is
    --  an interference.
    --      LoopClassifier  is an algorithm  used to test
    --  if a Loop is inside  another  Loop.
    --  The  result of the  reconstruction is an iteration
    --  on the reconstructed areas.  An  area is described
    --  by a set of Loops.
    --      A AreaBuilder is built with :
    --    - a LoopSet describing the object to reconstruct.
    --    - a LoopClassifier providing the classification algorithm.

uses

    State from TopAbs,

    Loop                     from BOP,
    ListOfLoop               from BOP,
    ListIteratorOfListOfLoop from BOP,
    ListOfListOfLoop         from BOP,
    LoopSet                  from BOP,
    LoopClassifier           from BOP,
    LoopEnum                 from BOP, 
    ListIteratorOfListOfListOfLoop from BOP
    
is

    Create  
    	returns AreaBuilder;
    	---Purpose:  
    	--- Empty  Constructor 
    	---
    Create(LS :out LoopSet from BOP;  
    	   LC :out LoopClassifier from BOP;
    	   ForceClass : Boolean = Standard_False)  
    	returns AreaBuilder;
    	---Purpose:  
    	--- Creates the objectr to build the areas on
    	--- the shapes described by <LS> using the classifier <LC>.
    	---
    Delete(me:out) is virtual;
    	---C++: alias "Standard_EXPORT virtual ~BOP_AreaBuilder(){Delete() ; }"
    	---Purpose:  
    	--- Destructor
    	---
    InitAreaBuilder(me :out;
    	    	    LS :out LoopSet from BOP;  
    	    	    LC :out LoopClassifier;
    	    	    ForceClass : Boolean from Standard = Standard_False) 
    	is virtual;
    	---Purpose:  
    	--- Sets a AreaBuilder to find the areas on
    	--- the shapes described by <LS> using the classifier <LC>.
    	---
    CompareLoopWithListOfLoop(me;
    	    	    	      LC  : out LoopClassifier from BOP;
    	    	    	      L   : Loop from BOP;
    	    	    	      LOL : ListOfLoop from BOP;
    	    	    	      aWhat  : LoopEnum from BOP) 
    	returns State from TopAbs  
    	is static protected;
    	---Purpose:  
    	--- Compare position of the Loop <L> with the Area <LOL>
    	--- using the Loop Classifier <LC>.
    	---       According to <aWhat>, Loops of <LOL> are selected or not
    	---       during <LOL> exploration. 
    	---
    	-- Result : TopAbs_OUT     if <LOL> is empty
    	---      TopAbs_UNKNOWN if position undefined
    	---      TopAbs_IN      if <L> is inside all the selected Loops of <LOL>
    	---      TopAbs_OUT     if <L> is outside one of the selected Loops of <LOL>
    	---      TopAbs_ON      if <L> is on one of the selected Loops of <LOL>	
    	---
    	---

    --- Iteration on Areas   
    --
    InitArea(me:out)  
    	returns Integer from Standard is static;
    	---Purpose:  
    	--- Initialize iteration on areas.
    	---
    MoreArea(me)  
    	returns Boolean from Standard is static;
     
    NextArea(me:out)  
    	is static;

    -- 
    --  Iteration on Loops inside the Area   
    --
    InitLoop(me:out)  
    	returns Integer from Standard is static;
    	---Purpose:  
    	--- Initialize iteration on loops of current Area. 
    	---
    MoreLoop(me)  
    	returns Boolean from Standard is static;
     
    NextLoop(me:out)  
    	is static;
     
    Loop(me)  
    	returns Loop from BOP is static; 
    	---C++: return const&
    	---Purpose:  
    	--- Returns the current Loop in the current area.
    	---
    ---
    --- 
    ---  Methods that are not for public usage 
    ---	     
    ADD_Loop_TO_LISTOFLoop  (me;  
    	    	    	     L  : Loop from BOP;
    	    	    	     LOL: out ListOfLoop from BOP)  
    	is virtual;
    	---Purpose: 
    	--- Internal 
    	---
    REM_Loop_FROM_LISTOFLoop(me;  
    	    	    	     ITLOL: out ListIteratorOfListOfLoop from BOP; 
     	    	    	     LOL  : out ListOfLoop from BOP)
	 is virtual;
    	---Purpose: 
    	--- Internal 
    	---
    ADD_LISTOFLoop_TO_LISTOFLoop(me;  
    	    	    	    	 LOL1 : out ListOfLoop from BOP;
    	    	    	         LOL2 : out ListOfLoop from BOP)
    	is virtual;
    	---Purpose: 
    	--- Internal 
    	---
    Atomize(me; 
    	    state : in out State from TopAbs;  
    	    newstate : State from TopAbs)
    	is static protected;
    	---Purpose: 
    	--- Internal 
    	---
fields

    myArea         : ListOfListOfLoop               from BOP is protected;
    myAreaIterator : ListIteratorOfListOfListOfLoop from BOP is protected;
    myLoopIterator : ListIteratorOfListOfLoop       from BOP is protected;
    myUNKNOWNRaise : Boolean  from Standard is protected;
    
end AreaBuilder;

