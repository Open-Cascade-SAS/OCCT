-- Created on: 1995-09-18
-- Created by: Bruno DUMORTIER
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class MakeEvolved from BRepOffsetAPI inherits MakeShape from BRepBuilderAPI

	---Purpose: Describes functions to build evolved shapes.
    	-- An evolved shape is built from a planar spine (face or
    	-- wire) and a profile (wire). The evolved shape is the
    	-- unlooped sweep (pipe) of the profile along the spine.
    	-- Self-intersections are removed.
    	-- A MakeEvolved object provides a framework for:
    	-- - defining the construction of an evolved shape,
    	-- - implementing the construction algorithm, and
    	-- - consulting the result.
    	--        Computes an Evolved by 
	--             1 - sweeping a profil along a spine.
	--             2 - removing the self-intersections.
	--             
	--  The profile is defined in a Referential R. The position of
	--  the profile at the current point of the  spine is given by
	--  confusing R  and the local  referential given by (  D0, D1
	--  and the normal of the Spine)
	--  
	--  If the Boolean <AxeProf> is  true, R is  O,X,Y,Z 
	--  else R is defined as the local refential at the nearest 
	--  point of the profil to the spine.
	--  
	--   if <Solid> is TRUE the Shape result  is completed to be a
	--   solid or a compound of solids.



uses
    Evolved     from BRepFill,
    ListOfShape from TopTools,
    Shape       from TopoDS,	
    Face        from TopoDS,
    Wire        from TopoDS,
    JoinType    from GeomAbs
    
is
    Create returns MakeEvolved from BRepOffsetAPI;
    
    Create( Spine      : Wire      from TopoDS;
    	    Profil     : Wire      from TopoDS;
    	    Join       : JoinType  from GeomAbs  = GeomAbs_Arc;
	    AxeProf    : Boolean   from Standard = Standard_True;
    	    Solid      : Boolean   from Standard = Standard_False;
    	    ProfOnSpine: Boolean   from Standard = Standard_False;
    	    Tol        : Real      from Standard = 0.0000001)
	---Purpose: 
	---Level: Public 
    returns MakeEvolved from BRepOffsetAPI;

    Create( Spine      : Face      from TopoDS;
    	    Profil     : Wire      from TopoDS;
    	    Join       : JoinType  from GeomAbs  = GeomAbs_Arc;
	    AxeProf    : Boolean   from Standard = Standard_True;
    	    Solid      : Boolean   from Standard = Standard_False;
    	    ProfOnSpine: Boolean   from Standard = Standard_False;
    	    Tol        : Real      from Standard = 0.0000001)
	---Purpose: These constructors construct an evolved shape by sweeping the profile
    	-- Profile along the spine Spine.
    	--	The profile is defined in a coordinate system R.
    	-- The coordinate system is determined by AxeProf:
    	-- - if AxeProf is true, R is the global coordinate system,
    	-- - if AxeProf is false, R is computed so that:
    	--   - its origin is given by the point on the spine which is
    	--    closest to the profile,
    	--   - its "X Axis" is given by the tangent to the spine at this point, and
    	-- - its "Z Axis" is the normal to the plane which contains the spine.
    	--        The position of the profile at the current point of the
    	-- spine is given by making R coincident with the local
    	-- coordinate system given by the current point, the
    	-- tangent vector and the normal to the spine.
    	-- Join defines the type of pipe generated by the salient
    	-- vertices of the spine. The default type is GeomAbs_Arc
    	-- where the vertices generate revolved pipes about the
    	-- axis passing along the vertex and the normal to the
    	-- plane of the spine. At present, this is the only
    	-- construction type implemented.
    returns MakeEvolved from BRepOffsetAPI;

    Evolved(me) returns Evolved from BRepFill
	---C++: return const &
	---Level: Advanced
    is static;

    Build(me : in out)
    is redefined;
	---Purpose: Builds the resulting shape (redefined from MakeShape).
	---Level: Public    

    GeneratedShapes (me ;
    	    	     SpineShape : Shape from TopoDS;
    	    	     ProfShape  : Shape from TopoDS)
        ---Purpose: Returns   the  shapes  created  from   a  subshape
        --          <SpineShape>  of     the  spine   and   a subshape
        --          <ProfShape> on the profile.
        ---C++ : return const &          
    returns ListOfShape from TopTools
    is static;			 

    Top (me) returns Shape from TopoDS
       ---Purpose: Return the face Top if <Solid> is True in the constructor.
       ---C++ : return const &
    is static;

    Bottom (me) returns Shape from TopoDS
       ---Purpose: Return the face Bottom  if <Solid> is True in the constructor.
       ---C++ : return const &
    is static;
    
fields
    myEvolved : Evolved from BRepFill;
    
end MakeEvolved;
