-- Created on: 2001-12-19
-- Created by: Sergey KUUL
-- Copyright (c) 2001-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class MTHasher from MoniTool

	---Purpose: 
	-- The auxiliary class provides hash code for mapping objects   

is

    HashCode(myclass; Str : CString; Upper : Integer) returns Integer;
	---C++: inline
	---Purpose: Returns a HasCode value for the CString <Str>  in the
	-- range 0..Upper.
	-- Default ::HashCode(Str,Upper)
	
    IsEqual(myclass; Str1, Str2 : CString) returns Boolean;
	---C++: inline
	---Purpose: Returns True  when the two CString are the same. Two
	-- same strings must have the same hashcode, the
	-- contrary is not necessary.
	-- Default Str1 == Str2
	
end MTHasher;
