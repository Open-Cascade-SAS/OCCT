-- Created on: 1995-01-26
-- Created by: Mister rmi
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class SensitivePoint from Select2D inherits SensitiveEntity from Select2D

	---Purpose: A framework to define sensitive 2D points.

uses
    Integer from Standard,
    Pnt2d from gp,
    EntityOwner from SelectBasics,
    ListOfBox2d from SelectBasics  

is


    Create (OwnerId         : EntityOwner from SelectBasics;
    	    Location        : Pnt2d from gp;
    	    InitSensitivity : Real = 0)
    returns mutable SensitivePoint from Select2D;
    	---Purpose: Constructs the sensitive point object defined by the
    	-- owner OwnerId, the point Location and the sensitivity InitSensitivity.
    	-- InitSensitivity allows choice of dimensions in the
    	-- selectable box around the sensitive point. It is
    	-- initialized with a null value, and is given a working one by Set.
    
    
    Set(me:mutable; aSensitivity:Real) is static;
    	---Purpose: Sets the sensitivity aSensitivity for sensitive
    	-- primitives to find owners of points.

    Areas  (me:mutable ; aresul : in out ListOfBox2d from SelectBasics) is static;
    	---Level: Public 
    	---Purpose: Returns the 2Dbox around the point (this box) has to be enlarged (sensitivity = 0) 
    
    
    Location(me) returns Pnt2d from gp;
    	---Level: Public 
    	---C++: inline
    	---C++: return const&
    	---Purpose: returns the original point.
    
    
    
    Matches (me     : mutable ; 
    	     X,Y    : Real from Standard;
             aTol   : Real from Standard;
    	     DMin   : out Real from Standard) 
    returns Boolean
    is static;
    	---Purpose: if distance between P

    Matches (me  :mutable; 
             XMin,YMin,XMax,YMax : Real from Standard;
             aTol: Real from Standard) 
    returns Boolean
    is static;


fields
    
    mylocation    : Pnt2d from gp;
    mysensitivity : Real;

end SensitivePoint;

