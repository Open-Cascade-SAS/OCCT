-- Created on: 1999-02-12
-- Created by: Andrey BETENEV
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class TranslateCompositeCurve from StepToTopoDS 
    inherits Root from StepToTopoDS
	---Purpose: Translate STEP entity composite_curve to TopoDS_Wire
	--          If surface is given, the curve is assumed to lie on that
        --          surface and in case if any segment of it is a
	--          curve_on_surface, the pcurve for that segment will be taken.
	--          Note: a segment of composite_curve may be itself 
        --                composite_curve. Only one-level protection against 
        --                cyclic references is implemented.

uses
    TransientProcess from Transfer,
    CompositeCurve   from StepGeom,
    Surface          from StepGeom,
    Surface          from Geom,
    Wire             from TopoDS
    
is

    Create returns TranslateCompositeCurve;
        ---Purpose: Empty constructor
	
    Create (CC: CompositeCurve from StepGeom;
    	    TP: TransientProcess from Transfer)
    	returns TranslateCompositeCurve;
        ---Purpose: Translates standalone composite_curve

    Create (CC: CompositeCurve from StepGeom;
    	    TP: TransientProcess from Transfer;
    	    S : Surface from StepGeom;
    	    Surf: Surface from Geom)
    	returns TranslateCompositeCurve;
        ---Purpose: Translates composite_curve lying on surface 
	
    Init (me: in out;
          CC: CompositeCurve from StepGeom;
    	  TP: TransientProcess from Transfer)
    	returns Boolean;
        ---Purpose: Translates standalone composite_curve

    Init (me: in out;
          CC: CompositeCurve from StepGeom;
    	  TP: TransientProcess from Transfer;
    	  S : Surface from StepGeom;
    	  Surf: Surface from Geom)
    	returns Boolean;
        ---Purpose: Translates composite_curve lying on surface 

    Value (me) returns Wire from TopoDS;
        ---Purpose: Returns result of last translation or null wire if failed.
	---C++: return const &

    IsInfiniteSegment (me) returns Boolean;
        ---Purpose: Returns True if composite_curve contains a segment with infinite parameters.
        ---C++: inline 

fields

    myWire: Wire from TopoDS;
    myInfiniteSegment: Boolean;

end TranslateCompositeCurve;
