-- Created on: 1996-01-10
-- Created by: Denis PASCAL
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PlanarDistance from DrawDim inherits PlanarDimension from DrawDim

	---Purpose: PlanarDistance point/point
	--          PlanarDistance point/line
	--          PlanarDistance line/line

uses Face    from TopoDS,
     Pnt     from gp,
     Shape   from TopoDS,
     Edge    from TopoDS,
     Color   from Draw,
     Display from Draw

is

    Create (plane  : Face from TopoDS;
            point1 : Shape from TopoDS;
            point2 : Shape from TopoDS)
    returns PlanarDistance from DrawDim;
    
    Create (geom1 : Shape from TopoDS;
            geom2 : Shape from TopoDS)
    returns PlanarDistance from DrawDim; 
    
    DrawOn(me; dis : in out Display);

    ---Purpose: private
    Draw (me; p : Pnt from gp;
              e : Edge from TopoDS;
              d : in out Display) is private;
    
fields

    myGeom1 : Shape from TopoDS;
    myGeom2 : Shape from TopoDS;
    
end PlanarDistance;
