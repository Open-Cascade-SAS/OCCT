-- Created on: 2003-02-10
-- Created by: Sergey KUUL
-- Copyright (c) 2003-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class ConversionBasedUnitAndMassUnit from StepBasic inherits ConversionBasedUnit from StepBasic 

	--- This classe is an implementation of EXPRESS
	--  ANDOR Subtype Declaration.
uses

    MassUnit from StepBasic, 
    DimensionalExponents from StepBasic, 
    HAsciiString from TCollection, 
    MeasureWithUnit from StepBasic
    
is

    Create returns mutable ConversionBasedUnitAndMassUnit;
	---Purpose: Returns a ConversionBasedUnitAndLengthUnit

    Init (me: mutable; aDimensions: mutable DimensionalExponents from StepBasic)
    is redefined;

    Init (me: mutable; aDimensions: mutable DimensionalExponents from StepBasic;
	               aName      : mutable HAsciiString from TCollection;
	               aConversionFactor: mutable MeasureWithUnit from StepBasic) is redefined;

    -- Specific Methods for Field Data Access --

    SetMassUnit(me: mutable; aMassUnit: mutable MassUnit);
    
    MassUnit (me) returns mutable MassUnit;

    -- Specific Methods for ANDOR Field Data Access --

fields

    massUnit: MassUnit from StepBasic;

end ConversionBasedUnitAndMassUnit;
