-- Created on: 2003-04-29
-- Created by: Michael KLOKOV
-- Copyright (c) 2003-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class SectionHistoryCollector from BOP inherits HistoryCollector from BOP

uses
    Shape from TopoDS,
    Operation from BOP,
    PDSFiller from BOPTools,
    ListOfShape from TopTools,
    IndexedMapOfShape from TopTools, 
    IndexedDataMapOfShapeListOfShape from TopTools

is
    Create(theShape1   : Shape from TopoDS;
    	   theShape2   : Shape from TopoDS)
    	returns SectionHistoryCollector from BOP;

    SetResult(me: mutable; theResult: Shape from TopoDS;
    	    	    	   theDSFiller: PDSFiller from BOPTools)
    	is redefined virtual;


    -- private
    FillFaceSection(me: mutable; theDSFiller : PDSFiller from BOPTools;
    	    	    	    	 theResultMap: IndexedMapOfShape from TopTools) 
    is private;
    
    FillEdgeSection(me: mutable; theEdge     : Shape                            from TopoDS; 
    	    	    	    	 theDSFiller : PDSFiller                        from BOPTools; 
    	    	    	    	 theResultMap: IndexedMapOfShape                from TopTools; 
    	    	    	    	 theVEMapRes : IndexedDataMapOfShapeListOfShape from TopTools; 
    	    	    	    	 theEFMap    : IndexedDataMapOfShapeListOfShape from TopTools) 
    is private;

end SectionHistoryCollector from BOP;
