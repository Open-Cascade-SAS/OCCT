-- File:	StepData_SelectMember.cdl
-- Created:	Mon Dec 16 16:01:41 1996
-- Author:	Christian CAILLET
--		<cky@heliox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1996


class SelectMember  from StepData    inherits TShared

    ---Purpose : The general form for a Select Member. A Select Member can,
    --           either define a value of a basic type (such as an integer)
    --           with an additional information : a name or list of names
    --           which precise the meaning of this value
    --           or be an alternate value in a select, which also accepts an
    --           entity (in this case, the name is not mandatory)
    --           
    --           Several sub-types of SelectMember are defined for integer and
    --           real value, plus an "universal" one for any, and one more to
    --           describe a select with several names
    --           
    --           It is also possible to define a specific subtype by redefining
    --           virtual method, then give a better control
    --           
    --           Remark : this class itself could be deferred, because at least
    --           one of its virtual methods must be redefined to be usable

uses CString, ParamType from Interface, Logical from StepData

is

    Create returns mutable SelectMember;
    --  this constructor is useless, the class is empty

    HasName (me) returns Boolean  is virtual;
    ---Purpose : Tells if a SelectMember has a name. Default is False

    Name (me) returns CString  is virtual;
    ---Purpose : Returns the name of a SelectMember. Default is empty

    SetName (me : mutable; name : CString)  returns Boolean  is virtual;
    ---Purpose : Sets the name of a SelectMember, returns True if done, False
    --           if no name is allowed
    --           Default does nothing and returns False

    Matches (me; name : CString) returns Boolean  is virtual;
    ---Purpose : Tells if the name of a SelectMember matches a given one
    --           By default, compares the strings, can be redefined (optimised)

    Kind (me) returns Integer  is virtual;
    --  see Field for Kind (same codes)

    SetKind  (me : mutable; kind : Integer)  is virtual;
    --  called by various Set*

    ParamType (me) returns ParamType from Interface;
    ---Purpose : Returns the Kind of the SelectMember, under the form of an
    --           enum ParamType

    Int (me) returns Integer  is virtual;
    ---Purpose : This internal method gives access to a value implemented by an
    --           Integer (to read it)

    SetInt (me : mutable; val : Integer)  is virtual;
    ---Purpose : This internal method gives access to a value implemented by an
    --           Integer (to set it)

    Integer (me) returns Integer;
    ---Purpose : Gets the value as an Integer

    SetInteger (me : mutable; val : Integer);

    Boolean (me) returns Boolean;

    SetBoolean (me : mutable; val : Boolean);

    Logical (me) returns Logical;

    SetLogical (me : mutable; val : Logical);

    Real (me) returns Real  is virtual;

    SetReal (me : mutable; val : Real)  is virtual;

    String (me) returns CString  is virtual;

    SetString (me : mutable; val : CString)  is virtual;

    Enum (me) returns Integer;
    EnumText (me) returns CString  is virtual;
    --  By default, returns the String
    --  Can be redefined to return a String for instance bound with int value

    SetEnum (me : mutable; val : Integer; text : CString = "");
    --  calls SetInt (for val) and SetEnumText (see below)

    SetEnumText (me : mutable; val : Integer; text : CString)  is virtual;
    --  By default, calls SetString and disregards val
    --  It is enough for standard subtypes
    --  Can be redefined for a check on text and/or control of val and/or set
    --  val according to text

end SelectMember;
