-- Created on: 1991-05-13
-- Created by: Laurent PAINNOT
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class FunctionRoots from math
    ---Purpose:
    -- This class implements an algorithm which finds all the real roots of
    -- a function with derivative within a given range.
    -- Knowledge of the derivative is required.

uses FunctionWithDerivative from math,
     SequenceOfReal         from TColStd,
     SequenceOfInteger      from TColStd,
     OStream                from Standard

raises RangeError from Standard,
       NotDone from StdFail

is

    Create(F: in out FunctionWithDerivative; A, B: Real;
    	   NbSample: Integer; EpsX, EpsF, EpsNull, K : Real= 0.0) 

    ---Purpose: Calculates all the real roots of a function F-K within the range 
    -- A..B. whithout conditions on A and B
    -- A solution X is found when
    --   abs(Xi - Xi-1) <= Epsx and abs(F(Xi)-K) <= EpsF.
    -- The function is considered as null between A and B if
    -- abs(F-K) <= EpsNull within this range.
    
    returns FunctionRoots;
    
    IsDone(me)
    	---Purpose: Returns true if the computations are successful, otherwise returns false.
    	---C++: inline
    returns Boolean
    is static;


    IsAllNull(me)
    	---Purpose:
        -- returns true if the function is considered as null between A and B.
    	-- Exceptions
    	-- StdFail_NotDone if the algorithm fails (and IsDone returns false).	
    	---C++: inline
    returns Boolean
    raises NotDone
    is static;
    
    
    NbSolutions(me)
    	---Purpose: Returns the number of solutions found.
    	-- Exceptions
    	-- StdFail_NotDone if the algorithm fails (and IsDone returns false).
    	---C++: inline
    returns Integer
    raises NotDone
    is static;


    Value(me; Nieme: in Integer)
    	---Purpose: Returns the Nth value of the root of function F.
    	-- Exceptions
    	-- StdFail_NotDone if the algorithm fails (and IsDone returns false).
    	---C++: inline

    returns Real
    raises NotDone, RangeError
    is static;
    
    
    StateNumber(me; Nieme: in Integer)
    	---Purpose:
        -- returns the StateNumber  of the Nieme root.
        -- Exception RangeError is raised if Nieme is < 1
        --  or Nieme > NbSolutions.
    	---C++: inline

    returns Integer
    raises NotDone
    is static;

    
    Dump(me; o: in out OStream)
	---Purpose: Prints on the stream o information on the current state 
    	--          of the object.

    is static;


fields

Done:       Boolean;
AllNull:    Boolean;
Sol:        SequenceOfReal    from TColStd;
NbStateSol: SequenceOfInteger from TColStd;

end FunctionRoots;
