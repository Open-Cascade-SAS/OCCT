-- Created on: 1996-11-25
-- Created by: Philippe MANGIN
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class AppFunc from BRepBlend inherits AppFuncRoot from BRepBlend

	---Purpose: Function to approximate by AppSurface
	---Level: Advanced

uses
 Line        from BRepBlend,
 Point       from Blend,
 AppFunction from Blend,
 Function    from Blend,
 Vector      from math
 
raises OutOfRange

is
   Create(Line : in out Line from BRepBlend;
    	  Func : in out Function from Blend;
          Tol3d: Real;
          Tol2d: Real)
   ---Warning: The Object Func cannot be killed before me. 
   returns AppFunc; 

   Point(me;
    	 Func  : AppFunction from Blend; 
	 Param : Real;
	 Sol   : Vector from math;
	 Pnt   : in out Point from Blend);
	
   Vec(me;
       Sol : in out Vector from math;
       Pnt : Point from Blend);
	
end AppFunc;
