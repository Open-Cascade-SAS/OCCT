-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class CartesianTransformationOperator3d from StepGeom 

inherits CartesianTransformationOperator from StepGeom 

uses

	Direction from StepGeom, 
	Boolean from Standard, 
	HAsciiString from TCollection, 
	CartesianPoint from StepGeom, 
	Real from Standard
is

	Create returns CartesianTransformationOperator3d;
	---Purpose: Returns a CartesianTransformationOperator3d


	Init (me : mutable;
	      aName : HAsciiString from TCollection;
	      hasAaxis1 : Boolean from Standard;
	      aAxis1 : Direction from StepGeom;
	      hasAaxis2 : Boolean from Standard;
	      aAxis2 : Direction from StepGeom;
	      aLocalOrigin : CartesianPoint from StepGeom;
	      hasAscale : Boolean from Standard;
	      aScale : Real from Standard) is redefined;

	Init (me : mutable;
	      aName : HAsciiString from TCollection;
	      hasAaxis1 : Boolean from Standard;
	      aAxis1 : Direction from StepGeom;
	      hasAaxis2 : Boolean from Standard;
	      aAxis2 : Direction from StepGeom;
	      aLocalOrigin : CartesianPoint from StepGeom;
	      hasAscale : Boolean from Standard;
	      aScale : Real from Standard;
	      hasAaxis3 : Boolean from Standard;
	      aAxis3 : Direction from StepGeom) is virtual;

	-- Specific Methods for Field Data Access --

	SetAxis3(me : mutable; aAxis3 : Direction);
	UnSetAxis3 (me:mutable);
	Axis3 (me) returns Direction;
	HasAxis3 (me) returns Boolean;

fields

	axis3 : Direction from StepGeom;   -- OPTIONAL can be NULL
	hasAxis3 : Boolean from Standard;

end CartesianTransformationOperator3d;
