-- File:        ProductDefinitionFormation.cdl
-- Created:     Mon Dec  4 12:02:29 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWProductDefinitionFormation from RWStepBasic

	---Purpose : Read & Write Module for ProductDefinitionFormation

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     ProductDefinitionFormation from StepBasic,
     EntityIterator from Interface

is

	Create returns RWProductDefinitionFormation;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable ProductDefinitionFormation from StepBasic);

	WriteStep (me; SW : in out StepWriter; ent : ProductDefinitionFormation from StepBasic);

	Share(me; ent : ProductDefinitionFormation from StepBasic; iter : in out EntityIterator);

end RWProductDefinitionFormation;
