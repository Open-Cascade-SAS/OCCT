-- Created on: 1998-02-27
-- Created by: Christian CAILLET
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ModifEditForm  from IFSelect  inherits Modifier

    ---Purpose : This modifier applies an EditForm on the entities selected

uses CString, AsciiString from TCollection,
     InterfaceModel, CopyTool, Protocol from Interface, ContextModif,
     EditForm

is

    Create (editform : EditForm) returns mutable ModifEditForm;
    ---Purpose : Creates a ModifEditForm. It may not change the graph

    EditForm (me) returns EditForm;
    ---Purpose : Returns the EditForm

    Perform (me; ctx  : in out ContextModif;
    	     target   : mutable InterfaceModel;
    	     protocol : Protocol from Interface;
    	     TC       : in out CopyTool);
    ---Purpose : Acts by applying an EditForm to entities, selected or all model

    Label (me) returns AsciiString from TCollection;
    ---Purpose : Returns Label as "Apply EditForm <+ label of EditForm>"

fields

    theedit : EditForm;

end ModifEditForm;
