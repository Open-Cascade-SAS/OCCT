-- Created on: 1998-06-23
-- Created by: Stephanie HUMEAU
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class  GuideTrihedronAC  from  GeomFill   


inherits  TrihedronWithGuide  from  GeomFill  

---Purpose:   Trihedron in  the  case of a sweeping along a guide  curve.
--            defined by curviline  absciss


uses  
    Shape  from  GeomAbs, 
    Array1OfReal   from TColStd, 
    Vec  from  gp,  
    Curve  from  Geom, 
    HCurve  from  Adaptor3d, 
    TrihedronLaw  from  GeomFill, 
    CurvlinFunc from  Approx   

raises
    OutOfRange,  ConstructionError

is 
    Create(guide  :  HCurve  from  Adaptor3d)
    returns  GuideTrihedronAC  from  GeomFill; 

    SetCurve(me:mutable;  C  :  HCurve  from  Adaptor3d) 
    is  redefined; 

    Copy(me)  returns  TrihedronLaw  from  GeomFill          
     is  redefined;
     
    Guide(me)   
    returns  HCurve  from  Adaptor3d 
    is  redefined;      
      
    D0( me : mutable;  
        Param  : Real; 
        Tangent    : out  Vec  from  gp; 
        Normal     : out  Vec  from  gp;  
        BiNormal   : out  Vec  from  gp)        
    returns Boolean  is  redefined;    

    D1( me : mutable;  
        Param  : Real; 
        Tangent    : out  Vec  from  gp; 
    	DTangent   : out  Vec  from  gp; 
        Normal     : out  Vec  from  gp;  
        DNormal    : out  Vec  from  gp;  
        BiNormal   : out  Vec  from  gp; 
        DBiNormal  : out  Vec  from  gp)        
    returns Boolean  is  redefined;  
    
    D2( me : mutable;  
        Param  : Real; 
        Tangent    : out  Vec  from  gp; 
    	DTangent   : out  Vec  from  gp; 
    	D2Tangent  : out  Vec  from  gp; 
        Normal     : out  Vec  from  gp;  
        DNormal    : out  Vec  from  gp;  
        D2Normal   : out  Vec  from  gp;  
        BiNormal   : out  Vec  from  gp; 
        DBiNormal  : out  Vec  from  gp; 
        D2BiNormal : out  Vec  from  gp)        
    returns Boolean  is  redefined;  

       
--
--  =================== Management  of  continuity  ===================
--                 
    NbIntervals(me; S : Shape from GeomAbs) 
	---Purpose: Returns  the number  of  intervals for  continuity
	--          <S>. 
        --          May be one if Continuity(me) >= <S>
    returns Integer  is  redefined;
 
    Intervals(me; T : in out Array1OfReal from TColStd; 
    	         S : Shape from GeomAbs)
	---Purpose: Stores in <T> the  parameters bounding the intervals
	--          of continuity <S>.
	--          
	--          The array must provide  enough room to  accomodate
	--          for the parameters. i.e. T.Length() > NbIntervals()
    raises
    	OutOfRange from Standard 
    is redefined;  

    SetInterval(me: mutable; First, Last: Real from Standard)    
	---Purpose: Sets the bounds of the parametric interval on 
	--          the function
	--          This determines the derivatives in these values if the
	--          function is not Cn.
   is redefined; 
   
--  ===================  To help   computation of  Tolerance   ===============	 
    GetAverageLaw(me  :  mutable;
      ATangent    : out  Vec  from  gp; 
      ANormal     : out  Vec  from  gp; 
      ABiNormal   : out  Vec  from  gp) 
     ---Purpose: Get average value of M(t) and V(t) it is usfull to 
     --          make fast approximation of rational  surfaces.        
  is  redefined;

--   =================== To help Particular case   ===============	 
    IsConstant(me) 
    ---Purpose: Say if the law is Constant

    --          Return False by Default.        
    returns  Boolean   
    is redefined;  
     
     
    IsOnlyBy3dCurve(me) 
     ---Purpose: Say if the law is defined, only by the 3d Geometry of
     --          the setted Curve  
     --          Return False by Default.        
    returns  Boolean   
    is redefined;           

    Origine(me  :  mutable; 
    	    OrACR1  :  Real; 
    	    OrACR2  :  Real) 
    is  redefined;

fields 
    myGuideAC   :   CurvlinFunc from  Approx; 
    Lguide      :   Real  from  Standard; 
    myCurveAC   :   CurvlinFunc from  Approx; 
    L           :   Real  from  Standard;  
    myCurve     :   HCurve from  Adaptor3d;  
    UTol,  STol :   Real;     
    Orig1  :  Real  from  Standard;
    Orig2  :  Real  from  Standard;
end  GuideTrihedronAC; 
