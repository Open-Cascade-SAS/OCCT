-- Created on: 1994-02-14
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred generic class CSFunction from IntImp 
    (ThePSurface as any;
     TheCurve as any
    )
    
inherits FunctionSetWithDerivatives from math

      	---Purpose: This class is the template function for the intersection
      	--          between a curve and a surface.
      	--          It is possible to implement such a function with an
      	--          instantiation of :
      	--           - ZerCSParFunc for the intersection between a 3d curve
      	--             and a surface.
      	--           - ZerCOnSSParFunc for the intersection between a curve
      	--             on surface and another surface.
    	

uses Vector from math,
     Matrix from math,
     Pnt from gp

is
	    
    NbVariables(me) returns Integer from Standard
    ---Purpose: Returns 3.
    is static;
    
    NbEquations(me) returns Integer from Standard
    ---Purpose: Returns 3.
    is static;
    
    Value(me : in out; X : in Vector from math;
    	    	       F : out Vector from math)
    returns Boolean from Standard
    is static;
    
    Derivatives(me : in out;X : in  Vector from math;
    	    	    	    D : out Matrix from math)
    returns Boolean from Standard
    is static;
    
    Values(me : in out;
    	   X  : in Vector from math;
	   F  : out Vector from math; D: out Matrix from math)
    returns Boolean from Standard
    is static;

    Point(me)
    	---C++: return const&
    	returns Pnt from gp
    	is static;
    
    Root(me) returns Real from Standard
    is static;
    
    AuxillarSurface(me)
    	---C++: return const&
    	returns ThePSurface
    	is static;

    AuxillarCurve(me)
    	---C++: return const&
    	returns TheCurve
    	is static;
     
end CSFunction;
