-- Created on: 1992-08-24
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



package IntSurf 

	---Purpose: This package provides resources for
	--          all the packages concerning the intersection
	--          between surfaces. 

        ---Level: Internal
        --
        -- All the methods of all the classes of this package are Internal.
        -- 


uses Standard, MMgt, StdFail, GeomAbs, TCollection, gp, TColgp

is

    class PntOn2S;
    
    imported Allocator;
    
    imported SequenceOfPntOn2S;

    class Couple;

    class SequenceOfCouple instantiates Sequence from TCollection
                (Couple from IntSurf);
    
    
    class LineOn2S;
    
    class Quadric;
    
    class QuadricTool;
    
    class PathPoint;
    
    class SequenceOfPathPoint instantiates Sequence from TCollection
    	(PathPoint from IntSurf);

    class PathPointTool;
    
    class InteriorPoint;
    
    class SequenceOfInteriorPoint instantiates Sequence from TCollection
    	(InteriorPoint from IntSurf);
    
    class InteriorPointTool;

    class Transition;    

    --amv    
    class ListOfPntOn2S instantiates List from TCollection
    	(PntOn2S from IntSurf);
    
    enumeration TypeTrans is In, Out, Touch, Undecided;
    
    enumeration Situation is Inside, Outside, Unknown;


    MakeTransition(TgFirst,TgSecond: Vec from gp; Normal: Dir from gp;
                   TFirst,TSecond: out Transition from IntSurf);

	---Purpose: Computes the transition of the intersection point
	--          between the two lines.
	--          TgFirst is the tangent vector of the first line.
	--          TgSecond is the tangent vector of the second line.
	--          Normal is the direction used to orientate the cross
	--          product TgFirst^TgSecond.
	--          TFirst is the transition of the point on the first line.
	--          TSecond is the transition of the point on the second line.


end IntSurf;
