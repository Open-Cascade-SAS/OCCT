-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Torus from StepShape 

inherits GeometricRepresentationItem from StepGeom

uses

	Axis1Placement from StepGeom,
	Real from Standard, 
	HAsciiString from TCollection
is

	Create returns mutable Torus;
	---Purpose: Returns a Torus


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aPosition : mutable Axis1Placement from StepGeom;
	      aMajorRadius : Real from Standard;
	      aMinorRadius : Real from Standard) is virtual;

	-- Specific Methods for Field Data Access --

	SetPosition(me : mutable; aPosition : mutable Axis1Placement);
	Position (me) returns mutable Axis1Placement;
	SetMajorRadius(me : mutable; aMajorRadius : Real);
	MajorRadius (me) returns Real;
	SetMinorRadius(me : mutable; aMinorRadius : Real);
	MinorRadius (me) returns Real;

fields

	position : Axis1Placement from StepGeom;
	majorRadius : Real from Standard;
	minorRadius : Real from Standard;

end Torus;
