-- Created on: 1999-09-24
-- Created by: Sergey ZARITCHNY
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class TopNaming from QANewBRepNaming 

    ---Purpose: The root class for all the primitives, features, ...

uses 
 
    Label from TDF

is 
 
    Initialize;

    Initialize(Label : Label from TDF); 
     
    ResultLabel(me) returns Label from TDF; 
    ---C++: inline  
    ---C++: return const& 
    ---Purpose : Returns the result label. 
    
fields  

    myResultLabel : Label from TDF  is  protected; 
      
end TopNaming;
