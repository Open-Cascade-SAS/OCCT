-- File:        ConnectedFaceSet.cdl
-- Created:     Mon Dec  4 12:02:24 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWConnectedFaceSet from RWStepShape

	---Purpose : Read & Write Module for ConnectedFaceSet

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     ConnectedFaceSet from StepShape,
     EntityIterator from Interface

is

	Create returns RWConnectedFaceSet;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable ConnectedFaceSet from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : ConnectedFaceSet from StepShape);

	Share(me; ent : ConnectedFaceSet from StepShape; iter : in out EntityIterator);

end RWConnectedFaceSet;
