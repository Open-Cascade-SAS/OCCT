-- Created on: 1993-06-03
-- Created by: fid
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



package PColPGeom 

        ---Purpose : This package  is used to  instantiate of  several
        --         generic classes from  the package  PCollection with
        --         objects from the package PGeom.

uses PCollection, PGeom

is


    class HArray1OfCurve 
    	instantiates HArray1 from PCollection (Curve from PGeom);
    class HArray1OfBoundedCurve 
    	instantiates HArray1 from PCollection (BoundedCurve from PGeom);
    class HArray1OfBezierCurve 
    	instantiates HArray1 from PCollection (BezierCurve from PGeom);
    class HArray1OfBSplineCurve 
    	instantiates HArray1 from PCollection (BSplineCurve from PGeom);
    class HArray1OfSurface 
    	instantiates HArray1 from PCollection (Surface from PGeom);
    class HArray1OfBoundedSurface 
    	instantiates HArray1 from PCollection (BoundedSurface from PGeom);



    class HArray2OfSurface 
    	instantiates HArray2 from PCollection (Surface from PGeom);
    class HArray2OfBoundedSurface 
    	instantiates HArray2 from PCollection (BoundedSurface from PGeom);
    class HArray2OfBezierSurface 
    	instantiates HArray2 from PCollection (BezierSurface from PGeom);
    class HArray2OfBSplineSurface 
    	instantiates HArray2 from PCollection (BSplineSurface from PGeom);



--    class HSequenceOfCurve  
--    	instantiates HSequence from PCollection (Curve from PGeom);
--    class HSequenceOfBoundedCurve  
--    	instantiates HSequence from PCollection (BoundedCurve from PGeom);
--    class HSequenceOfSurface 
--    	instantiates HSequence from PCollection (Surface from PGeom);
--    class HSequenceOfBoundedSurface 
--    	instantiates HSequence from PCollection (BoundedSurface from PGeom);


end PColPGeom;
