-- Created on: 1995-12-04
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.





package RWStepAP214 

uses

	StepData, Interface, TCollection, TColStd, StepAP214

is


class ReadWriteModule;

class GeneralModule;

class RWAutoDesignActualDateAndTimeAssignment;
class RWAutoDesignActualDateAssignment;
class RWAutoDesignApprovalAssignment;
class RWAutoDesignDateAndPersonAssignment;
class RWAutoDesignGroupAssignment;
class RWAutoDesignNominalDateAndTimeAssignment;
class RWAutoDesignNominalDateAssignment;
class RWAutoDesignOrganizationAssignment;
class RWAutoDesignPersonAndOrganizationAssignment;
class RWAutoDesignPresentedItem;
class RWAutoDesignSecurityClassificationAssignment;
-- Removed from Rev2 to Rev4 : class RWAutoDesignViewArea;

-- Added from STEP214-CC1 to CC2
class RWAutoDesignDocumentReference;
--Added from CC2 to DIS

class RWAppliedDateAndTimeAssignment;
class RWAppliedDateAssignment;
class RWAppliedApprovalAssignment;
class RWAppliedGroupAssignment;
class RWAppliedOrganizationAssignment;
class RWAppliedPersonAndOrganizationAssignment;
class RWAppliedPresentedItem;
class RWAppliedSecurityClassificationAssignment;
class RWAppliedDocumentReference;

-- added for external references (CAX-IF TRJ4)
class RWAppliedExternalIdentificationAssignment;
class RWClass;
class RWExternallyDefinedClass;
class RWExternallyDefinedGeneralProperty;
class RWRepItemGroup;

	Init;
	---Purpose: enforced the initialisation of the  libraries

end RWStepAP214;
