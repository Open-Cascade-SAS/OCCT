-- Created on: 2004-05-20
-- Created by: Sergey ZARITCHNY <szy@opencascade.com>
-- Copyright (c) 2004-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class CurveSet from BinTools 

	---Purpose: Stores a set of Curves from Geom in binary format.

uses
    Curve from Geom,
    IndexedMapOfTransient from TColStd
    
raises
    OutOfRange from Standard

is

    Create returns CurveSet from BinTools;
	---Purpose: Returns an empty set of Curves.
	
    Clear(me : in out)
	---Purpose: Clears the content of the set.
    is static;
	
    Add(me : in out; C : Curve from Geom) returns Integer
	---Purpose: Incorporate a new Curve in the  set and returns
	--          its index.
    is static;
    
    Curve(me; I : Integer) returns Curve from Geom
	---Purpose: Returns the Curve of index <I>.
    raises
    	OutOfRange from Standard
    is static;

    Index(me; C : Curve from Geom) returns Integer
	---Purpose: Returns the index of <L>.
    is static;
    	
    Write(me; OS : in out OStream)
	---Purpose: Writes the content of  me  on the stream <OS> in a
	--          format that can be read back by Read.
    is static;
	
    Read(me : in out; IS : in out IStream)
	---Purpose: Reads the content of me from the  stream  <IS>. me
	--          is first cleared.
	--          
    is static;
	
    --
    -- 	class methods to write an read curves
    -- 	
    
    WriteCurve(myclass; C  : Curve from Geom;
    	    	    	OS : in out OStream);
	---Purpose: Dumps the curve on the stream in binary format
	--          that can be read back.
	
    ReadCurve(myclass; IS : in out IStream;
    	    	       C  : in out Curve from Geom)
    returns IStream;
	---Purpose: Reads the curve  from  the stream.  The  curve  is
	--          assumed  to have  been  written  with  the Write
	--          method
	--          
	---C++: return &
	
fields

    myMap : IndexedMapOfTransient from TColStd;

end CurveSet;
