-- Created on: 2000-08-11
-- Created by: data exchange team
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Driver from XCAFPrs inherits Driver from TPrsStd

    ---Purpose: Implements a driver for presentation of shapes in DECAF 
    --          document. Its the only purpose is to initialize and return 
    --          XCAFPrs_AISObject object on request

uses
    Label             from TDF,
    InteractiveObject from AIS

is

    Update (me : mutable ; L   :        Label from TDF;
	                   ais : in out InteractiveObject from AIS)
    returns Boolean from Standard is redefined;

    GetID (myclass) returns GUID;
    	---Purpose: returns GUID of the driver
	---C++: return const &
    
end Driver;
