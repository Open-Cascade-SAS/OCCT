-- File:	IGESSolid_ToolSelectedComponent.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolSelectedComponent  from IGESSolid

    ---Purpose : Tool to work on a SelectedComponent. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses SelectedComponent from IGESSolid,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolSelectedComponent;
    ---Purpose : Returns a ToolSelectedComponent, ready to work


    ReadOwnParams (me; ent : mutable SelectedComponent;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : SelectedComponent;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : SelectedComponent;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a SelectedComponent <ent>, from
    --           its specific (own) parameters

    DirChecker (me; ent : SelectedComponent) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : SelectedComponent;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : SelectedComponent; entto : mutable SelectedComponent;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : SelectedComponent;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolSelectedComponent;
