-- File:	RWStepFEA_RWParametricSurface3dElementCoordinateSystem.cdl
-- Created:	Thu Dec 12 17:51:07 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWParametricSurface3dElementCoordinateSystem from RWStepFEA

    ---Purpose: Read & Write tool for ParametricSurface3dElementCoordinateSystem

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    ParametricSurface3dElementCoordinateSystem from StepFEA

is
    Create returns RWParametricSurface3dElementCoordinateSystem from RWStepFEA;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : ParametricSurface3dElementCoordinateSystem from StepFEA);
	---Purpose: Reads ParametricSurface3dElementCoordinateSystem

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: ParametricSurface3dElementCoordinateSystem from StepFEA);
	---Purpose: Writes ParametricSurface3dElementCoordinateSystem

    Share (me; ent : ParametricSurface3dElementCoordinateSystem from StepFEA;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWParametricSurface3dElementCoordinateSystem;
