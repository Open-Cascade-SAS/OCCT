-- Created on: 1999-06-24
-- Created by: Sergey ZARITCHNY
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class TranslateTool from TNaming inherits  TShared from MMgt

	---Purpose: The TranslateTool class is provided to support the          
        --          translation of topological data structures  Transient 
    	--  .       to  Transient.

uses 
     Shape                  from TopoDS, 
     IndexedDataMapOfTransientTransient  from TColStd 
      
raises

    TypeMismatch from Standard 
    
is

    Add(me;
    	S1 : in out Shape from TopoDS;
    	S2 :        Shape from TopoDS)
	---Level: Internal 
    raises
    	TypeMismatch from Standard;
    
    --
    --       The Make methods should create a new empty  object of the
    --       given type with  the given Model.   They should raise the
    --       TypeMismatch   exception  if  the Model   is  not of  the
    --       expected type.
    --       


    MakeVertex(me; 
    	       S  : out Shape from TopoDS) 
	---Level: Internal 
    raises
    	TypeMismatch from Standard;
    
    MakeEdge(me; 
    	     S  : out Shape from TopoDS) 
	---Level: Internal 
    raises
    	TypeMismatch from Standard;
    
    MakeWire(me; 
    	     S  : out Shape from TopoDS) 
	---Level: Internal 
    raises
    	TypeMismatch from Standard;
    
    MakeFace(me; 
    	     S  : out Shape from TopoDS) 
	---Level: Internal 
    raises
    	TypeMismatch from Standard;
    
    MakeShell(me; 
    	      S  : out Shape from TopoDS) 
	---Level: Internal 
    raises
    	TypeMismatch from Standard;
    
    MakeSolid(me; 
    	      S  : out Shape from TopoDS) 
	---Level: Internal 
    raises
    	TypeMismatch from Standard;
    
    MakeCompSolid(me; 
    	    	  S  : out Shape from TopoDS) 
	---Level: Internal 
    raises
    	TypeMismatch from Standard;
    
    MakeCompound(me; 
    	    	 S  : out Shape from TopoDS) 
	---Level: Internal 
    raises
    	TypeMismatch from Standard;
    
    --
    --     The Update methods should transfer the data from  the first
    --     shape to the second.
    --     
    
    UpdateVertex(me;
    	         S1 :         Shape                  from TopoDS;
		 S2 : in out  Shape                  from TopoDS;
		 M  : in out  IndexedDataMapOfTransientTransient  from TColStd);
	---Level: Internal 
        
    UpdateEdge  (me;
    	         S1 :         Shape                  from TopoDS;
	         S2 : in out  Shape                  from TopoDS;
	         M  : in out  IndexedDataMapOfTransientTransient  from TColStd);
	---Level: Internal 
    
    UpdateFace  (me;
    	         S1 :         Shape                  from TopoDS;
	         S2 : in out  Shape                  from TopoDS;
	         M  : in out  IndexedDataMapOfTransientTransient  from TColStd);
	---Level: Internal  
    UpdateShape (me; 
    	    	 S1 :         Shape                  from TopoDS;
	         S2 : in out  Shape                  from TopoDS); 
	---Level: Internal 
	     
end TranslateTool;
