-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ViewVolume from StepVisual 

inherits TShared from MMgt

uses

	CentralOrParallel from StepVisual, 
	CartesianPoint from StepGeom, 
	Real from Standard, 
	Boolean from Standard, 
	PlanarBox from StepVisual
is

	Create returns ViewVolume;
	---Purpose: Returns a ViewVolume

	Init (me : mutable;
	      aProjectionType : CentralOrParallel from StepVisual;
	      aProjectionPoint : CartesianPoint from StepGeom;
	      aViewPlaneDistance : Real from Standard;
	      aFrontPlaneDistance : Real from Standard;
	      aFrontPlaneClipping : Boolean from Standard;
	      aBackPlaneDistance : Real from Standard;
	      aBackPlaneClipping : Boolean from Standard;
	      aViewVolumeSidesClipping : Boolean from Standard;
	      aViewWindow : PlanarBox from StepVisual) is virtual;

	-- Specific Methods for Field Data Access --

	SetProjectionType(me : mutable; aProjectionType : CentralOrParallel);
	ProjectionType (me) returns CentralOrParallel;
	SetProjectionPoint(me : mutable; aProjectionPoint : CartesianPoint);
	ProjectionPoint (me) returns CartesianPoint;
	SetViewPlaneDistance(me : mutable; aViewPlaneDistance : Real);
	ViewPlaneDistance (me) returns Real;
	SetFrontPlaneDistance(me : mutable; aFrontPlaneDistance : Real);
	FrontPlaneDistance (me) returns Real;
	SetFrontPlaneClipping(me : mutable; aFrontPlaneClipping : Boolean);
	FrontPlaneClipping (me) returns Boolean;
	SetBackPlaneDistance(me : mutable; aBackPlaneDistance : Real);
	BackPlaneDistance (me) returns Real;
	SetBackPlaneClipping(me : mutable; aBackPlaneClipping : Boolean);
	BackPlaneClipping (me) returns Boolean;
	SetViewVolumeSidesClipping(me : mutable; aViewVolumeSidesClipping : Boolean);
	ViewVolumeSidesClipping (me) returns Boolean;
	SetViewWindow(me : mutable; aViewWindow : PlanarBox);
	ViewWindow (me) returns PlanarBox;

fields

	projectionType : CentralOrParallel from StepVisual; -- an Enumeration
	projectionPoint : CartesianPoint from StepGeom;
	viewPlaneDistance : Real from Standard;
	frontPlaneDistance : Real from Standard;
	frontPlaneClipping : Boolean from Standard;
	backPlaneDistance : Real from Standard;
	backPlaneClipping : Boolean from Standard;
	viewVolumeSidesClipping : Boolean from Standard;
	viewWindow : PlanarBox from StepVisual;

end ViewVolume;
