-- File:	GeomFill_Curved.cdl
-- Created:	Tue Sep 28 16:24:04 1993
-- Author:	Bruno DUMORTIER
--		<dub@sdsun1>
---Copyright:	 Matra Datavision 1993

class Curved from GeomFill inherits Filling from GeomFill

uses
    Array1OfPnt  from TColgp,
    Array1OfReal from TColStd

is
    Create;
    
    Create(P1, P2, P3, P4 : Array1OfPnt from TColgp)
    returns Curved from GeomFill;
    
    Create(P1, P2, P3, P4 : Array1OfPnt  from TColgp;
    	   W1, W2, W3, W4 : Array1OfReal from TColStd)
    returns Curved from GeomFill;
    

    Create(P1, P2, P3 : Array1OfPnt from TColgp)
    returns Curved from GeomFill;
    
    Create(P1, P2, P3 : Array1OfPnt  from TColgp;
    	   W1, W2, W3 : Array1OfReal from TColStd)
    returns Curved from GeomFill;
    

    Create(P1, P2 : Array1OfPnt from TColgp)
    returns Curved from GeomFill;
    
    Create(P1, P2 : Array1OfPnt  from TColgp;
    	   W1, W2 : Array1OfReal from TColStd)
    returns Curved from GeomFill;
    

    Init(me : in out;
    	 P1, P2, P3, P4 : Array1OfPnt from TColgp)
    is static;

    Init(me : in out;
    	 P1, P2, P3, P4 : Array1OfPnt  from TColgp;
    	 W1, W2, W3, W4 : Array1OfReal from TColStd)
    is static;

    Init(me : in out;
    	 P1, P2, P3 : Array1OfPnt from TColgp)
    is static;

    Init(me : in out;
    	 P1, P2, P3 : Array1OfPnt  from TColgp;
    	 W1, W2, W3 : Array1OfReal from TColStd)
    is static;

    Init(me : in out;
    	 P1, P2 : Array1OfPnt from TColgp)
    is static;

    Init(me : in out;
    	 P1, P2 : Array1OfPnt  from TColgp;
    	 W1, W2 : Array1OfReal from TColStd)
    is static;

end Curved;
