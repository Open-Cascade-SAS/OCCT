-- Created on: 1999-11-26
-- Created by: Andrey BETENEV
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0

class RWCurveBoundedSurface from RWStepGeom

    ---Purpose: Read & Write tool for CurveBoundedSurface

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    CurveBoundedSurface from StepGeom

is
    Create returns RWCurveBoundedSurface from RWStepGeom;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : CurveBoundedSurface from StepGeom);
	---Purpose: Reads CurveBoundedSurface

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: CurveBoundedSurface from StepGeom);
	---Purpose: Writes CurveBoundedSurface

    Share (me; ent : CurveBoundedSurface from StepGeom;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWCurveBoundedSurface;
