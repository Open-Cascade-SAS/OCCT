-- Created on: 1995-03-02
-- Created by: Christian CAILLET
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class AddGroup  from IGESSelect  inherits ModelModifier from IGESSelect

    ---Purpose : Adds a Group to contain the entities designated by the
    --           Selection. If no Selection is given, nothing is done

uses AsciiString from TCollection,
     IGESModel, CopyTool, ContextModif

is

    Create returns mutable AddGroup;
    ---Purpose : Creates an AddGroup

    Performing (me; ctx : in out ContextModif;
    	        target  : mutable IGESModel;
                TC      : in out CopyTool);
    ---Purpose : Specific action : Adds a new group

    Label (me) returns AsciiString from TCollection;
    ---Purpose : Returns a text which is
    --           "Add Group"

end AddGroup;
