-- Created on: 2001-11-02
-- Created by: Peter KURNEV
-- Copyright (c) 2001-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class BuilderTools from BOP 

    ---Purpose: 
    	--  Some  handy tools used by classes    
	--  BOP_ShellShell, 
	--  BOP_ShellSolid, 
	--  BOP_SolidSolid  
	--  to build a result  

uses
  
    IndexedMapOfInteger from TColStd,  
     
    State     from TopAbs,  
    ShapeEnum from TopAbs, 
     
    Face from TopoDS, 
    Edge from TopoDS,   
     
    ListOfShape from TopTools, 
      
    StateOfShape from BooleanOperations, 
      
    IndexedDataMapOfIntegerIndexedMapOfInteger from BOPTColStd, 	
     
    CArray1OfSSInterference from BOPTools,  
     
    Operation            from BOP,
    ListOfConnexityBlock from BOP     
    
    
is

    StateToCompare(myclass; 
	    iRank :Integer from Standard; 
	    anOp  :Operation from BOP) 
	returns StateOfShape from BooleanOperations;  
    
    ToReverseSection(myclass; 
	    iRank :Integer from Standard; 
	    anOp  :Operation from BOP) 
	returns Boolean from Standard;   
	 
    ToReverseFace(myclass; 
	    iRank :Integer from Standard; 
	    anOp  :Operation from BOP) 
	returns Boolean from Standard;  
	 
    OrientSectionEdgeOnF1(myclass; 
	    aF1   :Face from TopoDS; 
	    aF2   :Face from TopoDS;  
    	    iRank :Integer from Standard;  
	    anOp  :Operation from BOP;
	    aE    :out Edge from TopoDS); 
	 
    IsSameDomainFaceWithF1(myclass; 
    	    nF1 :Integer from Standard; 
    	    nF2 :Integer from Standard; 
    	    aFFM:IndexedMapOfInteger from TColStd; 
	    aFFs:out CArray1OfSSInterference from BOPTools)  
	returns Boolean from Standard;     

    IsPartIN2DToKeep(myclass;  
    	    aSt   :State from TopAbs;
	    iRank :Integer from Standard;  
	    anOp  :Operation from BOP)	
	returns Boolean from Standard;   	 

    IsPartOn2dToKeep(myclass;  
    	    aSt   :State from TopAbs;
	    iRank :Integer from Standard;  
	    anOp  :Operation from BOP)	
	returns Boolean from Standard;  
	 
    DoMap(myclass;  
    	    aFFs  :out  CArray1OfSSInterference from BOPTools; 
    	    aFFMap:out  IndexedDataMapOfIntegerIndexedMapOfInteger from BOPTColStd);      

    MakeConnexityBlocks(myclass;  
    	    aLE        :  ListOfShape from TopTools;  
	    aType      :  ShapeEnum   from TopAbs;  
	    aLConBlks  : out ListOfConnexityBlock from BOP); 

end BuilderTools;
