-- Created on: 2001-04-24
-- Created by: Christian CAILLET
-- Copyright (c) 2001-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MeasureQualification  from StepShape    inherits TShared

    ---Purpose : Added for Dimensional Tolerances

uses
    HAsciiString from TCollection,
    MeasureWithUnit from StepBasic,
    ValueQualifier from StepShape,
    HArray1OfValueQualifier from StepShape

is

    Create returns mutable MeasureQualification;

    Init (me : mutable; name : HAsciiString from TCollection;
    	    description : HAsciiString from TCollection;
	    qualified_measure : MeasureWithUnit from StepBasic;
	    qualifiers : HArray1OfValueQualifier from StepShape);

    Name (me) returns HAsciiString from TCollection;
    SetName (me : mutable; name : HAsciiString from TCollection);

    Description (me) returns HAsciiString from TCollection;
    SetDescription (me : mutable; description : HAsciiString from TCollection);

    QualifiedMeasure (me) returns MeasureWithUnit from StepBasic;
    SetQualifiedMeasure (me : mutable; qualified_measure : MeasureWithUnit from StepBasic);

    Qualifiers (me) returns HArray1OfValueQualifier from StepShape;
    NbQualifiers (me) returns Integer;
    SetQualifiers (me : mutable; qualifiers : HArray1OfValueQualifier from StepShape);
    QualifiersValue (me; num : Integer) returns ValueQualifier from StepShape;
    SetQualifiersValue (me : mutable; num : Integer; aqualifier : ValueQualifier from StepShape);

fields

    theName : HAsciiString from TCollection;
    theDescription : HAsciiString from TCollection;
    theQualifiedMeasure : MeasureWithUnit from StepBasic;
    theQualifiers : HArray1OfValueQualifier from StepShape;

end MeasureQualification;
