-- Created on: 1996-04-01
-- Created by: Philippe MANGIN
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

private class DistributionOfJerk from FairCurve inherits  DistributionOfEnergy  from FairCurve

	---Purpose: Compute the "Jerk" distribution.

uses  Vector        from math, 
      FunctionSet   from math,
      HArray1OfReal  from TColStd,
      HArray1OfPnt2d from TColgp,
      BattenLaw  from FairCurve


is
    Create( BSplOrder :  Integer;
            FlatKnots :  HArray1OfReal;
	    Poles     :  HArray1OfPnt2d;
	    DerivativeOrder : Integer; 
	    Law       :  BattenLaw;
            NbValAux  : Integer = 0) returns DistributionOfJerk;
	    

    Value(me: in out; X: Vector; F: out Vector)
    	---Purpose: computes the values <F> of the functions for the 
    	--          variable <X>.
    	--          returns True if the computation was done successfully, 
    	--          False otherwise.

    returns Boolean is redefined;
    

fields
    MyLaw           : BattenLaw;
end DistributionOfJerk;
