-- Created on: 1998-12-29
-- Created by: Joelle CHAUVET
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class NSections from BRepFill inherits  SectionLaw  from  BRepFill

	---Purpose: Build Section Law, with N Sections
	--          
        ---Level: Advanced
       
uses 
 SectionLaw          from  GeomFill,  
 HArray1OfSectionLaw from  GeomFill,
 SequenceOfTrsf      from  GeomFill,
 BSplineSurface      from  Geom, 
 HArray2OfShape      from  TopTools,  
 SequenceOfReal      from  TColStd,  
 SequenceOfShape     from  TopTools,  
 Shape               from  GeomAbs,
 Vertex              from  TopoDS, 
 Wire                from  TopoDS,  
 Edge                from  TopoDS,  
 Shape               from  TopoDS, 
 Function            from  Law

is  
  Create (S:SequenceOfShape  from  TopTools;   
          Build :  Boolean = Standard_True)   
     ---Purpose: Construct    
  returns NSections from BRepFill;  
   
  Create (S      :  SequenceOfShape from  TopTools; 
  	  Trsfs  :  SequenceOfTrsf  from  GeomFill; 
  	  P      :  SequenceOfReal  from  TColStd; 
	  VF,VL  :  Real; 
          Build  :  Boolean = Standard_True)   
     ---Purpose: Construct    
  returns NSections from BRepFill;  
   

  IsVertex(me) 
    ---Purpose: Say if the input shape is a  vertex. 
  returns  Boolean   
  is  redefined; 
   
  IsConstant(me) 
    ---Purpose: Say if the Law is  Constant.        
  returns  Boolean   
  is  redefined;        

  ConcatenedLaw(me)  
   ---Purpose: Give the law build on a concatened section         
  returns SectionLaw from GeomFill 
  is  redefined;    
  
  Continuity(me; Index  :  Integer; 
    	         TolAngular  :  Real)
  returns  Shape  from  GeomAbs  
  is  redefined;  
   
  VertexTol(me; Index  :  Integer;   
                Param  :  Real) 
  returns  Real   
  is  redefined;  
  
  Vertex(me;  Index  :  Integer; 
              Param  :  Real) 
  returns Vertex  from  TopoDS 
  is  redefined;	    
   
  D0(me:mutable;  Param  :  Real;   
     S  :  out  Shape  from  TopoDS)   
    is  redefined;  
   
  Init(me  :  mutable;  P  : SequenceOfReal  from  TColStd; 
    	    	    	B  : Boolean  from  Standard )  is  private;
   
fields
  VFirst,  VLast : Real;
  myShapes:  SequenceOfShape  from  TopTools;
  myTrsfs:   SequenceOfTrsf   from  GeomFill;
  myParams:  SequenceOfReal   from  TColStd;   
  myEdges:  HArray2OfShape from  TopTools;   
  mySurface:  BSplineSurface from  Geom;   
end NSections;
