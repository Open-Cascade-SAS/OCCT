-- Created on: 1993-09-28
-- Created by: Bruno DUMORTIER
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Filling from GeomFill


uses
    Array1OfPnt    from TColgp,
    Array2OfPnt    from TColgp,
    HArray2OfPnt   from TColgp,
    Array1OfReal   from TColStd,
    Array2OfReal   from TColStd,
    HArray2OfReal  from TColStd
    
raises
    NoSuchObject from Standard

is
    Create;
    
    NbUPoles(me) returns Integer from Standard
    is static;
    
    NbVPoles(me) returns Integer from Standard
    is static;

    Poles(me; Poles : in out Array2OfPnt from TColgp)
    is static;
    
    isRational(me) returns Boolean from Standard
    is static;
    
    Weights(me; Weights : in out Array2OfReal from TColStd)
    raises
    	NoSuchObject from Standard
    is static;    
    
    
fields
    
    IsRational : Boolean        from Standard is protected;
    myPoles    : HArray2OfPnt   from TColgp   is protected;
    myWeights  : HArray2OfReal  from TColStd  is protected;

end Filling;
