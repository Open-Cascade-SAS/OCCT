-- File:	 SphereToBSplineSurface.cdl
-- Created:	 Thu Oct 10 15:43:43 1991
-- Author:	 Jean Claude VAUTHIER
---Copyright:	 Matra Datavision 1991, 1992





class SphereToBSplineSurface   from Convert

        --- Purpose :
        --  This algorithm converts a bounded Sphere into a rational 
        --  B-spline surface. The sphere is a Sphere from package gp. 
        --  The parametrization of the sphere is
        --  P (U, V) = Loc  + Radius * Sin(V) * Zdir +
        --             Radius * Cos(V) * (Cos(U)*Xdir + Sin(U)*Ydir)
        --  where Loc is the center of the sphere Xdir, Ydir and Zdir are the
        --  normalized directions of the local cartesian coordinate system of
        --  the sphere. The parametrization range is U [0, 2PI] and
        --  V [-PI/2, PI/2].
        --- KeyWords :
        --  Convert, Sphere, BSplineSurface.

inherits ElementarySurfaceToBSplineSurface

uses Sphere from gp

raises DomainError from Standard

is

  Create (Sph : Sphere; U1, U2, V1, V2 : Real)  returns SphereToBSplineSurface
       --- Purpose : 
       --  The equivalent B-spline surface as the same orientation as the 
       --  sphere in the U and V parametric directions.
     raises DomainError;
       --- Purpose :
       --  Raised if U1 = U2 or U1 = U2 + 2.0 * Pi
       --  Raised if V1 = V2.


  Create (Sph : Sphere; 
          Param1, Param2 : Real; 
          UTrim : Boolean = Standard_True) 
        returns SphereToBSplineSurface
       --- Purpose : 
       --  The equivalent B-spline surface as the same orientation
       --  as the sphere in the U and V parametric directions.
     raises DomainError;
       --- Purpose :
       --  Raised if UTrim = True and Param1 = Param2 or 
       --            Param1 = Param2 + 2.0 * Pi
       --  Raised if UTrim = False and Param1 = Param2 


  Create (Sph : Sphere)   returns SphereToBSplineSurface;
       --- Purpose : 
       --  The equivalent B-spline surface as the same orientation
       --  as the sphere in the U and V parametric directions.



end SphereToBSplineSurface;




