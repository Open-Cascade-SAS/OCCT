-- Created on: 1993-06-17
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package TopOpeBRepDS

    ---Purpose: This package provides services used by the TopOpeBRepBuild
    --          package performing topological operations on the BRep
    --          data structure.

uses

    MMgt,
    Standard,
    TopAbs,
    TopoDS,
    TopTools,
    TCollection,
    TColStd,
    TopExp,
    gp,
    BRep,
    Geom,
    Geom2d,
    TopOpeBRepTool,
    
    -- for HDataStructure and relevant classes 
    TopTrans
    
is
    enumeration Kind is 
    POINT,CURVE,SURFACE,VERTEX,EDGE,WIRE,FACE,SHELL,SOLID,COMPSOLID,COMPOUND,UNKNOWN
    end Kind;
    ---Purpose: different types of objects in DataStructure

    enumeration Config is
    UNSHGEOMETRY, SAMEORIENTED, DIFFORIENTED
    end Config;

    enumeration CheckStatus is
    OK,NOK
    end CheckStatus;

    imported DataMapOfCheckStatus;

    imported DataMapIteratorOfDataMapOfCheckStatus;

    class Interference;
    imported ListOfInterference;
    imported ListIteratorOfListOfInterference;
    class InterferenceIterator;
    imported DataMapOfInterferenceListOfInterference;
    imported DataMapIteratorOfDataMapOfInterferenceListOfInterference;

    imported DataMapOfInterferenceShape;

    imported DataMapIteratorOfDataMapOfInterferenceShape;

    imported DataMapOfIntegerListOfInterference;

    imported DataMapIteratorOfDataMapOfIntegerListOfInterference;
    
    imported Array1OfDataMapOfIntegerListOfInterference;

    imported transient class HArray1OfDataMapOfIntegerListOfInterference;
        
    class TKI;
    class Transition;

    class CurvePointInterference;

    class SurfaceCurveInterference;

    class SolidSurfaceInterference;

    class ShapeShapeInterference;

    class EdgeVertexInterference;

    class FaceEdgeInterference;

    class Surface;
    class Curve;
    class Point;
    	
    imported IndexedDataMapOfVertexPoint;

    class GeometryData;
    
    class SurfaceData;
    imported MapOfSurface;
    imported DataMapIteratorOfMapOfSurface;

    class CurveData;
    imported MapOfCurve;
    imported DataMapIteratorOfMapOfCurve;

    class PointData;
    imported MapOfPoint;
    imported DataMapIteratorOfMapOfPoint;

    class ShapeData;
    imported MapOfShapeData;

    imported ShapeSurface;

    imported DataMapIteratorOfShapeSurface;
    
    imported DoubleMapOfIntegerShape;
    
    imported DoubleMapIteratorOfDoubleMapOfIntegerShape; -- for DSS

    imported MapOfIntegerShapeData;

    imported DataMapIteratorOfMapOfIntegerShapeData; -- for DSS

    class DSS; -- (DataStructure Shape) NYI
    
    class DataStructure;
    pointer PDataStructure to DataStructure from TopOpeBRepDS; 
    
    class SurfaceIterator;
    class CurveIterator;
    class PointIterator;

    class SurfaceExplorer;
    class CurveExplorer;
    class PointExplorer;
    
    class InterferenceTool;
    class BuildTool;    
    class Dumper;
    class Marker;
    
    class HDataStructure;
    class EdgeInterferenceTool;
    class Edge3dInterferenceTool;
    class FaceInterferenceTool;

    class Filter;
    class Reducer;
    class TOOL;
    class FIR;
    class EIR;
    class Check;
    
    class GapFiller;
    class GapTool;
    class Association;
    
    class ListOfShapeOn1State;
    imported DataMapOfShapeListOfShapeOn1State;
    imported DataMapIteratorOfDataMapOfShapeListOfShapeOn1State;

    class Explorer;

--modified by NIZNHY-PKV Mon Sep 20 11:49:15 1999  f 
	 
    class  ShapeWithState; 
    imported IndexedDataMapOfShapeWithState; 

    imported DataMapOfShapeState;

    imported DataMapIteratorOfDataMapOfShapeState;
        	 
--modified by NIZNHY-PKV Mon Sep 20 11:49:20 1999  t	     
    




    SPrint(S:State from TopAbs) 
    returns AsciiString from TCollection; ---Purpose: IN OU ON UN
    Print(S:State from TopAbs; OS:in out OStream) returns OStream; ---C++: return &

    SPrint(K:Kind) returns AsciiString from TCollection; ---Purpose: <K>
    SPrint(K:Kind;I:Integer;
    	   B:AsciiString from TCollection = "";A:AsciiString from TCollection = "")
    returns AsciiString from TCollection; ---Purpose: S1(<K>,<I>)S2
    Print(K:Kind;S:in out OStream) returns OStream; ---C++: return &
    Print(K:Kind;I:Integer;S:in out OStream;
    	  B:AsciiString from TCollection = "";A:AsciiString from TCollection = "")
    returns OStream; ---C++: return &

    SPrint(T:ShapeEnum from TopAbs) returns AsciiString from TCollection;
    SPrint(T:ShapeEnum from TopAbs;I:Integer) 
    returns AsciiString from TCollection; ---Purpose: (<T>,<I>)
    Print(T:ShapeEnum from TopAbs;I:Integer;S:in out OStream) returns OStream; ---C++: return &

    SPrint(O:Orientation from TopAbs) returns AsciiString from TCollection;
    SPrint(C:Config) returns AsciiString from TCollection;
    Print(C:Config;S:in out OStream) returns OStream; ---C++: return &

    IsGeometry(K:Kind) returns Boolean;
    IsTopology(K:Kind) returns Boolean;
    KindToShape(K:Kind) returns ShapeEnum from TopAbs;
    ShapeToKind(S:ShapeEnum from TopAbs) returns Kind;

end TopOpeBRepDS;
