-- Created on: 2002-12-14
-- Created by: data exchange team
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class FreedomAndCoefficient from StepFEA
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity FreedomAndCoefficient

uses
    DegreeOfFreedom from StepFEA,
    MeasureOrUnspecifiedValue from StepElement

is
    Create returns FreedomAndCoefficient from StepFEA;
	---Purpose: Empty constructor

    Init (me: mutable; aFreedom: DegreeOfFreedom from StepFEA;
                       aA: MeasureOrUnspecifiedValue from StepElement);
	---Purpose: Initialize all fields (own and inherited)

    Freedom (me) returns DegreeOfFreedom from StepFEA;
	---Purpose: Returns field Freedom
    SetFreedom (me: mutable; Freedom: DegreeOfFreedom from StepFEA);
	---Purpose: Set field Freedom

    A (me) returns MeasureOrUnspecifiedValue from StepElement;
	---Purpose: Returns field A
    SetA (me: mutable; A: MeasureOrUnspecifiedValue from StepElement);
	---Purpose: Set field A

fields
    theFreedom: DegreeOfFreedom from StepFEA;
    theA: MeasureOrUnspecifiedValue from StepElement;

end FreedomAndCoefficient;
