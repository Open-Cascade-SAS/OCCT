-- Created on: 2003-03-05
-- Created by: Sergey KUUL
-- Copyright (c) 2003-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Material from XCAFDoc inherits Attribute from TDF
uses
    Label from TDF,
    RelocationTable from TDF,
    HAsciiString from TCollection

is
    Create returns Material from XCAFDoc;
    
    ---Category: class methods
    --           =============

    GetID (myclass)   
    	---C++: return const &  
    returns GUID from Standard;
    
    Set (myclass; label : Label from TDF;
    	    	  aName : HAsciiString from TCollection;
    	    	  aDescription : HAsciiString from TCollection;
    	    	  aDensity : Real from Standard;
    	    	  aDensName : HAsciiString from TCollection;
    	    	  aDensValType : HAsciiString from TCollection)
    returns Material from XCAFDoc;

    Set (me : mutable; aName : HAsciiString from TCollection;
    	    	       aDescription : HAsciiString from TCollection;
    	    	       aDensity : Real from Standard;
    	    	       aDensName : HAsciiString from TCollection;
    	    	       aDensValType : HAsciiString from TCollection);
	     
    GetName (me) returns HAsciiString from TCollection;

    GetDescription (me) returns HAsciiString from TCollection;

    GetDensity (me) returns Real from Standard;

    GetDensName (me) returns HAsciiString from TCollection;

    GetDensValType (me) returns HAsciiString from TCollection;

    ID (me)
    	---C++: return const & 
    returns GUID from Standard;

    Restore (me: mutable; With : Attribute from TDF);

    NewEmpty (me)
    returns Attribute from TDF;

    Paste (me; Into : Attribute from TDF;
	       RT   : RelocationTable from TDF);    

fields
    myName        : HAsciiString from TCollection;
    myDescription : HAsciiString from TCollection;
    myDensity     : Real from Standard;
    myDensName    : HAsciiString from TCollection;
    myDensValType : HAsciiString from TCollection;

end Material;
