-- Created on: 1993-06-23
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Point from TopOpeBRepDS

    ---Purpose: A Geom point and a tolerance.

uses

    Pnt from gp,
    Shape from TopoDS
    
is

    Create returns Point from TopOpeBRepDS; 

    Create(P : Pnt from gp; T : Real from Standard)
    returns Point from TopOpeBRepDS; 

    Create(S : Shape from TopoDS)
    returns Point from TopOpeBRepDS;

    IsEqual(me; other : Point from TopOpeBRepDS)
    returns Boolean from Standard
    is static;

    Point(me) returns Pnt from gp
    ---C++: return const &
    is static;
    
    ChangePoint(me : in out) returns Pnt from gp
    ---C++: return &
    is static;
    
    Tolerance(me) returns Real from Standard
    is static;

    Tolerance(me : in out; Tol : Real from Standard)
    is static;

    Keep(me) returns Boolean from Standard
    is static;
    ChangeKeep(me : in out; B : Boolean from Standard)
    is static;

fields

    myPoint     : Pnt from gp;
    myTolerance : Real from Standard;
    myKeep      : Boolean from Standard;
    
end Point from TopOpeBRepDS;
