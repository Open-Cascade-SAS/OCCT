-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class LocalTime from StepBasic 

inherits TShared from MMgt

uses

	Integer from Standard, 
	Real from Standard, 
	CoordinatedUniversalTimeOffset from StepBasic, 
	Boolean from Standard
is

	Create returns mutable LocalTime;
	---Purpose: Returns a LocalTime

	Init (me : mutable;
	      aHourComponent : Integer from Standard;
	      hasAminuteComponent : Boolean from Standard;
	      aMinuteComponent : Integer from Standard;
	      hasAsecondComponent : Boolean from Standard;
	      aSecondComponent : Real from Standard;
	      aZone : mutable CoordinatedUniversalTimeOffset from StepBasic) is virtual;

	-- Specific Methods for Field Data Access --

	SetHourComponent(me : mutable; aHourComponent : Integer);
	HourComponent (me) returns Integer;
	SetMinuteComponent(me : mutable; aMinuteComponent : Integer);
	UnSetMinuteComponent (me:mutable);
	MinuteComponent (me) returns Integer;
	HasMinuteComponent (me) returns Boolean;
	SetSecondComponent(me : mutable; aSecondComponent : Real);
	UnSetSecondComponent (me:mutable);
	SecondComponent (me) returns Real;
	HasSecondComponent (me) returns Boolean;
	SetZone(me : mutable; aZone : mutable CoordinatedUniversalTimeOffset);
	Zone (me) returns mutable CoordinatedUniversalTimeOffset;

fields

	hourComponent : Integer from Standard;
	minuteComponent : Integer from Standard;   -- OPTIONAL can be NULL
	secondComponent : Real from Standard;   -- OPTIONAL can be NULL
	zone : CoordinatedUniversalTimeOffset from StepBasic;
	hasMinuteComponent : Boolean from Standard;
	hasSecondComponent : Boolean from Standard;

end LocalTime;
