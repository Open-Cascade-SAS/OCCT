-- Created on: 1994-11-21
-- Created by: CAL
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


-- Modified: TCL G002A, 28-11-00, new section "inquire methods"


class ImageFile from Graphic2d inherits Primitive from Graphic2d

	---Version:

	---Purpose: The primitive ImageFile

	---Keywords: Primitive, ImageFile
	---Warning:
	---References:

uses

	File		from OSD,
	AsciiString	from TCollection,
	Drawer          from Graphic2d,
	GraphicObject	from Graphic2d,
	Factor          from Quantity,
	Length          from Quantity,
	CardinalPoints  from Aspect, 
	FStream         from Aspect,
	IFStream	from Aspect

raises
	ImageDefinitionError from Graphic2d

is
	-------------------------
	-- Category: Constructors
	-------------------------

	Create (aGraphicObject: GraphicObject from Graphic2d;
		aFile: in out File from OSD;
		X, Y: Length from Quantity;
		adx: Length from Quantity = 0.0;
		ady: Length from Quantity = 0.0;
		aTypeOfPlacement: CardinalPoints
				from Aspect = Aspect_CP_Center;
		aScale: Factor from Quantity = 1.0)
	returns mutable ImageFile from Graphic2d
	---Level: Public
	---Purpose: Defines an image with its center location;
	--	    <X>, <Y> defines the position in the space model.
	--	    <adx>, <ady> defines an offset in the device space.
	--	    <ascale> defines a scale factor applied to the
	--	    original size of the image.
	--	    The image will be placed at this offset
	--	    according to the type of placement.
	--
	--	    CardinalPoints values :
	--		- CP_North
	--		- CP_NorthEast
	--		- CP_East
	--		- CP_SouthEast
	--		- CP_South
	--		- CP_SouthWest
	--		- CP_West
	--		- CP_NorthWest
	--		- CP_Center
	raises ImageDefinitionError;
	---Trigger:
	--	If the file don't exist or has a null size.	
	---Category: Constructors

	--------------------------
	-- Category: Draw and Pick
	--------------------------

	Draw (me : mutable; aDrawer: Drawer from Graphic2d)
	is static protected;
	---Level: Internal
	---Purpose: Draws the image at the required center location
	--	    defined by the SetCenter method.
	---Category: Draw and Pick

	Pick (me : mutable;
		X, Y: ShortReal from Standard;
		aPrecision: ShortReal from Standard;
		aDrawer: Drawer from Graphic2d)
	returns Boolean from Standard
	is static protected;
	---Purpose: Returns Standard_True if the image <me> is picked,
	--          Standard_False if not.
	---Category: Draw and Pick

    ---------------------------------------------------
	-- Category: Methods to modify the class definition
	---------------------------------------------------

	SetCenter (me: mutable;
		X, Y: Length from Quantity)
	is static;
	---Level: Public
	---Purpose: Modifies the center location of the image <me>.
	---Category: Methods to modify the class definition

	SetOffset (me: mutable;
		dx, dy: Length from Quantity)
	is static;
	---Level: Public
	---Purpose: Modifies the offset of the image <me>.
	---Category: Methods to modify the class definition

	SetPlacement (me: mutable; aPlacement: CardinalPoints from Aspect)
	is  static;
	---Level: Public
	---Purpose: Modifies the type of placement of the image <me>.
	--
	--	    CardinalPoints values :
	--		- CP_North
	--		- CP_NorthEast
	--		- CP_East
	--		- CP_SouthEast
	--		- CP_South
	--		- CP_SouthWest
	--		- CP_West
	--		- CP_NorthWest
	--		- CP_Center
	---Category: Methods to modify the class definition

	Translate (me: mutable;
	           DX, DY: Length from Quantity)
	is static;
	---Level: Public
	---Purpose: Modifies the center location of the image <me>
	--          by translating it.
	---Category: Methods to modify the class definition

	SetScale (me: mutable; aScale: Factor from Quantity) is static;
	---Level: Public
	---Purpose: Changes the scale factor of the image.
	---Category: Methods to modify the class definition 

	SetZoomable (me: mutable; aFlag: Boolean from Standard = Standard_False)
	is static;
	---Level: Public
	---Purpose: The image <me> follows the scale factor of the view
	--	    if the flag is Standard_True.
	---Category: Zoom management

        Clear (me: mutable) is static; 
        ---Level: Public 
        ---Purpose: Clear the reference to this imagefile if something 
        --         inside have changed,Forced the reload of this at Draw()
        --         time.
        ---Category: Methods to modify the class definition
 
	----------------------------
	-- Category: Zoom management
	----------------------------

	Scale (me)
		returns Factor from Quantity;
	---Level: Internal
	---Purpose: Returns the original scale factor applied to
	--	    the image <me>.
	---Category: Zoom management

	IsZoomable (me)
		returns Boolean from Standard is static;
	---Level: Internal
	---Purpose: Returns Standard_True if the image <me> follows
	--	    the scale factor of the view.
	---Category: Zoom management

	----------------------------
	-- Category: Inquire methods
	----------------------------

    Position( me; X, Y: out Length from Quantity );  
	---Level: Public
	---Purpose: returns the position in the space model
	
	Offset( me; aX, aY: out Length from Quantity );
	---Level: Public
	---Purpose: returns the offset in the device space
	
    Placement( me ) returns CardinalPoints from Aspect;
	---Level: Public
	---Purpose: returns the type of placement
	
	ImageFile( me ) returns File from OSD;
	---Level: Public
	---Purpose: returns the image file


	Values (myclass;
		aFile: in out File from OSD;
		aWidth, aHeight: out Integer from Standard;
		aDepth: out Integer from Standard)
	returns Boolean from Standard;
	---Level: Internal
	---Purpose: Returns Standard_True, the Image pixel size
	--	    and the Image planes depth, if the image file :
	--		- is not open
	--		- exists
	--		- have the extension .xwd
	--	    NOTE that only XWD image file type are recognized.
	---Category: Inquire methods

	----------------------------
	-- Category: Private methods
	----------------------------

	ComputeCenterAndSize (me : mutable;
		aDrawer: Drawer from Graphic2d;
		cx, cy, width, height: out ShortReal from  Standard)
	returns Boolean from Standard is static private;
	---Level: Internal
	---Purpose: Evaluates the center of the image in the device space.
	--	    Called by the methods :
	--		- Graphic2d_ImageFile::Draw
	--		- Graphic2d_ImageFile::Pick
	--		- Graphic2d_ImageFile::FillAndDraw
    	--Returns FALSE if the size cann't gbe evaluated.
	---Category: Private methods

	SwapLong (myclass;
		anAddress: Address from Standard;
		aNumOfBytes: Integer from  Standard);
	---Level: Internal
	---Purpose: Swaps long ints
	---Category: Private methods

	----------------------------------------------------------------------

	Save( me; aFStream: in out FStream from Aspect ) is virtual;
--	Retrieve( me; aIFStream: in out IFStream from AIS2D ) is virtual;

fields

	myFile:		       File from OSD;
	myFileName:	       AsciiString from TCollection;
	myX, myY:	       ShortReal from Standard;
	mydx, mydy:        ShortReal from Standard;
	myWidth, myHeight: Integer from Standard;
	myPlacement:	   CardinalPoints from Aspect;
	myIsZoomable:	   Boolean from Standard;
	myScale:	       ShortReal from Standard;
	myIsModified:	   Boolean from Standard;

end ImageFile from Graphic2d;
