-- Created on: 1996-09-17
-- Created by: Odile Olivier
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class ShapeTypeFilter from StdSelect inherits Filter from SelectMgr

	--- Purpose: A filter framework which allows you to define a filter
    	-- for a specific shape type. The types available include:
    	-- -   compound
    	-- -   compsolid
    	-- -   solid
    	-- -   shell
	-- -   face
    	-- -   wire
    	-- -   edge
    	-- -   vertex.

uses
    Shape from TopoDS,
    EntityOwner from SelectMgr,
    ShapeEnum from TopAbs
is

    Create (aType: ShapeEnum from TopAbs)
    returns mutable ShapeTypeFilter from StdSelect;
    	---Purpose: Constructs a filter object defined by the shape type aType.
    
    IsOk (me;anobj : EntityOwner from SelectMgr) 
    returns Boolean from Standard is redefined virtual;

    Type(me) returns ShapeEnum from TopAbs;
    	---Purpose: Returns the type of shape selected by the filter.
    	---C++: inline

    ActsOn(me; aStandardMode : ShapeEnum from TopAbs)
    returns Boolean from Standard is redefined virtual;

fields

    myType : ShapeEnum from TopAbs;

end ShapeTypeFilter;
