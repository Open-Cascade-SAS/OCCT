-- Created on: 1994-06-07
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SurfaceIterator from TopOpeBRepDS 
    inherits InterferenceIterator from TopOpeBRepDS

uses

    State               from TopAbs,
    Orientation         from TopAbs,
    ListOfInterference  from TopOpeBRepDS
    
is
    Create(L : ListOfInterference from TopOpeBRepDS) 
    returns SurfaceIterator;
    ---Purpose: Creates an  iterator on the  Surfaces on solid
    --          described by the interferences in <L>.
    
    Current(me) returns Integer from Standard
    ---Purpose: Index of the surface in the data structure.
    is static;
    
    Orientation(me; S : State from TopAbs) 
    returns Orientation from TopAbs
    is static;
    
end SurfaceIterator from TopOpeBRepDS;
