-- Created on: 1993-06-22
-- Created by: Martine LANGLOIS
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class MakeSurface from GeomToStep inherits Root from GeomToStep

    ---Purpose: This class implements the mapping between classes 
    --          Surface from Geom and the class Surface from StepGeom which
    --          describes a Surface from prostep. As Surface is an abstract
    --          Surface this class is an access to the sub-class required.
  
uses Surface from Geom,
     Surface from StepGeom
     
raises NotDone from StdFail
     
is 

Create ( C : Surface from Geom ) returns MakeSurface;

Value (me) returns Surface from StepGeom
    raises NotDone
    is static;
    ---C++: return const&

fields

    theSurface : Surface from StepGeom;
    	-- The solution from StepGeom
    	
end MakeSurface;



