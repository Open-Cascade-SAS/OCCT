-- Created on: 2002-01-04
-- Created by: data exchange team
-- Copyright (c) 2002-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1

class SeamEdge from StepShape
inherits OrientedEdge from StepShape

    ---Purpose: Representation of STEP entity SeamEdge

uses
    HAsciiString from TCollection,
    Vertex from StepShape,
    Edge from StepShape,
    Pcurve from StepGeom

is
    Create returns SeamEdge from StepShape;
	---Purpose: Empty constructor

    
		       
    Init (me: mutable; aRepresentationItem_Name: HAsciiString from TCollection;	       
                       aOrientedEdge_EdgeElement: Edge from StepShape;
                       aOrientedEdge_Orientation: Boolean;
                       aPcurveReference: Pcurve from StepGeom);
	---Purpose: Initialize all fields (own and inherited)

    PcurveReference (me) returns Pcurve from StepGeom;
	---Purpose: Returns field PcurveReference
    SetPcurveReference (me: mutable; PcurveReference: Pcurve from StepGeom);
	---Purpose: Set field PcurveReference

fields
    thePcurveReference: Pcurve from StepGeom;

end SeamEdge;
