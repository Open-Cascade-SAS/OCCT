-- File:	IGESSelect_FloatFormat.cdl
-- Created:	Wed Jun  1 16:04:47 1994
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1994


class FloatFormat  from IGESSelect    inherits FileModifier  from IGESSelect

    ---Purpose : This class gives control out format for floatting values :
    --           ZeroSuppress or no, Main Format, Format in Range (for values
    --           around 1.), as IGESWriter allows to manage it.
    --           Formats are given under C-printf form

uses CString, AsciiString from TCollection,
     IGESWriter , ContextWrite

is

    Create returns mutable FloatFormat;
    ---Purpose : Creates a new FloatFormat, with standard options :
    --           ZeroSuppress, Main Format = %E,
    --           Format between 0.001 and 1000. = %f

    SetDefault (me : mutable; digits : Integer = 0);
    ---Purpose : Sets FloatFormat to default value (see Create) but if <digits>
    --           is given positive, it commands Formats (main and range) to
    --           ensure <digits> significant digits to be displayed

    SetZeroSuppress (me : mutable; mode : Boolean);
    ---Purpose : Sets ZeroSuppress mode to a new value

    SetFormat (me : mutable; format : CString = "%E");
    ---Purpose : Sets Main Format to a new value
    --           Remark : SetFormat, SetZeroSuppress and SetFormatForRange are
    --           independant

    SetFormatForRange (me : mutable; format : CString = "%f";
    	    	       Rmin : Real = 0.1; Rmax : Real = 1000.0);
    ---Purpose : Sets Format for Range to a new value with its range of
    --           application.
    --           To cancel it, give format as "" (empty string)
    --           Remark that if the condition (0. < Rmin < Rmax)  is not
    --           verified, this secondary format will be ignored.
    --           Moreover, this secondary format is intended to be used in a
    --           range around 1.


    Format (me; zerosup  : out Boolean;
    	    	mainform : out AsciiString from TCollection;
		hasrange : out Boolean;
		forminrange : out AsciiString from TCollection;
		rangemin, rangemax : out Real);
    ---Purpose : Returns all recorded parameters :
    --           zerosup  : ZeroSuppress status
    --           mainform : Main Format (which applies out of the range, or
    --                       for every real if no range is set)
    --           hasrange : True if a FormatInRange is set, False else
    --                      (following parameters do not apply if it is False)
    --           forminrange : Secondary Format (it applies inside the range)
    --           rangemin, rangemax : the range in which the secondary format
    --                                applies


    Perform (me; ctx : in out ContextWrite;
    	     writer : in out IGESWriter);
    ---Purpose : Sets the Floatting Formats of IGESWriter to the recorded
    --           parameters

    Label (me) returns AsciiString from TCollection;
    ---Purpose : Returns specific Label : for instance,
    --           "Float Format [ZeroSuppress] %E [, in range R1-R2 %f]"

fields

    thezerosup   : Boolean;
    themainform  : AsciiString from TCollection;
    theformrange : AsciiString from TCollection;
    therangemin  : Real;
    therangemax  : Real;

end FloatFormat;

