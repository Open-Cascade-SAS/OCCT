-- Created on: 1994-06-17
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class FacetedBrepAndBrepWithVoids from StepShape 

inherits ManifoldSolidBrep from StepShape 


	--- This class is an implementation of EXPRESS
	--  ANDOR Subtype Declaration.
uses

	FacetedBrep from StepShape, 
	BrepWithVoids from StepShape, 
	ClosedShell from StepShape, 
	HArray1OfOrientedClosedShell from StepShape, 
	OrientedClosedShell from StepShape,
	HAsciiString from TCollection
is

	Create returns mutable FacetedBrepAndBrepWithVoids;
	---Purpose: Returns a FacetedBrepAndBrepWithVoids


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aOuter : mutable ClosedShell from StepShape) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aOuter : mutable ClosedShell from StepShape;
	      aFacetedBrep : mutable FacetedBrep from StepShape;
	      aBrepWithVoids : mutable BrepWithVoids from StepShape);

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aOuter : mutable ClosedShell from StepShape;
	      aVoids : mutable HArray1OfOrientedClosedShell from StepShape);

	-- Specific Methods for Field Data Access --

	SetFacetedBrep(me : mutable; aFacetedBrep : mutable FacetedBrep);
	FacetedBrep (me) returns mutable FacetedBrep;
	SetBrepWithVoids(me : mutable; aBrepWithVoids : mutable BrepWithVoids);
	BrepWithVoids (me) returns mutable BrepWithVoids;

	-- Specific Methods for ANDOR Field Data Access --

	SetVoids(me : mutable; aVoids : mutable HArray1OfOrientedClosedShell);
	Voids (me) returns mutable HArray1OfOrientedClosedShell;
	VoidsValue (me; num : Integer) returns mutable OrientedClosedShell;
	NbVoids (me) returns Integer;

	-- Specific Methods for ANDOR Field Data Access --


fields

	facetedBrep : FacetedBrep from StepShape;
	brepWithVoids : BrepWithVoids from StepShape;

end FacetedBrepAndBrepWithVoids;
