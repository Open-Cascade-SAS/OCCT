-- Created on: 1999-04-15
-- Created by: Denis PASCAL
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DocumentStorageDriver from MDocStd inherits StorageDriver from PCDM

	---Purpose: storage driver for  a standard document


uses Document           from TDocStd,
     Document           from PDocStd,
     SRelocationTable   from MDF,
     Document           from CDM, 
     MessageDriver      from CDM,       
     Document           from PCDM,
     ExtendedString from  TCollection,
     ASDriverTable from MDF


is


    Create
    returns  DocumentStorageDriver from MDocStd;
    
    CreateDocument (me: mutable) returns Document from PCDM
    ---Purpose: returns an empty PDocStd_Document. may be redefined;
    is virtual;
    	     
    Paste (me : mutable; TDOC   : Document from TDocStd;
                         PDOC   : Document from PDocStd;
			 aReloc : SRelocationTable from MDF);
  

    ---Purpose: virtual  methods of StorageDriver from PCDM
    --          ============================================
    
    Make (me: mutable; aDocument: Document from CDM)
    returns Document from PCDM 
    is redefined;
    
    ---Purpose: virtual methods (may be redefined by specialized application)
    --          =============================================================
    
    SchemaName(me) 
    returns   ExtendedString from  TCollection
    is virtual;
    
    AttributeDrivers(me : mutable; theMessageDriver : MessageDriver from CDM)
    returns ASDriverTable from MDF
    is virtual;
    
fields

    myDrivers : ASDriverTable from MDF;
    
end DocumentStorageDriver;
