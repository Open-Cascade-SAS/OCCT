-- Created on: 1997-03-03
-- Created by: Yves FRICAUD
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

private class Identifier from TNaming 

	---Purpose: 

uses

    Label            from TDF,
    Shape            from TopoDS,
    NamedShape       from TNaming,
    ListOfNamedShape from TNaming,
    ListOfShape      from TopTools,
    NameType         from TNaming,
    Localizer        from TNaming
is

    Create (Lab     : Label   from TDF;
    	    S	    : Shape   from TopoDS;
	    Context     : Shape   from TopoDS;
	    Geom        : Boolean from Standard)
    returns Identifier from TNaming;	    
    
    Create (Lab     : Label      from TDF;
    	    S	    : Shape      from TopoDS;
	    ContextNS   : NamedShape from TNaming;
	    Geom        : Boolean    from Standard)
    returns Identifier from TNaming;	    
    
    
    
    ---Category: Querying

    IsDone (me) returns Boolean from Standard;

    Type (me) returns NameType from TNaming;

    IsFeature (me : in out) returns Boolean from Standard;
  
    Feature   (me) returns NamedShape  from TNaming;
    
    
    InitArgs (me : in out);
    
    MoreArgs (me) returns Boolean from Standard;
    
    NextArg (me : in out);
    
    ArgIsFeature(me) returns Boolean from Standard;	
    
    FeatureArg (me : in out) returns NamedShape from TNaming;

    ShapeArg (me : in out) returns Shape from TopoDS;
    
    ShapeContext (me) returns Shape from TopoDS;

    NamedShapeOfGeneration  (me) returns NamedShape from TNaming;

    ---Category: Private methods.

    AncestorIdentification(me        : in out; 
    	    	    	   Localizer : in out Localizer from TNaming;
    	    	    	   Context   :        Shape     from TopoDS);
			   
    PrimitiveIdentification(me        : in out; 
    	    	    	    Localizer : in out Localizer  from TNaming;
    	    	    	    NS        :        NamedShape from TNaming);

    GeneratedIdentification(me        : in out; 
    	    	    	    Localizer : in out Localizer  from TNaming;
			    NS        :        NamedShape from TNaming);


    Identification(me        : in out; 
    	    	   Localizer : in out Localizer  from TNaming;	
    	    	   NS        :        NamedShape from TNaming);


    Init(me : in out; Context : Shape   from TopoDS) is private;
		  
fields
    
    myTDFAcces       : Label   from TDF;	
    myShape          : Shape   from TopoDS;
    
    myDone           : Boolean from Standard;

    myIsFeature      : Boolean          from Standard;
    myType           : NameType         from TNaming;
    myFeature        : NamedShape       from TNaming;
    myPrimitiveArgs  : ListOfNamedShape from TNaming;	
    myShapeArgs      : ListOfShape      from TopTools;
    myNSContext      : NamedShape       from TNaming;
    
end Identifier;


