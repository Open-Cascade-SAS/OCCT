-- Created on: 1994-10-03
-- Created by: Christian CAILLET
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class TransientListBinder  from Transfer  inherits Binder from Transfer

    ---Purpose : This binder binds several (a list of) Transients with a starting
    --           entity, when this entity itself corresponds to a simple list
    --           of Transients. Each part is not seen as a sub-result of an
    --           independant componant, but as an item of a built-in list

uses CString, Type,
	      HSequenceOfTransient from TColStd

raises TypeMismatch, OutOfRange

is

    Create returns mutable TransientListBinder;

    Create (list : mutable HSequenceOfTransient from TColStd)
    	 returns mutable TransientListBinder;

    IsMultiple (me) returns Boolean  is redefined;
    -- returns True if more than one result

    ResultType (me) returns Type;
    -- returns Standard_Transient

    ResultTypeName (me) returns CString;
    -- returns list(Standard_Transient)

    AddResult (me : mutable; res : Transient);
    ---Purpose : Adds an item to the result list

    Result (me) returns HSequenceOfTransient from TColStd;

    SetResult (me : mutable; num : Integer; res : Transient);
    ---Purpose : Changes an already defined sub-result

    NbTransients (me) returns Integer;

    Transient (me; num : Integer) returns Transient
    	raises OutOfRange;
    ---C++ : return const &


fields

    theres :  HSequenceOfTransient from TColStd;

end TransientListBinder;
