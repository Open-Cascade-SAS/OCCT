-- Created on: 1999-11-03
-- Created by: Denis PASCAL
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



private class Scope from TNaming 


    ---Purpose: this class manage a scope of labels
    --          ===================================


uses Label      from TDF,
     LabelMap   from TDF,
     NamedShape from TNaming,
     Shape      from TopoDS

is

    Create
    ---Purpose: WithValid = FALSE
    returns Scope from TNaming;

    Create (WithValid : Boolean from Standard)
    ---Purpose: if <WithValid> the scope is defined by the map. If not
    --          on the whole framework.
    returns Scope from TNaming;    

    Create (valid : in out LabelMap from TDF)
    ---Purpose: create a scope with a map. WithValid = TRUE.
    returns Scope from TNaming;

    WithValid (me)
    returns Boolean from Standard;  

    WithValid (me : in out; mode : Boolean from Standard);

    ClearValid (me :  in  out);

    Valid (me : in  out; L :Label from TDF);
    
    ValidChildren (me : in  out; L        : Label from TDF;
                                 withroot : Boolean from Standard = Standard_True);    

    Unvalid (me : in  out; L :Label from TDF);
    
    UnvalidChildren (me : in  out; L        : Label from TDF;
                                   withroot : Boolean from Standard = Standard_True);
    
    IsValid (me; L :Label from TDF) 
    returns Boolean  from  Standard; 
    
    GetValid (me)
    ---C++: return const &
    returns LabelMap from TDF;    

    ChangeValid (me : in out)
    ---C++: return &
    returns LabelMap from TDF;

    CurrentShape (me ; NS : NamedShape from TNaming)
    ---Purpose:  Returns  the current  value of  <NS> according to the
    --          Valid Scope.
    returns Shape from TopoDS;			    


fields
   
    myWithValid  : Boolean  from Standard;
    myValid      : LabelMap from TDF;

end Scope;
