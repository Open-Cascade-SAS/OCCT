-- Created on: 1998-06-03
-- Created by: data exchange team
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package ShapeUpgrade 

    	---Purpose:  This package provides tools
    	-- for splitting and converting shapes by some criteria. It
    	-- provides modifications of the kind when one topological
    	-- object can be converted or splitted to several ones. In
    	-- particular this package contains high level API classes which perform: 
    	--      converting geometry of shapes up to given continuity, 
    	--      splitting revolutions by U to segments less than given value, 
    	--      converting to beziers, 
    	--      splitting closed faces. 
    
uses
    gp,
    Geom,
    Geom2d,
    GeomAbs,
    Adaptor3d,
    GeomAdaptor,
    Geom2dAPI,
    TopLoc,
    TColStd,
    TColGeom,
    TColGeom2d,
    TCollection,
    TopoDS,
    TopTools,
    TopAbs,
    ShapeExtend,
    ShapeBuild,
    ShapeAnalysis,
    BRepBuilderAPI

is

    --- Instanciation of generic classes (tools)
    
    private class Tool;
    
    	class EdgeDivide;
	
	    class ClosedEdgeDivide;
	    
    	class WireDivide;
    
    	class FaceDivide;
    
    	    class ClosedFaceDivide;
	    class FaceDivideArea;
    
    class ShapeDivide;
    	class ShapeDivideArea;
    
    class ShapeDivideContinuity;    
    	---Purpose: API Tool for converting shapes with C0 geometry into C1 ones
    
    class ShapeDivideAngle;
    	---Purpose: API Class for splitting revolutions to segments less than 90

    class ShapeConvertToBezier;
    	---Purpose: API Class for convering curves to beziers.
	
    class ShapeDivideClosed;
    	---Purpose:
	
    class ShapeDivideClosedEdges;
    	---Purpose:
	
    class SplitCurve;
	class SplitCurve2d;
    	    class SplitCurve2dContinuity;
	    class ConvertCurve2dToBezier;
    	class SplitCurve3d;
    	    class SplitCurve3dContinuity;
	    class ConvertCurve3dToBezier;
	
    class SplitSurface;
    	class SplitSurfaceContinuity;
	class SplitSurfaceAngle;
	class ConvertSurfaceToBezierBasis;
	class SplitSurfaceArea;
	
    class ShellSewing;
    	---Purpose: Provides access to a sewing algorithms from BRepOffsetAPI
    class FixSmallCurves;
    ---Purpose:
    class FixSmallBezierCurves;
    ---Purpose:
    
    class RemoveLocations;
    ---Purpose: Removes all locations sub-shapes of specified shape
    
    class RemoveInternalWires;
    ---Purpose: Removes all internal wires having area less than specified min area
    
    class UnifySameDomain;
    ---Purpose: Unifies same domain faces and edges of specified shape
    
    C0BSplineToSequenceOfC1BSplineCurve (BS   : BSplineCurve from Geom;
    	    	    	    	         seqBS: out HSequenceOfBoundedCurve from TColGeom)
    returns Boolean;
				      
    C0BSplineToSequenceOfC1BSplineCurve (BS   : BSplineCurve from Geom2d;
    	    	    	    	         seqBS: out HSequenceOfBoundedCurve from TColGeom2d)
    returns Boolean;
    --- Purpose: Converts C0 B-Spline curve into sequence of C1 B-Spline curves.
    --           This method splits B-Spline at the knots with multiplicities
    --           equal to degree, i.e. unlike method
    --           GeomConvert::C0BSplineToArrayOfC1BSplineCurve this one does not
    --           use any tolerance and therefore does not change the geometry of
    --           B-Spline.
    --           Returns True if C0 B-Spline was successfully splitted, else
    --           returns False (if BS is C1 B-Spline).

end ShapeUpgrade;
