-- Created on: 1994-01-10
-- Created by: Yves FRICAUD
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class PointOnBis from Bisector 

	---Purpose: 
    
uses 
    Pnt2d from gp

is
    Create returns PointOnBis from Bisector;
    
    Create ( Param1, Param2, ParamBis, Distance : Real; Point : Pnt2d) 
    returns PointOnBis from Bisector; 
    
    ParamOnC1 (me : in out; Param : Real)
    is static;
    
    ParamOnC2 (me : in out; Param : Real)
    is static;
    
    ParamOnBis (me : in out; Param : Real)
    is static;
    
    Distance (me : in out; Distance : Real)
    is static;
    
    IsInfinite (me : in out; Infinite : Boolean)
    is static;

    Point (me : in out ; P :Pnt2d)
    is static;
    
    ParamOnC1 (me) returns Real
    is static;
    
    ParamOnC2 (me) returns Real
    is static;

    ParamOnBis (me) returns Real
    is static;
        
    Distance (me) returns Real
    is static;
    
    Point (me) returns Pnt2d
    is static;
    
    IsInfinite (me) returns Boolean 
    is static;
    
    Dump (me) is static;
    
fields

    param1   : Real;
    param2   : Real;
    paramBis : Real;
    distance : Real;
    infinite : Boolean;	
    point    : Pnt2d from gp;
    
end PointOnBis;
