-- Created by: CAL
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Vertex from Graphic2d

	---Version:

	---Purpose: This class allows the creation and update of a
	--	    2D point.

	---Keywords: Vertex, Coordinate, Point
	---Warning:
	---References:

uses
	Drawer	from Graphic2d,
	Length	from Quantity

is
	-------------------------
	-- Category: Constructors
	-------------------------

	Create
	returns Vertex from Graphic2d;
	---Level: Public
	---Purpose: Creates a point with 0.0, 0.0 coordinates.

	Create (AX, AY: Real from Standard)
	returns Vertex from Graphic2d;
	---Level: Public
	---Purpose: Creates a point with <AX>, <AY> coordinates.

	Create (AX, AY: ShortReal from Standard)
	returns Vertex from Graphic2d;
	---Level: Public
	---Purpose: Creates a point with <AX>, <AY> coordinates.

	---------------------------------------------------
	-- Category: Methods to modify the class definition
	---------------------------------------------------

	SetCoord (me: in out;
		  Xnew, Ynew: Length from Quantity)
	is static;
	---Level: Public
	---Purpose: Modifies the coordinates of the point <me>.
	---Category: Methods to modify the class definition

	SetXCoord (me: in out;
		   Xnew: Length from Quantity)
	is static;
	---Level: Public
	---Purpose: Modifies the X coordinate of the point <me>.
	---Category: Methods to modify the class definition

	SetYCoord (me: in out;
		   Ynew: Length from Quantity)
	is static;
	---Level: Public
	---Purpose: Modifies the Y coordinate of the point <me>.
	---Category: Methods to modify the class definition

	----------------------------
	-- Category: Inquire methods
	----------------------------

	Coord (me;
		AX, AY: out Length from Quantity)
	is static;
	---Level: Public
	---Purpose: Returns the coordinates of the point <me>.
	---Category: Inquire methods

	X (me) returns Length from Quantity
	is static;
	---Level: Public
	---Purpose: Returns the X coordinates of the point <me>.
	---Category: Inquire methods

	Y (me) returns Length from Quantity
	is static;
	---Level: Public
	---Purpose: Returns the Y coordinate of the point <me>.
	---Category: Inquire methods

   	IsEqual (me ; other : Vertex) returns Boolean
   	is static;
   	---Level: Public
   	---Purpose: Test if <me> and <other> are the the same vertex.
   	---C++: alias operator ==

	--------------------------
	-- Category: Class methods
	--------------------------

	Distance (myclass;
		   AV1, AV2: Vertex from Graphic2d)
	returns Length from Quantity;
	---Level: Public
	---Purpose: Returns the distance between <AV1> and <AV2>.
	---Category: Class methods

fields
	myX:	ShortReal from Standard;
	myY:	ShortReal from Standard;

end Vertex from Graphic2d;
