-- Created on: 1991-04-04
-- Created by: Remi GILET
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


package GccIter

    ---Purpose :
    --           This package provides an implementation of analytics 
    --           algorithms (using only non persistant entities) used 
    --           to create 2d lines or circles with geometric constraints.
    --
    -- Exceptions :
    -- 	            IsParallel which inherits DomainError. This exception 
    -- 	            is raised in the class Lin2dTanObl when we want to 
    -- 	            find the intersection point between the solution and 
    -- 	            the second argument with a null angle.

uses GccEnt,
     GccInt,
     GccAna,
     StdFail,
     gp,
     math

is

enumeration Type1 is CuCuCu,CiCuCu,CiCiCu,CiLiCu,LiLiCu,LiCuCu;

enumeration Type2 is CuCuOnCu,CiCuOnCu,LiCuOnCu,CuPtOnCu,
                     CuCuOnLi,CiCuOnLi,LiCuOnLi,CuPtOnLi,
		     CuCuOnCi,CiCuOnCi,LiCuOnCi,CuPtOnCi;

enumeration Type3 is CuCu,CiCu;

generic class FunctionTanCuCu;

generic class FunctionTanCirCu;

generic class FunctionTanCuCuCu;

generic class FunctionTanCuCuOnCu;

generic class FunctionTanCuPnt;

generic class FunctionTanObl;

generic class Lin2dTanObl, FuncTObl;
    -- Create a 2d line TANgent to a 2d curve and OBLic to a 2d line.

generic class Lin2d2Tan, FuncTCuCu, FuncTCirCu, FuncTCuPt;
    -- Create a 2d line TANgent to 2 2d entities.

generic class Circ2d3Tan, FuncTCuCuCu;
    -- Create a 2d circle TANgent to 3 2d entities.

generic class Circ2d2TanOn, FuncTCuCuOnCu;
    -- Create a 2d circle TANgent to a 2d entity and centered ON a 2d 
    -- entity (not a point).

exception IsParallel inherits DomainError from Standard;

end GccIter;
