-- Created on: 1993-09-29
-- Created by: Isabelle GRIGNON
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class GeomTool from BRepMesh
       	---Purpose: 

uses 
     Pnt                  from gp,
     Vec                  from gp,
     Dir                  from gp,
     Pnt2d                from gp,
     IsoType              from GeomAbs,
     TangentialDeflection from GCPnts,
     Curve                from BRepAdaptor,
     HSurface             from BRepAdaptor
     


is

    Create (C : in out Curve from BRepAdaptor;
            Ufirst,Ulast,AngDefl, Deflection : Real;
            nbpointsmin: Integer = 2)
    	returns GeomTool;
    
    Create (S        : HSurface from BRepAdaptor;
            ParamIso : Real;
            Type     : IsoType  from GeomAbs;
    	    Ufirst,Ulast,AngDefl,Deflection : Real;
    	    nbpointsmin: Integer = 2) returns GeomTool;

    AddPoint(me : in out; thePnt : in Pnt from gp;
                          theParam : in Real;
                          theIsReplace : in Boolean = Standard_True)
    returns Integer from Standard;
    ---Purpose: Add point to already calculated points (or replace existing)
    --          Returns index of new added point
    --           or founded with parametric tolerance (replaced if theIsReplace is true)
	    
    NbPoints(me) returns Integer from Standard;
    
    Value(me; IsoParam : Real ; Index : Integer ; 
          W : out Real; P : out Pnt from gp; UV : out Pnt2d from gp);
	      
    Value(me;C : Curve from BRepAdaptor;
             S : HSurface from BRepAdaptor;
             Index : Integer from Standard; 
    	     W : out Real; P : out Pnt from gp; UV : out Pnt2d from gp);    
	
    D0(myclass; F : HSurface  from BRepAdaptor;U,V : Real; P : out Pnt);
	
    Normal(myclass; F : HSurface from BRepAdaptor;U,V : Real ; P : out Pnt from gp; 
    	    	    	    	    	   Nor : out  Dir from gp)
    returns Boolean from Standard;
    ---Purpose: return false if the normal can not be computed 

fields

pnts                : TangentialDeflection from GCPnts;
parametric          : IsoType           from GeomAbs;

end GeomTool;
