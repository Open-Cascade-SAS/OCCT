-- Created on: 1993-09-29
-- Created by: Denis PASCAL
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class RGNode from GraphTools

uses SC                from GraphTools,
     SequenceOfInteger from TColStd

is

    Create returns RGNode;
    
    Reset (me : in out);
    
    SetVisited (me : in out; v : Integer from Standard);
    
    GetVisited (me) 
    returns Integer from Standard;
    
    AddAdj (me : in out; adj : Integer from Standard);
    
    NbAdj (me) 
    returns Integer from Standard;
    
    GetAdj (me; index : Integer from Standard)
    returns Integer from Standard;

    SetSC (me : in out; SC : SC from GraphTools);

    GetSC (me) 
    returns SC from GraphTools;

fields

    visited : Integer from Standard;
    myAdj   : SequenceOfInteger from TColStd;
    mySC    : SC from GraphTools;

end RGNode;      	

