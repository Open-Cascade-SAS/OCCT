-- Created on: 1998-08-27
-- Created by: Robert COUBLANC
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class EventManager from ViewerTest inherits TShared from MMgt

	---Purpose: used to manage mouse event (move,select,shiftselect)
  --          By default the events are transmitted to interactive context.


uses
    View                from V3d,
    InteractiveContext  from AIS,
    Array1OfPnt2d       from TColgp
is

    Create (aView: View from V3d;
            aCtx :InteractiveContext from AIS)
    returns EventManager from ViewerTest;
    
    MoveTo (me:mutable;
            xpix, ypix  : Integer from Standard) is virtual;
    
    Select(me:mutable) is virtual;
    
    ShiftSelect(me:mutable) is virtual;

    Select(me:mutable;xmin,ymin,xmax,ymax:Integer) is virtual;
    
    ShiftSelect(me:mutable;xmin,ymin,xmax,ymax:Integer) is virtual;
    
    Select(me:mutable;thePolyline:Array1OfPnt2d from TColgp) is virtual;
    
    ShiftSelect(me:mutable;thePolyline:Array1OfPnt2d from TColgp) is virtual;

    Context(me) returns InteractiveContext from AIS;
    ---C++: inline
    ---C++: return const&

fields

    myCtx : InteractiveContext  from AIS;
    myView: View                from V3d;
    myX   : Integer             from Standard;
    myY   : Integer             from Standard;
    
end EventManager;
