-- Created on: 1995-12-06
-- Created by: Frederic MAUPAS
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DirectionCountSelect from StepVisual

    -- a Select Type (hand generated)

uses

    Integer from Standard
    
is

    Create returns DirectionCountSelect;
    
    SetTypeOfContent(me : in out; aTypeOfContent : Integer);

    TypeOfContent(me) returns Integer;
	--        1 -> UDirectionCount
	--        2 -> VDirectionCount

    UDirectionCount(me) returns Integer from Standard;
    
    SetUDirectionCount(me : in out; aUDirectionCount : Integer from Standard);
    
    VDirectionCount(me) returns Integer from Standard;
    
    SetVDirectionCount(me : in out; aUDirectionCount : Integer from Standard);


fields

    theUDirectionCount : Integer from Standard;
    theVDirectionCount : Integer from Standard;
    theTypeOfContent   : Integer from Standard;

end DirectionCountSelect;
