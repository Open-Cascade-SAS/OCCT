-- Created on: 2012-08-06
-- Created by: jgv@ROLEX
-- Copyright (c) 2012-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MiddlePath from BRepOffsetAPI inherits MakeShape from BRepBuilderAPI

    	---Purpose: Describes functions to build a middle path of a
    	--          pipe-like shape

uses

    Shape from TopoDS,
    Wire  from TopoDS,
    Edge  from TopoDS,
    Face  from TopoDS,
    MapOfShape from TopTools,
    SequenceOfSequenceOfShape from BRepOffsetAPI
    
is
    --Create(aShape    : Shape from TopoDS;
    	--   StartWire : Wire from TopoDS)
    --returns MiddlePath from BRepOffsetAPI;
    
    --Create(aShape    : Shape from TopoDS;
    	--   StartEdge : Edge from TopoDS)
    --returns MiddlePath from BRepOffsetAPI;
    
    Create(aShape     : Shape from TopoDS;
    	   StartShape : Shape from TopoDS;
	   EndShape   : Shape from TopoDS)
    ---Purpose: General constructor.
    --          StartShape and EndShape may be
    --          a wire or a face
    returns MiddlePath from BRepOffsetAPI;

    Build(me: in out)
    is redefined;

fields
    
    myInitialShape : Shape from TopoDS;
    myStartWire    : Wire  from TopoDS;
    myEndWire      : Wire  from TopoDS;
    myClosedSection  : Boolean from Standard;
    myClosedRing     : Boolean from Standard;
    
    myStartWireEdges : MapOfShape from TopTools;
    myEndWireEdges   : MapOfShape from TopTools;
    
    myPaths        : SequenceOfSequenceOfShape from BRepOffsetAPI;
    
end MiddlePath;
