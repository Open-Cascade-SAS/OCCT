-- Created on: 1991-03-05
-- Created by: Philippe DAUTRY
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package GccAna 

    ---Purpose : This package provides an implementation of analytics 
    --         algorithms (using only non persistant entities) used 
    --         to create 2d lines or circles with geometric constraints.

uses Standard,
     StdFail,
     gp,
     TColStd,
     TColgp,
     GccInt,
     GccEnt
     

is

    -- Exceptions :

exception NoSolution inherits Failure from Standard;

class Lin2dTanPar;

class Lin2dTanPer;

class Lin2dTanObl;

class Lin2d2Tan;

class Lin2dBisec;

class Circ2dTanCen;

class Circ2d3Tan;

class Circ2d2TanRad;

class Circ2d2TanOn;

class Circ2dTanOnRad;

class Pnt2dBisec;

class Circ2dBisec;

class CircLin2dBisec;

class CircPnt2dBisec;

class LinPnt2dBisec;

end GccAna;
