-- Created on: 1997-03-05
-- Created by: Joelle CHAUVET
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class PlateG0Criterion from GeomPlate inherits Criterion from AdvApp2Var


uses
    SequenceOfXY,SequenceOfXYZ from TColgp,
    Patch,Context from AdvApp2Var,
    CriterionType,CriterionRepartition from AdvApp2Var


is

    Create( Data : SequenceOfXY;
    	    G0Data : SequenceOfXYZ;
            Maximum : Real;
    	    Type : CriterionType  = AdvApp2Var_Absolute;
    	    Repart : CriterionRepartition  = AdvApp2Var_Regular)  returns PlateG0Criterion;
	    
    Value(me; P : in out Patch; C : Context )
    is redefined;
    
    IsSatisfied(me; P : Patch ) returns Boolean
    is redefined;
    

    
fields
    myData : SequenceOfXY;
    myXYZ : SequenceOfXYZ;
    
end PlateG0Criterion;

