-- Created on: 2000-12-25
-- Created by: Igor FEOKTISTOV <ifv@nnov.matra-dtv.fr>
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

class Intersection from QANewModTopOpe inherits BooleanOperation from BRepAlgoAPI 

---Purpose: provides  intersection  of  two  shapes;
 
uses

    Shape from TopoDS, 
    DataMapOfShapeListOfShape from TopTools,
    ListOfShape from TopTools
     
is 
  
    Create(theObject1,  theObject2 : Shape from TopoDS )
    ---Purpose: 
    
    returns Intersection  from QANewModTopOpe;   

    Generated (me: in out; theS : Shape from TopoDS)
    	---Purpose: Returns the list  of shapes generated from the shape <S>. 
        ---C++: return const & 
        ---Level: Public
    returns ListOfShape from TopTools
    is redefined; 

    HasGenerated (me)
    	returns Boolean from Standard
	is redefined;
    	---Purpose: Returns true if there is at least one generated shape.
    	---         For use in BRepNaming.

    IsDeleted (me: in out;  
    	    aS : Shape from TopoDS)
    	returns Boolean
    	is redefined;


    HasDeleted (me)
    	returns Boolean from Standard
	is redefined;
    	---Purpose: Returns true if there is at least one deleted shape.
    	---         For use in BRepNaming.

fields
    
    myMapGener: DataMapOfShapeListOfShape from TopTools;

end  Intersection;
