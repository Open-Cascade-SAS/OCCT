-- Created on: 1994-06-16
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ReadWriteModule from RWHeaderSection  inherits ReadWriteModule from StepData

	---Purpose : General module to read and write HeaderSection entities

uses Transient,
     SequenceOfAsciiString    from TColStd,
     AsciiString              from TCollection,
     Check                    from Interface,
     StepReaderData           from StepData,
     StepWriter               from StepData

is

	Create returns mutable ReadWriteModule from RWHeaderSection;

	CaseStep (me; atype : AsciiString from TCollection) returns Integer;
	---Purpose : associates a positive Case Number to each type of HeaderSection entity,
	-- given as a String defined in the EXPRESS form

	CaseStep(me; types : SequenceOfAsciiString from TColStd) returns Integer is redefined;
	---Purpose : associates a positive Case Number to each type of HeaderSection Complex entity,
	-- given as a String defined in the EXPRESS form

	IsComplex (me; CN : Integer) returns Boolean is redefined;
	---Purpose : returns True if the Case Number corresponds to a Complex Type

	StepType (me; CN : Integer) returns AsciiString from TCollection;
	---Purpose : returns a StepType (defined in EXPRESS form which belongs to a 
	-- Type of Entity, identified by its CaseNumber determined by Protocol
	---C++ : return const &

	ReadStep (me; CN : Integer; data : StepReaderData; num : Integer;
	            ach : in out Check; ent : mutable Transient);

	WriteStep (me; CN : Integer; SW : in out StepWriter; ent : Transient);

end ReadWriteModule;
