-- File:	Select2D_SensitiveSegment.cdl
-- Created:	Thu Jan 26 11:45:23 1995
-- Author:	Mister rmi
--		<rmi@photon>
---Copyright:	 Matra Datavision 1995


class SensitiveSegment from Select2D 
inherits SensitiveEntity from Select2D


	---Purpose: A framework to define sensitive areas along a line segment.

uses
    Pnt2d from gp,
    EntityOwner from SelectBasics,
    ListOfBox2d from SelectBasics    

is


    Create (OwnerId      : EntityOwner from SelectBasics;
    	    FirstP,LastP : Pnt2d from gp;
    	    MaxRect      : Integer = 3)
     returns mutable SensitiveSegment;
    	---Purpose: Constructs the sensitive line segment object defined
    	-- by the owner OwnerId, the 2D starting and ending
    	-- points FirstPoint and LastPoint and the maximum
    	-- number of sensitive bounding boxes MaxRect.
    	-- The parameters can be modified using the functions provided.	    
	    
    Set (me:mutable; MaxRect : Integer) is static;
    	---Purpose: Sets the maximum number of 2D sensitive bounding boxes - MaxRect.
    
    
    
    StartPoint (me : mutable ; aPt : Pnt2d from gp) is static;
    	---Level: Public 
    	---C++: inline
    	---Purpose: changes the start Point of the Segment;
    


    EndPoint (me : mutable ; aPt : Pnt2d from gp) is static;
    	---Level: Public 
    	---C++: inline
    	---Purpose: changes the end point of the segment
    
    
    StartPoint (me) returns Pnt2d from gp;
    	---Level: Public 
    	---Purpose: gives the 3D start Point of the Segment
    	---C++: return const&
    	---C++: inline
    
    
    EndPoint(me) returns Pnt2d from gp;
    	---Level: Public 
    	---Purpose: Returnes the 3D start Point of the Segment
    	---C++: return const&
    	---C++: inline
    
    
    Areas   (me:mutable;aSeq : in out ListOfBox2d from SelectBasics) is static;
    
    
    Matches (me   : mutable; 
    	     X,Y  : Real from Standard;
    	     aTol : Real from Standard;
    	     DMin : out Real from Standard)
    returns Boolean is static;

    Matches (me  :mutable; 
             XMin,YMin,XMax,YMax : Real from Standard;
             aTol: Real from Standard) 
    returns Boolean
    is static;
    

    MaxBoxes(me) returns Integer is redefined static;
    	---Level: Public 
    	---Purpose: Returns the max number of sensitive aeas describing the sensitive segment
    	---C++: inline

fields

    mymaxrect : Integer;
    mystart   : Pnt2d from gp;
    myend     : Pnt2d from gp;

end SensitiveSegment;
