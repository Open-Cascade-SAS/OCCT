-- Created by: Peter KURNEV
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ShapeInfo from BOPDS 

	---Purpose: 
    	-- The class BOPDS_ShapeInfo is to store  
    	-- handy information about shape
uses 
    Box   from Bnd, 
    Shape from TopoDS, 
    BaseAllocator from BOPCol, 
    ListOfInteger from BOPCol, 
    ShapeEnum from TopAbs 
	
--raises

is
    Create 
    	returns ShapeInfo from BOPDS;  
    ---C++: alias "virtual ~BOPDS_ShapeInfo();" 
    ---C++: inline 
     	---Purpose:  
    	--- Empty contructor  
    	---    
    Create (theAllocator: BaseAllocator from BOPCol) 
    	returns ShapeInfo from BOPDS;
    ---C++: inline 
    	---Purpose:   
     	---  Contructor    
    	---  theAllocator - the allocator to manage the memory     
    	---   
    SetShape(me:out; 
    	    theS: Shape from TopoDS); 
    ---C++: inline  
    	---Purpose: 
    	--- Modifier   
	--- Sets the shape <theS>
    Shape(me) 
       returns Shape from TopoDS; 
    ---C++: return const &       
    ---C++: inline 
     	---Purpose: 
	--- Selector 
	--- Returns the shape    
     
    SetShapeType(me:out; 
    	    theType: ShapeEnum from TopAbs); 
    ---C++: inline  
      	---Purpose: 
    	--- Modifier   
	--- Sets the type of shape theType 
	
    ShapeType(me) 
    	returns ShapeEnum from TopAbs; 
    ---C++: inline  
    	---Purpose: 
	--- Selector 
        --- Returns the type of shape   
     
    SetBox(me:out; 
    	    theBox:Box from Bnd); 
    ---C++: inline 
    	---Purpose:      
     	--- Modifier   
	--- Sets the boundung box of the shape theBox
	
	
    Box(me) 
    	returns Box from Bnd; 
    ---C++: return const &    
    ---C++: inline 
    	---Purpose: 
	--- Selector 
        --- Returns the boundung box of the shape  
     
    ChangeBox(me:out) 
    	returns Box from Bnd; 
    ---C++: return  &    
    ---C++: inline   
    	---Purpose: 
	--- Selector/Modifier 
        --- Returns the boundung box of the shape 
    
    SubShapes(me) 
    	returns ListOfInteger from BOPCol;  
    ---C++: return const & 
    ---C++: inline 
    	---Purpose: 
	--- Selector 
        --- Returns the list of indices of sub-shapes 

    ChangeSubShapes(me:out) 
    	returns ListOfInteger from BOPCol;  
    ---C++: return & 
    ---C++: inline 
    	---Purpose: 
	--- Selector/ Modifier
        --- Returns the list of indices of sub-shapes 
  
    HasSubShape(me; 
    	    theI:Integer from Standard) 
	returns Boolean from Standard;   
    ---C++: inline  
        ---Purpose: 
	--- Query
        --- Returns true if the shape has sub-shape with 
        --- index theI 
	 
    HasReference(me) 
     	returns Boolean from Standard;  
    ---C++: inline  
     	--- Query
        --- Returns true if the shape has a reference information 

    SetReference(me:out; 
     	   theI: Integer from Standard); 
    ---C++: inline    
	---Purpose:      
     	--- Modifier   
	--- Sets the index of a reference information 
	 
    Reference(me) 
     	returns Integer from Standard; 	     
    ---C++: inline   
     	---Purpose:      
     	--- Selector   
	--- Returns the index of a reference information 
     
    HasBRep(me) 
	returns Boolean from Standard;   
    ---C++: inline 
    	---Purpose: 
	--- Query
        --- Returns true if the shape has boundary representation    
     
    IsInterfering(me) 
	returns Boolean from Standard;   
    ---C++: inline 
    	---Purpose: 
        --- Returns true if the shape can be participant of  
        --- an interference 	  
    -- 
    ---  Flag 
    --  
    HasFlag(me) 
	returns Boolean from Standard;   
    ---C++: inline  
    	---Purpose: 
    	--- Query
        --- Returns true if there is flag.  
     
    HasFlag(me; 
    	    theFlag:out Integer from Standard) 
	returns Boolean from Standard;   
    ---C++: inline  
    	---Purpose: 
    	--- Query
        --- Returns true if there is flag.  
    	--- Returns the the  flag theFlag  
      
    SetFlag(me:out; 
    	    theI:Integer from Standard); 
    ---C++: inline  
    	---Purpose:      
     	--- Modifier   
	--- Sets the flag 
    Flag(me) 
     	returns Integer from Standard; 	     
    ---C++: inline 
     	---Purpose:  
    	--- Returns the flag  

    Dump(me); 

fields
    myShape    : Shape from TopoDS is protected; 
    myType     : ShapeEnum from TopAbs is protected;         
    myBox      : Box from Bnd is protected; 
    mySubShapes: ListOfInteger from BOPCol is protected; 
    myReference: Integer from Standard is protected; 
    myFlag     : Integer from Standard is protected;  
    
end ShapeInfo;
