-- Created on: 2008-05-30
-- Created by: Vladislav ROMASHKO
-- Copyright (c) 2008-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class FastConverter from Voxel

    ---Purpose: Converts a shape to voxel representation.
    --          It does it fast, but with less precision.
    --          Also, it doesn't fill-in volumic part of the shape.

uses

    Pnt     from gp,
    Pln     from gp,
    Shape   from TopoDS,
    BoolDS  from Voxel,
    ColorDS from Voxel,
    ROctBoolDS from Voxel

is

    Create(shape  :     Shape   from TopoDS;
    	   voxels : out BoolDS  from Voxel;
    	   deflection : Real    from Standard = 0.1;
	   nbx    :     Integer from Standard = 10;
    	   nby    :     Integer from Standard = 10;
    	   nbz    :     Integer from Standard = 10;
    	   nbthreads :  Integer from Standard = 1;
    	   useExistingTriangulation : Boolean from Standard = Standard_False)
    ---Purpose: A constructor for conversion of a shape into a cube of boolean voxels.
    --          It allocates the voxels in memory.
    --          "nbthreads" defines the number of threads used to convert the shape.
    returns FastConverter from Voxel;

    Create(shape  :     Shape   from TopoDS;
    	   voxels : out ColorDS from Voxel;
    	   deflection : Real    from Standard = 0.1;
	   nbx    :     Integer from Standard = 10;
    	   nby    :     Integer from Standard = 10;
    	   nbz    :     Integer from Standard = 10;
    	   nbthreads :  Integer from Standard = 1;
    	   useExistingTriangulation : Boolean from Standard = Standard_False)
    ---Purpose: A constructor for conversion of a shape into a cube of colored voxels.
    --          It allocates the voxels in memory.
    --          "nbthreads" defines the number of threads used to convert the shape.
    returns FastConverter from Voxel;

    Create(shape  :     Shape   from TopoDS;
    	   voxels : out ROctBoolDS from Voxel;
    	   deflection : Real    from Standard = 0.1;
	   nbx    :     Integer from Standard = 10;
    	   nby    :     Integer from Standard = 10;
    	   nbz    :     Integer from Standard = 10;
    	   nbthreads :  Integer from Standard = 1;
    	   useExistingTriangulation : Boolean from Standard = Standard_False)
    ---Purpose: A constructor for conversion of a shape into a cube of boolean voxels
    --          split into 8 sub-voxels recursively.
    --          It allocates the voxels in memory.
    --          "nbthreads" defines the number of threads used to convert the shape.
    returns FastConverter from Voxel;

    Convert(me : in out;
    	    progress : out Integer from Standard;
    	    ithread : Integer from Standard = 1)
    ---Purpose: Converts a shape into a voxel representation.
    --          It sets to 0 the outside volume of the shape and
    --          1 for surfacic part of the shape.
    --          "ithread" is the index of the thread for current call of ::Convert().
    --          Start numeration of "ithread" with 1, please.
    returns Boolean from Standard;
	
    ConvertUsingSAT(me : in out;
		    progress : out Integer from Standard;
    	    	    ithread : Integer from Standard = 1)
    ---Purpose: Converts a shape into a voxel representation using separating axis theorem.
    --          It sets to 0 the outside volume of the shape and
    --          1 for surfacic part of the shape.
    --          "ithread" is the index of the thread for current call of ::Convert().
    --          Start numeration of "ithread" with 1, please.
    returns Boolean from Standard;

    FillInVolume(me : in out;
    	    	 inner : Byte from Standard;
    	    	 ithread : Integer from Standard = 1)
    ---Purpose: Fills-in volume of the shape by a value.
    returns Boolean from Standard;
    
    FillInVolume(me : in out;
                 inner : Byte from Standard;
                 shape : Shape   from TopoDS;
                 ithread : Integer from Standard = 1)
    ---Purpose: Fills-in volume of the shape by a value.
    --          Uses the topological information from the provided shape
    --          to judge whether points are inside the shape or not
    --          (only when processing vertical faces).
    --          The inner value has to be positive.
    returns Boolean from Standard;


    ---Category: Private area
    --           ============

    Destroy(me : in out);
    ---C++: alias ~
    ---Purpose: A destructor.

    Init(me : in out)
    is private;

    GetBndBox(me;
    	      p1   : Pnt      from gp;
    	      p2   : Pnt      from gp;
    	      p3   : Pnt      from gp;
	      xmin : out Real from Standard;
	      ymin : out Real from Standard;
	      zmin : out Real from Standard;
	      xmax : out Real from Standard;
	      ymax : out Real from Standard;
	      zmax : out Real from Standard)
    is private;

    ComputeVoxelsNearTriangle(me;
    	    	       	      plane :     Pln           from gp;
			      p1    :     Pnt           from gp;
			      p2    :     Pnt           from gp;
			      p3    :     Pnt           from gp;
		       	      hdiag :     Real          from Standard;
		       	      ixmin :     Integer       from Standard;
		       	      iymin :     Integer       from Standard;
		       	      izmin :     Integer       from Standard;
		       	      ixmax :     Integer       from Standard;
		       	      iymax :     Integer       from Standard;
		              izmax :     Integer       from Standard)
    is private;

	ComputeVoxelsNearTriangle(me;

			      p1    :     Pnt           from gp;
			      p2    :     Pnt           from gp;
			      p3    :     Pnt           from gp;
  			      extents    :     Pnt           from gp;
  			      extents2    :     Pnt           from gp;
  			      extents4    :     Pnt           from gp;
		       	      ixmin :     Integer       from Standard;
		       	      iymin :     Integer       from Standard;
		       	      izmin :     Integer       from Standard;
		       	      ixmax :     Integer       from Standard;
		       	      iymax :     Integer       from Standard;
		              izmax :     Integer       from Standard)
    is private;

fields

    myShape       : Shape   from TopoDS;
    myVoxels      : Address from Standard;
    myDeflection  : Real    from Standard;
    myIsBool      : Integer from Standard; -- 0 - ColorDS, 1 - BoolDS, 2 - ROctBoolDS
    myNbX         : Integer from Standard;
    myNbY         : Integer from Standard;
    myNbZ         : Integer from Standard;
    myNbThreads   : Integer from Standard;
    myNbTriangles : Integer from Standard;
    myUseExistingTriangulation : Boolean from Standard;

end FastConverter;
