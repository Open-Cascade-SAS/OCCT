-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package StepFEA


uses
    TCollection,
    TColStd,
    StepData,
    StepBasic,
    StepGeom,
    StepRepr,
    StepElement

is 

    enumeration ElementVolume is 
	Volume
    end;

    enumeration CurveEdge is 
	ElementEdge
    end;

    enumeration CoordinateSystemType is 
	Cartesian,
	Cylindrical,
	Spherical
    end;
    
    enumeration EnumeratedDegreeOfFreedom is 
	XTranslation,
	YTranslation,
	ZTranslation,
	XRotation,
	YRotation,
	ZRotation,
	Warp
    end;

    enumeration UnspecifiedValue is 
	Unspecified
    end;
    
    class AlignedCurve3dElementCoordinateSystem;
    class ArbitraryVolume3dElementCoordinateSystem;
    class Curve3dElementProperty;
    class Curve3dElementRepresentation;
    class CurveElementEndCoordinateSystem;
    class CurveElementEndOffset;
    class CurveElementEndRelease;
    class CurveElementInterval;
      class CurveElementIntervalConstant;
      class CurveElementIntervalLinearlyVarying; -- added 23.01.2003
    class CurveElementLocation;
    class DummyNode;
    class ElementGeometricRelationship;
    class ElementGroup;
    class ElementRepresentation;
    class FeaAreaDensity;
    class FeaAxis2Placement3d;
    class FeaGroup;
    class FeaLinearElasticity;
    class FeaMassDensity;
    class FeaMaterialPropertyRepresentation;
    class FeaMaterialPropertyRepresentationItem;
    class FeaModel;
    class FeaModel3d;
    class FeaMoistureAbsorption;
    class FeaParametricPoint;
    class FeaRepresentationItem;
    class FeaSecantCoefficientOfLinearThermalExpansion;
    class FeaShellBendingStiffness;
    class FeaShellMembraneBendingCouplingStiffness;
    class FeaShellMembraneStiffness;
    class FeaShellShearStiffness;
    class FeaTangentialCoefficientOfLinearThermalExpansion;
    class GeometricNode;
    class Node;
    class NodeGroup;
    class NodeRepresentation;
    class NodeSet;
    class NodeWithSolutionCoordinateSystem;
    class NodeWithVector;
    class ParametricCurve3dElementCoordinateDirection;
    class ParametricCurve3dElementCoordinateSystem;
    class ParametricSurface3dElementCoordinateSystem;
    class Surface3dElementRepresentation;
    class SymmetricTensor22d;
    class SymmetricTensor23d;
    	class SymmetricTensor23dMember;
    class SymmetricTensor42d;
    class SymmetricTensor43d;
    	class SymmetricTensor43dMember;
    class Volume3dElementRepresentation;
    class FeaModelDefinition;
    class DegreeOfFreedom;
    	class DegreeOfFreedomMember;
    class FreedomsList;
    class FreedomAndCoefficient;
    class NodeDefinition;
    class AlignedSurface3dElementCoordinateSystem;
    class ConstantSurface3dElementCoordinateSystem;
    class FeaCurveSectionGeometricRelationship;   -- added 23.01.2003
    class FeaSurfaceSectionGeometricRelationship; -- added 23.01.2003
    class ElementOrElementGroup;  -- added 04.02.2003
    
   
imported Array1OfNodeRepresentation;
imported transient class HArray1OfNodeRepresentation;

imported Array1OfCurveElementInterval;
imported transient class HArray1OfCurveElementInterval;

imported Array1OfCurveElementEndOffset;
imported transient class HArray1OfCurveElementEndOffset;

imported Array1OfCurveElementEndRelease;
imported transient class HArray1OfCurveElementEndRelease;

imported Array1OfElementRepresentation;
imported transient class HArray1OfElementRepresentation;

imported Array1OfDegreeOfFreedom;
imported transient class HArray1OfDegreeOfFreedom;

imported SequenceOfElementRepresentation;
imported transient class HSequenceOfElementRepresentation;

imported SequenceOfElementGeometricRelationship;
imported transient class HSequenceOfElementGeometricRelationship;

imported SequenceOfNodeRepresentation;
imported transient class HSequenceOfNodeRepresentation;

imported SequenceOfCurve3dElementProperty;
imported transient class HSequenceOfCurve3dElementProperty;

end;
