-- Created on: 1993-06-15
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class PaveSet from TopOpeBRepBuild 
    inherits LoopSet from TopOpeBRepBuild

---Purpose: 
-- class providing an exploration of a set of vertices to build edges.
-- It is similar to LoopSet from TopOpeBRepBuild where Loop is Pave.

uses 
    
    Shape from TopoDS,
    Edge from TopoDS,
    Loop from TopOpeBRepBuild,
    Pave from TopOpeBRepBuild,
    ListOfPave from TopOpeBRepBuild,
    ListIteratorOfListOfPave from TopOpeBRepBuild
    
is

    Create(E : Shape from TopoDS) returns PaveSet from TopOpeBRepBuild;
    ---Purpose: Create a Pave set on edge <E>. It contains <E> vertices. 

    RemovePV(me:in out; B : Boolean); -- particular case B = T/F : try/don't try
    -- to remove Pave in Prepare() (T by default)
		
    Append(me : in out; PV : Pave from TopOpeBRepBuild) is static;
    ---Purpose: Add <PV> in the Pave set.
    
    -- === start signature LoopSet
    InitLoop(me : in out) is redefined;
    MoreLoop(me) returns Boolean is redefined;
    NextLoop(me : in out) is redefined;
    Loop(me) returns Loop from TopOpeBRepBuild is redefined;
    ---C++: return const &
    -- === end signature LoopSet

    Edge(me) returns Edge from TopoDS is static;
    ---C++: return const &

    HasEqualParameters(me : in out) returns Boolean is static;
    EqualParameters(me) returns Real is static;
    ClosedVertices(me : in out) returns Boolean is static;

    Prepare(me : in out) is static private;
    SortPave(myclass; Lin:ListOfPave; Lout:out ListOfPave);
    
fields

    myEdge       : Edge from TopoDS;
    myVertices   : ListOfPave from TopOpeBRepBuild;
    myVerticesIt : ListIteratorOfListOfPave from TopOpeBRepBuild;
    myEdgeVertexIndex  : Integer from Standard;
    myEdgeVertexCount  : Integer from Standard;

    myHasEqualParameters : Boolean from Standard;
    myEqualParameters    : Real from Standard;
    myClosed             : Boolean from Standard;
    myPrepareDone        : Boolean from Standard;
    myRemovePV : Boolean;
    
end PaveSet from TopOpeBRepBuild;
