-- File:	IGESGraph_ToolTextFontDef.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolTextFontDef  from IGESGraph

    ---Purpose : Tool to work on a TextFontDef. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses TextFontDef from IGESGraph,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolTextFontDef;
    ---Purpose : Returns a ToolTextFontDef, ready to work


    ReadOwnParams (me; ent : mutable TextFontDef;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : TextFontDef;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : TextFontDef;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a TextFontDef <ent>, from
    --           its specific (own) parameters

    DirChecker (me; ent : TextFontDef) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : TextFontDef;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : TextFontDef; entto : mutable TextFontDef;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : TextFontDef;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolTextFontDef;
