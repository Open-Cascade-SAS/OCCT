-- Created on: 1995-06-12
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class ShapeListOfShape from TopOpeBRepBuild

---Purpose: represent shape + a list of shape

uses
    
    ListOfShape from TopTools,
    Shape from TopoDS
    
is

    Create returns ShapeListOfShape from TopOpeBRepBuild;

    Create(S : Shape from TopoDS)
    returns ShapeListOfShape from TopOpeBRepBuild;

    Create(S : Shape from TopoDS;
     	   L : ListOfShape from TopTools)
    returns ShapeListOfShape from TopOpeBRepBuild;

    List(me)
    returns ListOfShape from TopTools is static;
    ---C++: return const &

    ChangeList(me : in out)
    returns ListOfShape from TopTools is static;
    ---C++: return &

    Shape(me) 
    returns Shape from TopoDS is static;
    ---C++: return const &

    ChangeShape(me : in out) 
    returns Shape from TopoDS is static;
    ---C++: return &

fields

    myList : ListOfShape from TopTools;
    myShape : Shape from TopoDS;

end ShapeListOfShape from TopOpeBRepBuild;
