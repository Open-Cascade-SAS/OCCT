-- File:	RWStepShape_RWConnectedFaceShapeRepresentation.cdl
-- Created:	Fri Dec 28 16:02:00 2001 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class RWConnectedFaceShapeRepresentation from RWStepShape

    ---Purpose: Read & Write tool for ConnectedFaceShapeRepresentation

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    ConnectedFaceShapeRepresentation from StepShape

is
    Create returns RWConnectedFaceShapeRepresentation from RWStepShape;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : ConnectedFaceShapeRepresentation from StepShape);
	---Purpose: Reads ConnectedFaceShapeRepresentation

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: ConnectedFaceShapeRepresentation from StepShape);
	---Purpose: Writes ConnectedFaceShapeRepresentation

    Share (me; ent : ConnectedFaceShapeRepresentation from StepShape;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWConnectedFaceShapeRepresentation;
