-- Created on: 1993-09-14
-- Created by: Frederic MAUPAS
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class ContextTool from STEPConstruct

    ---Purpose : Gives access to Product Definition Context (one per Model)
    --           Maintains ApplicationProtocolDefinition entity (common for all
    --           products)
    --           Also maintains context specific for AP203 and provides set of
    --           methods to work with various STEP constructs as required 
    --           by Actor

uses
    SequenceOfInteger from TColStd,
    HSequenceOfTransient from TColStd,
    HAsciiString from TCollection,
    StepModel from StepData,
    ApplicationProtocolDefinition from StepBasic,
    ShapeDefinitionRepresentation from StepShape,
    Axis2Placement3d from StepGeom,
    AP203Context from STEPConstruct,
    Assembly from STEPConstruct,
    Part from STEPConstruct
    

is

    Create returns ContextTool from STEPConstruct;
    
    Create (aStepModel : StepModel from StepData) returns ContextTool from STEPConstruct;
    
    ---Management of ApplicationProtocolDefinition
    
    SetModel (me : in out; aStepModel : StepModel from StepData);
    	---Purpose: Initialize ApplicationProtocolDefinition by the first
	--          entity of that type found in the model

    GetAPD(me : in out) returns ApplicationProtocolDefinition from StepBasic;
    	---Purpose: 

    AddAPD(me : in out; enforce : Boolean = Standard_False);

    IsAP203 (me) returns Boolean;
    	---Purpose: Returns True if APD.schema_name is config_control_design

    IsAP214 (me) returns Boolean;
    	---Purpose: Returns True if APD.schema_name is automotive_design

    -- AC : Application Context

    GetACstatus(me : in out) returns HAsciiString from TCollection;
	
    GetACschemaName(me : in out) returns HAsciiString from TCollection;
	
    GetACyear(me : in out) returns Integer;

--    GetACapplication(me : in out)
--    	returns HAsciiString from TCollection;  via the SDR

    GetACname (me : in out) returns HAsciiString from TCollection;

    SetACstatus (me: in out; status: HAsciiString from TCollection);

    SetACschemaName(me: in out; schemaName: HAsciiString from TCollection);

    SetACyear (me: in out; year: Integer);

--    SetACapplication(me : in out;
--    	             application : HAsciiString from TCollection);

    SetACname (me: in out; name : HAsciiString from TCollection);

    -- Other context items

    GetDefaultAxis (me: in out) returns Axis2Placement3d from StepGeom;
    	---Purpose: Returns a default axis placement
    
    AP203Context (me: in out) returns AP203Context from STEPConstruct;
    	---Purpose: Returns tool which maintains context specific for AP203
	---C++: return &

    -- Management of assembly level for naming products
    
    Level (me) returns Integer;
        ---Purpose: Returns current assembly level

    NextLevel (me: in out);
    PrevLevel (me: in out);
    SetLevel (me: in out; lev: Integer );
        ---Purpose: Changes current assembly level

    Index (me) returns Integer;
        ---Purpose: Returns current index of assembly component on current level

    NextIndex (me: in out);
    PrevIndex (me: in out);
    SetIndex (me: in out; ind: Integer );
        ---Purpose: Changes current index of assembly component on current level

    GetProductName (me) returns HAsciiString from TCollection;
    	---Purpose: Generates a product name basing on write.step.product.name
	--          parameter and current position in the assembly structure

    -- Methods for collecting all roots corresponding to some constructs
    
    GetRootsForPart (me: in out; SDRTool: Part from STEPConstruct)
    returns HSequenceOfTransient from TColStd;
    	---Purpose: Produces and returns a full list of root entities required
	--          for part identified by SDRTool (including SDR itself)
    
    GetRootsForAssemblyLink (me: in out; assembly: Assembly from STEPConstruct)
    returns HSequenceOfTransient from TColStd;
    	---Purpose: Produces and returns a full list of root entities required
	--          for assembly link identified by assembly (including NAUO and CDSR)
    
fields

    myLevel  : SequenceOfInteger from TColStd; -- level of assembly for auto naming products
    theAPD   : ApplicationProtocolDefinition from StepBasic;
    theAP203 : AP203Context from STEPConstruct;
    myAxis   : Axis2Placement3d from StepGeom;

end ContextTool;
