-- Created on: 1998-09-07
-- Created by: Christian CAILLET
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class ActorWrite from IGESControl
    inherits ActorOfFinderProcess  from Transfer

    ---Purpose : Actor to write Shape to IGES

uses

    Finder from Transfer,
    FinderProcess from Transfer,
    Binder from Transfer

is

    Create returns ActorWrite;

    Recognize (me : mutable; start : Finder from Transfer)  returns Boolean
    	is redefined;
    ---Purpose : Recognizes a ShapeMapper

    Transfer  (me : mutable; start : Finder from Transfer;
    	       FP : mutable FinderProcess)  returns Binder  is redefined;
    ---Purpose : Transfers Shape to IGES Entities
    --         
    --           ModeTrans may be : 0 -> groups of Faces
    --           or 1 -> BRep

end ActorWrite;
