-- Created on: 2018-03-15
-- Created by: Stephan GARNAUD (ARM)
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


-- Updated:       J.P. TIRAULT August 1993
--                All methods are static methods.
--                the "Show" method returns the consumed CPU time in a Real
--                variable.
--                J.P. TIRAULT October 15 1994
--                We measure both user and system cpu time.
class Chronometer from OSD

 ---Purpose: This class measures CPU time (both user and system) consumed
 --          by current process or thread. The chronometer can be started
 --          and stopped multiple times, and measures cumulative time.
 --
 --          If only the thread is measured, calls to Stop() and Show()
 --          must occur from the same thread where Start() was called 
 --          (unless chronometer is stopped); otherwise measurement will 
 --          yield false values.

is

  Create (ThisThreadOnly: Boolean = Standard_False) returns Chronometer from OSD;
  ---Purpose: Initializes a stopped Chronometer.
  --
  --          If ThisThreadOnly is True, measured CPU time will account
  --          time of the current thread only; otherwise CPU of the 
  --          process (all threads, and completed children) is measured.
  --
  ---Level: Public

  Destroy ( me : out ) is virtual;
  ---C++: alias ~

  Reset (me : in out) is virtual;
  ---Purpose: Stops and Reinitializes the Chronometer.
  ---Level: Public

  Stop (me : in out) is virtual;
  ---Purpose: Stops the Chronometer. 
  ---Level: Public

  Start (me : in out) is virtual;
  ---Purpose: Starts (after Create or Reset) or restarts (after Stop)
  --          the chronometer.
  ---Level: Public

  Show (me : in out) is virtual;
  ---Purpose: Shows the current CPU user and system time on the 
  --          standard output stream <cout>.
  --          The chronometer can be running (laps Time) or stopped.
  ---Level: Public

  Show (me : in out; os : in out OStream from Standard) is virtual;
  ---Purpose: Shows the current CPU user and system time on the output 
  --          stream <os>.
  --          The chronometer can be running (laps Time) or stopped.
  ---Level: Public

  Show (me : in out; UserSeconds : in out Real from Standard) ;
  ---Purpose: Returns the current CPU user time in a variable.
  --          The chronometer can be running (laps Time) or stopped.
  ---Level: Public

  Show (me : in out; UserSeconds : in out Real from Standard;
                     SystemSeconds : in out Real from Standard) ;
  ---Purpose: Returns the current CPU user and system time in variables.
  --          The chronometer can be running (laps Time) or stopped.
  ---Level: Public

  GetProcessCPU (myclass; UserSeconds : out Real from Standard;
                          SystemSeconds : out Real from Standard);
  ---Purpose: Returns CPU time (user and system) consumed by the current
  --          process since its start, in seconds. The actual precision of 
  --          the measurement depends on granularity provided by the system,
  --          and is platform-specific.
  ---Level: Public
  
  GetThreadCPU (myclass; UserSeconds : out Real from Standard;
                         SystemSeconds : out Real from Standard);
  ---Purpose: Returns CPU time (user and system) consumed by the current
  --          thread since its start. Note that this measurement is
  --          platform-specific, as threads are implemented and managed 
  --          differently on different platforms and CPUs.
  ---Level: Advanced
  
fields

  Stopped    : Boolean is protected;
  ThreadOnly : Boolean;
  Start_user : Real;
  Start_sys  : Real;
  Cumul_user : Real;
  Cumul_sys  : Real;

end;


