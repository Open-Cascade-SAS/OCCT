-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ReversibleTopologyItem from StepShape inherits SelectType from StepData

	-- <ReversibleTopologyItem> is an EXPRESS Select Type construct translation.
	-- it gathers : Edge, Path, Face, FaceBound, ClosedShell, OpenShell

uses

	Edge,
	Path,
	Face,
	FaceBound,
	ClosedShell,
	OpenShell
is

	Create returns ReversibleTopologyItem;
	---Purpose : Returns a ReversibleTopologyItem SelectType

	CaseNum (me; ent : Transient) returns Integer;
	---Purpose: Recognizes a ReversibleTopologyItem Kind Entity that is :
	--        1 -> Edge
	--        2 -> Path
	--        3 -> Face
	--        4 -> FaceBound
	--        5 -> ClosedShell
	--        6 -> OpenShell
	--        0 else

	Edge (me) returns any Edge;
	---Purpose : returns Value as a Edge (Null if another type)

	Path (me) returns any Path;
	---Purpose : returns Value as a Path (Null if another type)

	Face (me) returns any Face;
	---Purpose : returns Value as a Face (Null if another type)

	FaceBound (me) returns any FaceBound;
	---Purpose : returns Value as a FaceBound (Null if another type)

	ClosedShell (me) returns any ClosedShell;
	---Purpose : returns Value as a ClosedShell (Null if another type)

	OpenShell (me) returns any OpenShell;
	---Purpose : returns Value as a OpenShell (Null if another type)


end ReversibleTopologyItem;

