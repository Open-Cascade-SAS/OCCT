-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class BSplineSurfaceWithKnotsAndRationalBSplineSurface from StepGeom 

inherits BSplineSurface from StepGeom 


	--- This classe is an implementation of EXPRESS
	--  ANDOR Subtype Declaration.
uses

	BSplineSurfaceWithKnots from StepGeom, 
	RationalBSplineSurface from StepGeom, 
	HAsciiString from TCollection, 
	Integer from Standard, 
	HArray2OfCartesianPoint from StepGeom, 
	BSplineSurfaceForm from StepGeom, 
	Logical from StepData, 
	HArray1OfInteger from TColStd, 
	HArray1OfReal from TColStd, 
	HArray2OfReal from TColStd, 
	KnotType from StepGeom
is

	Create returns BSplineSurfaceWithKnotsAndRationalBSplineSurface;
	---Purpose: Returns a BSplineSurfaceWithKnotsAndRationalBSplineSurface


	Init (me : mutable;
	      aName : HAsciiString from TCollection;
	      aUDegree : Integer from Standard;
	      aVDegree : Integer from Standard;
	      aControlPointsList : HArray2OfCartesianPoint from StepGeom;
	      aSurfaceForm : BSplineSurfaceForm from StepGeom;
	      aUClosed : Logical from StepData;
	      aVClosed : Logical from StepData;
	      aSelfIntersect : Logical from StepData) is redefined;

	Init (me : mutable;
	      aName : HAsciiString from TCollection;
	      aUDegree : Integer from Standard;
	      aVDegree : Integer from Standard;
	      aControlPointsList : HArray2OfCartesianPoint from StepGeom;
	      aSurfaceForm : BSplineSurfaceForm from StepGeom;
	      aUClosed : Logical from StepData;
	      aVClosed : Logical from StepData;
	      aSelfIntersect : Logical from StepData;
	      aBSplineSurfaceWithKnots : BSplineSurfaceWithKnots from StepGeom;
	      aRationalBSplineSurface : RationalBSplineSurface from StepGeom) is virtual;

	Init (me : mutable;
	      aName : HAsciiString from TCollection;
	      aUDegree : Integer from Standard;
	      aVDegree : Integer from Standard;
	      aControlPointsList : HArray2OfCartesianPoint from StepGeom;
	      aSurfaceForm : BSplineSurfaceForm from StepGeom;
	      aUClosed : Logical from StepData;
	      aVClosed : Logical from StepData;
	      aSelfIntersect : Logical from StepData;
	      aUMultiplicities : HArray1OfInteger from TColStd;
	      aVMultiplicities : HArray1OfInteger from TColStd;
	      aUKnots : HArray1OfReal from TColStd;
	      aVKnots : HArray1OfReal from TColStd;
	      aKnotSpec : KnotType from StepGeom;
	      aWeightsData : HArray2OfReal from TColStd) is virtual;

	-- Specific Methods for Field Data Access --

	SetBSplineSurfaceWithKnots(me : mutable; aBSplineSurfaceWithKnots : BSplineSurfaceWithKnots);
	BSplineSurfaceWithKnots (me) returns BSplineSurfaceWithKnots;
	SetRationalBSplineSurface(me : mutable; aRationalBSplineSurface : RationalBSplineSurface);
	RationalBSplineSurface (me) returns RationalBSplineSurface;

	-- Specific Methods for ANDOR Field Data Access --

	SetUMultiplicities(me : mutable; aUMultiplicities : HArray1OfInteger);
	UMultiplicities (me) returns HArray1OfInteger;
	UMultiplicitiesValue (me; num : Integer) returns Integer;
	NbUMultiplicities (me) returns Integer;
	SetVMultiplicities(me : mutable; aVMultiplicities : HArray1OfInteger);
	VMultiplicities (me) returns HArray1OfInteger;
	VMultiplicitiesValue (me; num : Integer) returns Integer;
	NbVMultiplicities (me) returns Integer;
	SetUKnots(me : mutable; aUKnots : HArray1OfReal);
	UKnots (me) returns HArray1OfReal;
	UKnotsValue (me; num : Integer) returns Real;
	NbUKnots (me) returns Integer;
	SetVKnots(me : mutable; aVKnots : HArray1OfReal);
	VKnots (me) returns HArray1OfReal;
	VKnotsValue (me; num : Integer) returns Real;
	NbVKnots (me) returns Integer;
	SetKnotSpec(me : mutable; aKnotSpec : KnotType);
	KnotSpec (me) returns KnotType;

	-- Specific Methods for ANDOR Field Data Access --

	SetWeightsData(me : mutable; aWeightsData : HArray2OfReal);
	WeightsData (me) returns HArray2OfReal;
	WeightsDataValue (me; num1 : Integer;  num2 : Integer) returns Real;
	NbWeightsDataI (me) returns Integer;
	NbWeightsDataJ (me) returns Integer;

fields

	bSplineSurfaceWithKnots : BSplineSurfaceWithKnots from StepGeom;
	rationalBSplineSurface : RationalBSplineSurface from StepGeom;

end BSplineSurfaceWithKnotsAndRationalBSplineSurface;
