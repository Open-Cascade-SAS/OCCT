--
-- File      :  OrderedGroupWithoutBackP.cdl
-- Created   :  Sat 9 Jan 1993
-- Author    : CKY / Contract Toubro-Larsen ( Arun MENON )
--
---Copyright : MATRA-DATAVISION  1993
--

class OrderedGroupWithoutBackP from IGESBasic  inherits Group

        ---Purpose: defines OrderedGroupWithoutBackP, Type <402> Form <15>
        --          in package IGESBasic
        --          
        --          It inherits from Group

uses

        Transient        ,
        HArray1OfIGESEntity from IGESData

raises OutOfRange

is

        Create returns mutable OrderedGroupWithoutBackP;

        -- Specific Methods pertaining to the class : see Group

--
-- Class    : IGESBasic_OrderedGroupWithoutBackP
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class OrderedGroupWithoutBackP.
--
-- Reminder : A OrderedGroupWithoutBackP instance is defined by :
--            - an array of entities
--            See Group

end OrderedGroupWithoutBackP;
