-- Created on: 1992-03-05
-- Created by: Herve LEGRAND
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred generic class SurfaceTool from LProp (Surface as any) 

uses Pnt from gp,
     Vec from gp

is

    Value(myclass; S : Surface; U, V : Real; P : out Pnt);
    ---Purpose: Computes the point <P> of parameter <U> and <V> on the 
    --          Surface <C>.
     	
    D1   (myclass; S : Surface; U, V : Real; P : out Pnt; D1U, D1V : out Vec);
    ---Purpose: Computes the point <P> and first derivative <D1*> of 
    --          parameter <U> and <V> on the Surface <C>.

    D2   (myclass; S : Surface; U, V : Real; 
              P : out Pnt; D1U, D1V, D2U, D2V, DUV : out Vec);
    ---Purpose: Computes the point <P>, the first derivative <D1*> and second
    --          derivative <D2*> of parameter <U> and <V> on the Surface <C>.
    
    DN  (myclass; S : Surface; U, V : Real;  IU,  IV  :  Integer) 
    returns  Vec;
    
    Continuity(myclass; S : Surface) returns Integer;
    ---Purpose: returns the order of continuity of the Surface <C>.
    --          returns 1 : first derivative only is computable
    --          returns 2 : first and second derivative only are computable.

    Bounds(myclass; S : Surface; U1, V1, U2, V2 : out Real);
    ---Purpose: returns the bounds of the Surface.

end SurfaceTool;


