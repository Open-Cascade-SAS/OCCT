-- File:	QANewModTopOpe_Glue.cdl
-- Created:	Fri May  3 18:01:59 2001
-- Author:	Michael SAZONOV <msv@nnov.matra-dtv.fr>
-- Copyright:	SAMTECH S.A. 2001


-- sccsid[] = "@(#) QANewModTopOpe_Glue.cdl 4.0-2, 07/01/03@(#)";

-- Lastly modified by :
-- +---------------------------------------------------------------------------+
-- !       msv ! Creation                                ! 3-05-2001! 3.0-00-2!
-- !       skv ! Add gluing Solid-Solid operation        ! 5-05-2001! 3.0-00-2!
-- !       skv ! Adaptation to OCC version 5.0           ! 6-05-2003! 3.0-00-2!
-- +---------------------------------------------------------------------------+



class Glue from QANewModTopOpe inherits BooleanOperation from BRepAlgoAPI

	---Purpose: Perform the gluing topological operation.

uses
    Boolean from Standard,
    Pnt from gp,
    Shape from TopoDS,
    Vertex from TopoDS,
    Edge from TopoDS,
    Face from TopoDS,
    ListOfShape from TopTools,
    State from TopAbs,
    Substitution from BRepTools,
    MapOfShape from TopTools,
    DataMapOfShapeShape from TopTools,
    DataMapOfShapeListOfShape from TopTools,
    IndexedDataMapOfShapeListOfShape from TopTools

is

    Create (theS1,theS2 : Shape from TopoDS;
    	    theAllowCutting: Boolean from Standard = Standard_False;
    	    thePerformNow: Boolean from Standard = Standard_True)
    returns Glue from QANewModTopOpe;  
    ---Purpose: Defines 2 operands.
    --          If one of operands is Solid and another is Shell and Shell
    --          goes inside Solid, the <allowCutting> determines what to do:
    --            if True, Shell is cut by Solid during the operation;
    --            if False, Null shape is returned, IsDone() returns False.
    --          If <thePerformNow> is False then does not compute immediately.
    ---Level: Public 

    Build (me: in out)
    is redefined static;
    ---Purpose: Computation; is usefull when Create was called with thePerformNow
    --          being False
    ---Level: Public

    Generated (me: in out; theS : Shape from TopoDS)
    returns ListOfShape from TopTools is redefined static;
    ---Purpose: Returns the  list   of shapes generated   from the
    --          shape <theS>. 
    ---C++: return const & 
    ---Level: Public

    Modified (me: in out; theS : Shape from TopoDS)
    returns ListOfShape from TopTools is redefined static;
    ---Purpose: Returns the list  of shapes modified from the shape
    --          <theS>. 
    ---C++: return const & 
    ---Level: Public

    IsDeleted (me: in out; theS : Shape from TopoDS)
    returns Boolean from Standard is redefined static;
    ---Purpose: Returns True if the shape <theS> existed in one of operands
    --          and is absent in the result.
    ---Level: Public 

    HasGenerated (me)
    returns Boolean  from  Standard 
    is redefined;
    ---Purpose: Returns True if there is at leat one generated shape
    ---Level: Public

    HasModified (me)
    returns Boolean  from  Standard 
    is redefined;
    ---Purpose: Returns True if there is at leat one modified shape
    ---Level: Public

    HasDeleted (me)
    returns Boolean  from  Standard 
    is redefined;
    ---Purpose: Returns True if there is at leat one deleted shape
    ---Level: Public 
     
    

    ------------------
    -- Private methods
    ------------------

    PerformShellWire (me: in out) is private;
    ---Purpose: Performs gluing Shell-Wire
    ---Level: Private

    PerformVertex (me: in out) is private;
    ---Purpose: Performs gluing Solid-Vertex and Shell-Vertex
    ---Level: Private

    PerformShell (me: in out) is private;
    ---Purpose: Performs gluing Solid-Shell and Shell-Shell
    ---Level: Private

    PerformWires (me: in out) is private;
    ---Purpose: Performs gluing Wire-Wire
    ---Level: Private

    SubstitudeSDFaces(me:  in  out; 
       theFirstSDFace      :           Shape                      from  TopoDS; 
       theSecondSDFace     :           Shape                      from  TopoDS; 
       theNewSolid1        :  in  out  Shape                      from  TopoDS;
       theNewSolid2        :  in  out  Shape                      from  TopoDS; 
       theMapOfChangedFaces:  in  out  DataMapOfShapeListOfShape  from  TopTools)
    ---Purpose: This function performs gluing operation of same domain
    --          faces theFirstSDFace and theSecondSDFace on shapes
    --          theNewSolid1 and theNewSolid2 and returns them.
    --          theMapOfChangedFaces contains changed faces as keys and
    --          lists of their splits as items.
    ---Level: Private
    returns  Boolean  from  Standard
    is  private;

    PerformSDFaces (me: in out) is private;
    ---Purpose: Performs gluing between same domain faces of object and tool
    ---Level: Private

    CutFace (me: in out; theFace: Face from TopoDS;
    	    	     	 theListSE: ListOfShape from TopTools)
    returns Boolean from Standard is private;
    ---Purpose: For the case Solid-Shell, <aFace> is from Shell.
    --          Splits <theFace> onto faces by section edges <theListSE> and
    --          add <theFace> for substitution by list of faces which are "out"
    --          of Solid
    ---Level: Private

    ClassifyFace (me: in; theFace: Face from TopoDS;
    	    	     	  theListSE: ListOfShape from TopTools)
    returns State from TopAbs is private;
    ---Purpose: For the case Solid-Shell, <theFace> is a split of Shell's face.
    --          Returns the state of <theFace> relatively Solid.
    ---Level: Private

    SectionInsideFace (me: in out; theFace: Face from TopoDS;
    	    	     	    	   theListSE: ListOfShape from TopTools;
    	    	    	    	   theShapeNum: Integer from Standard; 
    	    	    	    	   theGenEdges: MapOfShape from TopTools)
    is private;
    ---Purpose: Inserts "internal" elements (wires, edges, vertices) computed
    --          from a list of section edges <theListSE> into <theFace>.
    ---Level: Private

    ------------------
    -- Utilities
    ------------------
    ProjPointOnEdge (myclass; thePnt: Pnt from gp; theEdge: Edge from TopoDS;
    	    	     	      thePar, theDist: out Real from Standard)
    returns Boolean from Standard;

    InsertVertexInEdge (myclass; theEdge: Edge from TopoDS;
    	    	    	    	 theVer: Vertex from TopoDS;
				 thePar: Real from Standard;
				 theNewEdge: out Edge from TopoDS);

    SplitEdgeByVertex (myclass; theEdge: Edge from TopoDS;
    	    	    	    	theVer: Vertex from TopoDS;
				thePar: Real from Standard;
				theListE: out ListOfShape from TopTools);

    CompareVertices (myclass; theV1, theV2: Vertex from TopoDS;
			      theDist: out Real from Standard)
    returns Boolean from Standard;

    FindWireOrUpdateMap (myclass; theWire: Shape from TopoDS;
	      	  theMapELW: in out IndexedDataMapOfShapeListOfShape from TopTools)
    returns Shape from TopoDS is private;
    ---C++: return const &

fields

    myCompleted: Boolean from Standard;
    myAllowCutting: Boolean from Standard;
    mySubst : Substitution from BRepTools;
    -- Map: section edge => list of all faces-ancestors from corresponding shape
    myMapSEdgeFaces1: DataMapOfShapeListOfShape from TopTools;
    myMapSEdgeFaces2: DataMapOfShapeListOfShape from TopTools;
    -- Map: section edge => face crossed by this edge (i.e., edge lies
    --      inside the face, not on boundary)
    myMapSEdgeCrossFace1: DataMapOfShapeShape from TopTools;
    myMapSEdgeCrossFace2: DataMapOfShapeShape from TopTools;
    -- Map: internal edge => list of internal wires containing this edge;
    --      it is to share wires
    myMapEdgeWires: IndexedDataMapOfShapeListOfShape from TopTools;
    myEdgesToLeave: MapOfShape from TopTools;
    myMapModif: DataMapOfShapeListOfShape from TopTools;
    myMapGener: DataMapOfShapeListOfShape from TopTools;

end Glue;

-- @@SDM: begin

-- Copyright SAMTECH ..........................................Version    3.0-00
-- Lastly modified by : skv                                    Date :  6-05-2003

-- File history synopsis (creation,modification,correction)
-- +---------------------------------------------------------------------------+
-- ! Developer !              Comments                   !   Date   ! Version  !
-- +-----------!-----------------------------------------!----------!----------+
-- !       msv ! Creation                                ! 3-05-2001! 3.0-00-2!
-- !       skv ! Add gluing Solid-Solid operation        ! 5-05-2001! 3.0-00-2!
-- !       skv ! Adaptation to OCC version 5.0           ! 6-05-2003! 3.0-00-2!
-- !  vladimir ! adaptation to CAS 5.0                   !  07/01/03!    4.0-2!
-- +---------------------------------------------------------------------------+
--
-- @@SDM: end
