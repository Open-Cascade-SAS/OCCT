-- Created on: 2001-09-14
-- Created by: Alexander GRIGORIEV
-- Copyright (c) 2001-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class NamedShapeDriver from XmlMNaming inherits ADriver from XmlMDF

        ---Purpose: 


uses
    RRelocationTable    from XmlObjMgt,
    SRelocationTable    from XmlObjMgt,
    Persistent          from XmlObjMgt,
    Element             from XmlObjMgt,
    Attribute           from TDF,
    MessageDriver       from CDM,
    ShapeSet            from BRepTools,
    LocationSet         from TopTools

is
    Create (aMessageDriver: MessageDriver from CDM)
        returns mutable NamedShapeDriver from XmlMNaming;

    NewEmpty (me)
    returns mutable Attribute from TDF
        is redefined;

    Paste(me; theSource     : Persistent from XmlObjMgt;
              theTarget     : mutable Attribute from TDF;
              theRelocTable : out RRelocationTable from XmlObjMgt)
        returns Boolean from Standard
        is redefined;

    Paste(me; theSource     : Attribute from TDF;
              theTarget     : in out Persistent from XmlObjMgt;
              theRelocTable : out SRelocationTable from XmlObjMgt)
        is redefined;

    ReadShapeSection (me: mutable; anElement: Element from XmlObjMgt);
      ---Purpose: Input the shapes from DOM element

    WriteShapeSection (me: mutable; anElement: in out Element from XmlObjMgt);
      ---Purpose: Output the shapes into DOM element

    Clear (me:mutable);
      ---Purpose: Clear myShapeSet

    GetShapesLocations(me: mutable) returns LocationSet from TopTools; 
    ---Purpose: get the format of topology  
    ---C++: return &
    ---C++: inline 
    
fields
    myShapeSet          : ShapeSet from BRepTools;

end NamedShapeDriver;
