-- Created on: 2001-09-14
-- Created by: Alexander GRIGORIEV
-- Copyright (c) 2001-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class NamedShapeDriver from XmlMNaming inherits ADriver from XmlMDF

        ---Purpose: 


uses
    RRelocationTable    from XmlObjMgt,
    SRelocationTable    from XmlObjMgt,
    Persistent          from XmlObjMgt,
    Element             from XmlObjMgt,
    Attribute           from TDF,
    MessageDriver       from CDM,
    ShapeSet            from BRepTools,
    LocationSet         from TopTools

is
    Create (aMessageDriver: MessageDriver from CDM)
        returns mutable NamedShapeDriver from XmlMNaming;

    NewEmpty (me)
    returns mutable Attribute from TDF
        is redefined;

    Paste(me; theSource     : Persistent from XmlObjMgt;
              theTarget     : mutable Attribute from TDF;
              theRelocTable : out RRelocationTable from XmlObjMgt)
        returns Boolean from Standard
        is redefined;

    Paste(me; theSource     : Attribute from TDF;
              theTarget     : in out Persistent from XmlObjMgt;
              theRelocTable : out SRelocationTable from XmlObjMgt)
        is redefined;

    ReadShapeSection (me: mutable; anElement: Element from XmlObjMgt);
      ---Purpose: Input the shapes from DOM element

    WriteShapeSection (me: mutable; anElement: in out Element from XmlObjMgt);
      ---Purpose: Output the shapes into DOM element

    Clear (me:mutable);
      ---Purpose: Clear myShapeSet

    GetShapesLocations(me: mutable) returns LocationSet from TopTools; 
    ---Purpose: get the format of topology  
    ---C++: return &
    ---C++: inline 
    
fields
    myShapeSet          : ShapeSet from BRepTools;

end NamedShapeDriver;
