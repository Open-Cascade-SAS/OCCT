-- Created on: 2002-12-12
-- Created by: data exchange team
-- Copyright (c) 2002-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class FeaAxis2Placement3d from StepFEA
inherits Axis2Placement3d from StepGeom

    ---Purpose: Representation of STEP entity FeaAxis2Placement3d

uses
    HAsciiString from TCollection,
    CartesianPoint from StepGeom,
    Direction from StepGeom,
    CoordinateSystemType from StepFEA

is
    Create returns FeaAxis2Placement3d from StepFEA;
	---Purpose: Empty constructor

    Init (me: mutable; aRepresentationItem_Name: HAsciiString from TCollection;
                       aPlacement_Location: CartesianPoint from StepGeom;
                       hasAxis2Placement3d_Axis: Boolean;
                       aAxis2Placement3d_Axis: Direction from StepGeom;
                       hasAxis2Placement3d_RefDirection: Boolean;
                       aAxis2Placement3d_RefDirection: Direction from StepGeom;
                       aSystemType: CoordinateSystemType from StepFEA;
                       aDescription: HAsciiString from TCollection);
	---Purpose: Initialize all fields (own and inherited)

    SystemType (me) returns CoordinateSystemType from StepFEA;
	---Purpose: Returns field SystemType
    SetSystemType (me: mutable; SystemType: CoordinateSystemType from StepFEA);
	---Purpose: Set field SystemType

    Description (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Description
    SetDescription (me: mutable; Description: HAsciiString from TCollection);
	---Purpose: Set field Description

fields
    theSystemType: CoordinateSystemType from StepFEA;
    theDescription: HAsciiString from TCollection;

end FeaAxis2Placement3d;
