-- Created on: 1993-07-07
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ShapeScanner from TopOpeBRep
    
    ---Purpose: Find, among the  subshapes SS of a reference shape
    --          RS, the ones which 3D box interfers with the box of
    --          a shape S (SS and S are of the same type).

uses

    ShapeEnum from TopAbs,
    Shape from TopoDS,
    ListIteratorOfListOfInteger from TColStd,
    ShapeExplorer from TopOpeBRepTool,
    BoxSort from TopOpeBRepTool

is

    Create returns ShapeScanner from TopOpeBRep;
    Clear(me:in out);
    AddBoxesMakeCOB(me:in out;S:Shape;TS:ShapeEnum;TA:ShapeEnum=TopAbs_SHAPE);
    Init(me:in out;E:Shape);
    Init(me:in out;X:in out ShapeExplorer from TopOpeBRepTool);
    More(me) returns Boolean;
    Next(me:in out);
    Current(me) returns Shape;---C++: return const &
    BoxSort(me) returns BoxSort from TopOpeBRepTool;---C++:return const &
    ChangeBoxSort(me:in out) returns BoxSort from TopOpeBRepTool;---C++:return &
    Index(me) returns Integer;
    DumpCurrent(me; OS:in out OStream) returns OStream;---C++: return &
    
fields

    myBoxSort:BoxSort from TopOpeBRepTool;
    myListIterator:ListIteratorOfListOfInteger from TColStd;
    
end ShapeScanner from TopOpeBRep;

