-- Created on: 1994-06-27
-- Created by: Frederic MAUPAS
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class HeaderRecognizer         from HeaderSection
      inherits FileRecognizer  from StepData

    ---Purpose : Recognizes STEP Standard Header Entities
    --           (FileName, FileDescription, FileSchema)

uses AsciiString from TCollection

is

    Create returns mutable HeaderRecognizer ;

    Eval (me : mutable ; key : AsciiString from TCollection)  is protected;
    ---Purpose: Recognizes data types of Header STEP Standard

end HeaderRecognizer;
