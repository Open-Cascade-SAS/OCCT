-- Created on: 1992-05-22
-- Created by: Jean Claude VAUTHIER
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class BezierSurface 

from DrawTrSurf

inherits Surface from DrawTrSurf

uses BezierSurface from Geom,
     Color from Draw,
     MarkerShape from Draw,
     Display from Draw,
     Drawable3D from Draw

is


  Create (S : BezierSurface from Geom)
        --- Purpose :
        --  creates a drawable Bezier curve from a Bezier curve of 
        --  package Geom.
     returns mutable BezierSurface from DrawTrSurf;



  Create (S : BezierSurface from Geom;
          NbUIsos, NbVIsos : Integer;
          BoundsColor, IsosColor, PolesColor : Color from Draw;
          ShowPoles : Boolean; Discret : Integer;Deflection : Real;
          DrawMode : Integer)
     returns mutable BezierSurface from DrawTrSurf;


  DrawOn (me; dis : in out Display from Draw)
     is redefined static;


  ShowPoles  (me : mutable)
     is static;


  ClearPoles (me : mutable)
     is static;
  

  FindPole(me; X,Y : Real; D : Display from Draw; Prec : Real; 
           UIndex, VIndex : in out Integer)
  is static;
  

  SetPolesColor (me : mutable; aColor : Color from Draw)
        ---C++: inline
     is static;


  PolesColor (me)  returns Color from Draw
        ---C++: inline
     is static;
    
  Copy(me) returns mutable Drawable3D from Draw
	---Purpose: For variable copy.
  is redefined;
  
  
fields

  drawPoles   : Boolean;
  polesLook  : Color from Draw;

end BezierSurface;
