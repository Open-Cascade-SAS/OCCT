-- File:	GGraphic2d_Curve.cdl
-- Created:	Thu Jul  1 10:03:27 1993
-- Author:	Jean Louis FRENKEL
--		<jlf@stylox>
-- Modified: TCL G002A, 28-11-00, new method GeomCurve(...)

---Copyright:	 Matra Datavision 1993

class Curve from GGraphic2d inherits Line from Graphic2d

	---Version:

	---Purpose: The primitive Curve

	---Keywords: Primitive, Curve
	---Warning:
	---References:

uses
	Drawer		from Graphic2d,
	Curve		from Geom2d,
	GraphicObject	from Graphic2d,
	FStream		from Aspect,
	IFStream	from Aspect
is
	--------------------------------------
	-- Category: Constructors
	--------------------------------------

	Create (aGraphicObject: GraphicObject from Graphic2d;
		aCurve: Curve from Geom2d)
	returns mutable Curve from GGraphic2d;
	---Level: Public
	---Purpose: Creates a curve.
	---Category: Constructors

	--------------------------------------
	-- Category: Inquire methods
	--------------------------------------

	GeomCurve( me ) returns Curve from Geom2d;
	---Level: Internal
	---Purpose: returns the geometric curve

	--------------------------------------
	-- Category: Draw and Pick
	--------------------------------------

	Draw (me : mutable; aDrawer: Drawer from Graphic2d)
	is static protected;
	---Level: Internal
	---Purpose: Draws the curve <me>.

	Pick (me : mutable; X, Y: ShortReal from Standard;
		aPrecision: ShortReal from Standard;
		aDrawer: Drawer from Graphic2d)
	returns Boolean from Standard is static protected;
	---Level: Internal
	---Purpose: Returns Standard_True if the curve <me> is picked,
	--	    Standard_False if not.

	----------------------------------------------------------------

	Save( me; aFStream: in out FStream from Aspect ) is virtual protected;
	Retrieve(myclass; anIFStream: in out IFStream from Aspect;
		aGraphicObject: GraphicObject from Graphic2d);

fields
	myCurve:	Curve from Geom2d;

end Curve from GGraphic2d;
