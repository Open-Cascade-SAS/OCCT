-- Created on: 1995-07-24
-- Created by: Modelistation
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PoleCurve from StdPrs 

inherits Root from Prs3d
     
  	     
    	---Purpose: A framework to provide display of Bezier or BSpline curves.

uses
    Curve        from Adaptor3d,
    Presentation from Prs3d,
    Drawer       from Prs3d,
    Length       from Quantity 

is

    --- Purpose:
    
    Add(myclass; aPresentation: Presentation from Prs3d; 
    	    	 aCurve       : Curve        from Adaptor3d;
    	    	 aDrawer      : Drawer       from Prs3d);
    	---Purpose: Defines display of BSpline and Bezier curves.
    	-- Adds the 3D curve aCurve to the
    	-- StdPrs_PoleCurve algorithm. This shape is found in
    	-- the presentation object aPresentation, and its display
    	-- attributes are set in the attribute manager aDrawer.
    	-- The curve object from Adaptor3d provides data from
    	-- a Geom curve. This makes it possible to use the
    	-- surface in a geometric algorithm.

		 
    Match(myclass; X,Y,Z    : Length from Quantity;
                   aDistance: Length from Quantity;
    	    	   aCurve   : Curve  from Adaptor3d;
    	    	   aDrawer  : Drawer from Prs3d) 
    returns Boolean from Standard;
    	---Purpose: returns true if the distance between the point (X,Y,Z) and the
    	--          broken line made of the poles is less then aDistance.


    Pick(myclass; X,Y,Z    : Length from Quantity;
    	          aDistance: Length from Quantity;
                  aCurve   : Curve  from Adaptor3d;
    	          aDrawer  : Drawer from Prs3d)
    returns Integer from Standard;
    	---Purpose: returns the pole  the most near of the point (X,Y,Z) and
    	--          returns its range. The distance between the pole and
    	--          (X,Y,Z) must be less then aDistance. If no pole corresponds, 0 is returned.

end PoleCurve from StdPrs;



