-- Created on: 1997-04-01
-- Created by: Christian CAILLET
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MarkerMember  from StepVisual    inherits SelectInt  from StepData

    ---Purpose : Defines MarkerType as unique member of MarkerSelect
    --           Works with an EnumTool

uses CString, MarkerType from StepVisual

is

    Create returns mutable MarkerMember;

    HasName (me) returns Boolean  is redefined;
    -- returns True

    Name    (me) returns CString  is redefined;
    -- returns MARKER_TYPE

    SetName (me : mutable; name : CString)  returns Boolean  is redefined;
    -- does nothing and returns True

    EnumText (me) returns CString  is redefined;
    -- returns the string counterpart of a value

    SetEnumText (me : mutable; val : Integer; text : CString)  is redefined;
    -- considers text and interprets it to set val

    SetValue  (me : mutable; val : MarkerType from StepVisual);
    -- Sets directly the good value as enum

    Value     (me) returns MarkerType from StepVisual;

end MarkerMember;
