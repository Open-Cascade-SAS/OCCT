-- Created on: 1995-03-01
-- Created by: Arnaud BOUZY
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class RadiusPresentation from DsgPrs
    	---Purpose: A framework to define display of radii.
uses
    Presentation from Prs3d,
    Pnt from gp,
    Circ from gp,
    Drawer from Prs3d,
    ArrowSide from DsgPrs,
    ExtendedString from TCollection
    	
is  
    Add( myclass; aPresentation: Presentation from Prs3d;
    	    	  aDrawer: Drawer from Prs3d;
		  aText: ExtendedString from TCollection;
                  AttachmentPoint : Pnt from gp;
		  aCircle : Circ from gp;
		  firstparam : Real;
		  lastparam : Real;
		  drawFromCenter : Boolean = Standard_True;
    	    	  reverseArrow : Boolean = Standard_False);
	---Purpose: Adds the point AttachmentPoint, the circle aCircle,
    	-- the text aText, and the parameters firstparam and
    	-- lastparam to the presentation object aPresentation.
    	-- The display attributes of these elements is defined by
    	-- the attribute manager aDrawer.
    	-- If the Boolean drawFromCenter is false, the
    	-- arrowhead will point towards the center of aCircle.
    	-- If the Boolean reverseArrow is true, the arrowhead
    	-- will point away from the attachment point.

    Add( myclass; aPresentation: Presentation from Prs3d;
    	    	  aDrawer: Drawer from Prs3d;
		  aText: ExtendedString from TCollection;
                  AttachmentPoint : Pnt from gp;
		  aCircle : Circ from gp;
		  firstparam : Real;
		  lastparam : Real;
	          ArrowSide: ArrowSide from DsgPrs;
		  drawFromCenter : Boolean = Standard_True;
    	    	  reverseArrow : Boolean = Standard_False);
	---Purpose:  Adds the point AttachmentPoint, the circle aCircle,
    	-- the text aText, and the parameters firstparam and
    	-- lastparam to the presentation object aPresentation.
    	-- The display attributes of these elements is defined by
    	-- the attribute manager aDrawer.
    	-- The value of the enumeration Arrowside determines
    	-- the type of arrow displayed: whether there will be
    	-- arrowheads at both ends or only one, for example.
    	-- If the Boolean drawFromCenter is false, the
    	-- arrowhead will point towards the center of aCircle.
    	-- If the Boolean reverseArrow is true, the arrowhead
    	-- will point away from the attachment point.
   
    Add( myclass; aPresentation: Presentation from Prs3d;
    	    	  aDrawer: Drawer from Prs3d;
		  aText: ExtendedString from TCollection;
                  AttachmentPoint : Pnt from gp; 
		  Center          : Pnt from gp; 
		  EndOfArrow      : Pnt from gp;  
	          ArrowSide: ArrowSide from DsgPrs; 
		  drawFromCenter  : Boolean = Standard_True;
    	    	  reverseArrow : Boolean = Standard_False);
	---Purpose:  Adds the circle aCircle, the text aText, the points
    	-- AttachmentPoint, Center and EndOfArrow to the
    	-- presentation object aPresentation.
    	-- The display attributes of these elements is defined by
    	-- the attribute manager aDrawer.
    	-- The value of the enumeration Arrowside determines
    	-- the type of arrow displayed: whether there will be
    	-- arrowheads at both ends or only one, for example.
    	-- If the Boolean drawFromCenter is false, the
    	-- arrowhead will point towards the center of aCircle.
    	-- If the Boolean reverseArrow is true, the arrowhead
    	-- will point away from the attachment point.
    
     
end RadiusPresentation;
