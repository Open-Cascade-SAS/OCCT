-- Created on: 1992-05-27
-- Created by: Remi LEQUETTE
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class TVertex from BRep inherits TVertex from TopoDS

	---Purpose: The TVertex from  BRep inherits  from  the TVertex
	--          from TopoDS. It contains the geometric data.
	--          
	--          The  TVertex contains a 3d point and a tolerance.
	--            
uses
    Pnt    from gp,
    TShape from TopoDS,
    ListOfPointRepresentation from BRep

is
    Create returns mutable TVertex from BRep;

    Tolerance(me) returns Real
	---C++: inline
    is static;
    
    Tolerance(me : mutable; T : Real)
	---C++: inline
    is static;
    
    UpdateTolerance(me : mutable; T : Real)
	---Purpose: Sets the tolerance  to the   max  of <T>  and  the
	--          current  tolerance.
	--          
	---C++: inline
    is static;

    Pnt(me) returns Pnt from gp
	---C++: inline
	---C++: return const &
    is static;
    
    Pnt(me : mutable; P : Pnt from gp)
	---C++: inline
    is static;
    
    Points(me) returns ListOfPointRepresentation from BRep
	---C++: inline
	---C++: return const &
    is static;
    
    ChangePoints(me : mutable) returns ListOfPointRepresentation from BRep
	---C++: inline
	---C++: return &
    is static;
    
    EmptyCopy(me) returns mutable TShape from TopoDS;
	---Purpose: Returns a copy  of the  TShape  with no sub-shapes.
    
fields

    myPnt       : Pnt from gp;
    myTolerance : Real;
    myPoints    : ListOfPointRepresentation from BRep;

end TVertex;
