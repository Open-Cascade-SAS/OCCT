-- Created on: 1993-06-03
-- Created by: fid
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package PColPGeom2d 

        ---Purpose : This package  is used to  instantiate of  several
        --         generic classes from  the package  PCollection with
        --         objects from the package PGeom2d.

uses PCollection, PGeom2d

is



    class HArray1OfCurve 
    	instantiates HArray1 from PCollection (Curve from PGeom2d);
    class HArray1OfBoundedCurve 
    	instantiates HArray1 from PCollection (BoundedCurve from PGeom2d);
    class HArray1OfBezierCurve 
    	instantiates HArray1 from PCollection (BezierCurve from PGeom2d);
    class HArray1OfBSplineCurve 
    	instantiates HArray1 from PCollection (BSplineCurve from PGeom2d);



--    class HSequenceOfCurve  
--    	instantiates HSequence from PCollection (Curve from PGeom2d);
--    class HSequenceOfBoundedCurve  
--    	instantiates HSequence from PCollection (BoundedCurve from PGeom2d);


end PColPGeom2d;
