-- File:        MappedItem.cdl
-- Created:     Fri Dec  1 11:11:22 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class MappedItem from StepRepr 

inherits RepresentationItem from StepRepr 

uses

	RepresentationMap from StepRepr, 
	HAsciiString from TCollection
is

	Create returns mutable MappedItem;
	---Purpose: Returns a MappedItem


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aMappingSource : mutable RepresentationMap from StepRepr;
	      aMappingTarget : mutable RepresentationItem from StepRepr) is virtual;

	-- Specific Methods for Field Data Access --

	SetMappingSource(me : mutable; aMappingSource : mutable RepresentationMap);
	MappingSource (me) returns mutable RepresentationMap;
	SetMappingTarget(me : mutable; aMappingTarget : mutable RepresentationItem);
	MappingTarget (me) returns mutable RepresentationItem;

fields

	mappingSource : RepresentationMap from StepRepr;
	mappingTarget : RepresentationItem from StepRepr;

end MappedItem;
