-- Created on: 1998-02-11
-- Created by: Philippe MANGIN
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



private  class SectionPlacement from BRepFill 

	---Purpose: Place a shape in a local axis coordinate         

uses 
    LocationLaw  from  BRepFill,
    Shape        from  TopoDS, 
    Trsf   from  gp

is 
   Create(Law             :  LocationLaw  from  BRepFill; 
          Section         :  Shape        from  TopoDS;  
          WithContact     :  Boolean  =  Standard_False; 
          WithCorrection  :  Boolean  =  Standard_False)  
	   ---Purpose: Automatic placement         
   returns   SectionPlacement from  BRepFill;   
    
   Create(Law             :  LocationLaw  from  BRepFill; 
          Section         :  Shape        from  TopoDS; 
	  Vertex          :  Shape        from  TopoDS;   
          WithContact     :  Boolean  =  Standard_False; 
          WithCorrection  :  Boolean  =  Standard_False)  
	   ---Purpose: Placement on vertex       
   returns   SectionPlacement from  BRepFill;     
   
   Perform(me:in  out; 
           WithContact :  Boolean;  
           WithCorrection :  Boolean;
    	   Vertex         :  Shape        from  TopoDS)   
    is  private; 
    
   Transformation(me) 
   ---C++: return const &    
   returns  Trsf  from  gp;   
    
   AbscissaOnPath(me:in  out)   
   returns  Real;

fields
    myLaw :  LocationLaw  from  BRepFill; 
    mySection  :  Shape from  TopoDS; 
    myTrsf     :  Trsf  from  gp; 
    myParam    :  Real; 
    myIndex    :  Integer;
end SectionPlacement;
