-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class CsgPrimitive from StepShape inherits SelectType from StepData

	-- <CsgPrimitive> is an EXPRESS Select Type construct translation.
	-- it gathers : Sphere, Block, RightAngularWedge, Torus, RightCircularCone, RightCircularCylinder

uses

	Sphere,
	Block,
	RightAngularWedge,
	Torus,
	RightCircularCone,
	RightCircularCylinder
is

	Create returns CsgPrimitive;
	---Purpose : Returns a CsgPrimitive SelectType

	CaseNum (me; ent : Transient) returns Integer;
	---Purpose: Recognizes a CsgPrimitive Kind Entity that is :
	--        1 -> Sphere
	--        2 -> Block
	--        3 -> RightAngularWedge
	--        4 -> Torus
	--        5 -> RightCircularCone
	--        6 -> RightCircularCylinder
	--        0 else

	Sphere (me) returns any Sphere;
	---Purpose : returns Value as a Sphere (Null if another type)

	Block (me) returns any Block;
	---Purpose : returns Value as a Block (Null if another type)

	RightAngularWedge (me) returns any RightAngularWedge;
	---Purpose : returns Value as a RightAngularWedge (Null if another type)

	Torus (me) returns any Torus;
	---Purpose : returns Value as a Torus (Null if another type)

	RightCircularCone (me) returns any RightCircularCone;
	---Purpose : returns Value as a RightCircularCone (Null if another type)

	RightCircularCylinder (me) returns any RightCircularCylinder;
	---Purpose : returns Value as a RightCircularCylinder (Null if another type)


end CsgPrimitive;

