-- Created on: 1997-12-10
-- Created by: Denis PASCAL
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Variable from PDataStd inherits Attribute from PDF

	---Purpose: Persistant variable
	--          ===================

uses HAsciiString from PCollection
is

    Create returns mutable Variable from PDataStd;

    
    Create (constant : Boolean from Standard)
    returns mutable Variable from PDataStd;
    
    Constant (me : mutable; status : Boolean from Standard);    
    Constant (me)
    returns Boolean from Standard;

    Unit(me:mutable; unit : HAsciiString from PCollection);
    Unit(me) 
    returns HAsciiString from PCollection;

fields

    isConstant : Boolean      from Standard;
    myUnit     : HAsciiString from PCollection;

end Variable;
