-- Created on: 2002-12-15
-- Created by: data exchange team
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SiUnitAndThermodynamicTemperatureUnit from StepBasic inherits SiUnit from StepBasic 

	--- This class is an implementation of EXPRESS
	--  ANDOR Subtype Declaration.
uses

    ThermodynamicTemperatureUnit from StepBasic, 
    DimensionalExponents from StepBasic, 
    SiPrefix from StepBasic, 
    SiUnitName from StepBasic

is

    Create returns mutable SiUnitAndThermodynamicTemperatureUnit;
	---Purpose: Returns a SiUnitAndThermodynamicTemperatureUnit

    Init (me: mutable; aDimensions: mutable DimensionalExponents from StepBasic)
    is redefined;

    Init (me: mutable; hasAprefix: Boolean from Standard;
		       aPrefix   : SiPrefix from StepBasic;
		       aName     : SiUnitName from StepBasic) is redefined ;

    -- Specific Methods for Field Data Access --

    SetThermodynamicTemperatureUnit(me: mutable; aThermodynamicTemperatureUnit: mutable ThermodynamicTemperatureUnit);
    
    ThermodynamicTemperatureUnit (me) returns mutable ThermodynamicTemperatureUnit;

fields

    thermodynamicTemperatureUnit : ThermodynamicTemperatureUnit from StepBasic;

end SiUnitAndSolidAngleUnit;
