-- Created on: 1996-08-30
-- Created by: Yves FRICAUD
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

--  Modified by skv - Fri Dec 26 16:53:16 2003 OCC4455

class Inter2d from BRepOffset 

	---Purpose: Computes the intersections betwwen edges on a face
	--          stores result is SD as AsDes from BRepOffset.

uses
    AsDes               from BRepAlgo,
    Offset              from BRepOffset,
    Face                from TopoDS,
    IndexedMapOfShape          from TopTools,
    DataMapOfShapeShape from TopTools,
    Real                from Standard

is
    Compute(myclass ; AsDes    : mutable AsDes      from BRepAlgo;
    	    	      F        :         Face       from TopoDS;
       	    	      NewEdges :         IndexedMapOfShape from TopTools;
		      Tol      :         Real       from Standard);
		      
      	---Purpose: Computes the intersections between the edges stored
      	--          is AsDes as descendants of <F> . Intersections is computed
      	--          between two edges if one of them is bound in NewEdges.

    
    --  Modified by skv - Fri Dec 26 16:53:16 2003 OCC4455 Begin
    --  Add another parameter: offset value.
    ConnexIntByInt(myclass ; 
      	    	   FI    :          Face                from TopoDS;
    	    	   OFI   : in out   Offset              from BRepOffset;
		   MES   : in out   DataMapOfShapeShape from TopTools;  
		   Build :          DataMapOfShapeShape from TopTools;  
		   AsDes : mutable  AsDes               from BRepAlgo; 
    	    	   Offset:          Real                from Standard;
    	    	   Tol   :          Real                from Standard);
    --  Modified by skv - Fri Dec 26 16:53:16 2003 OCC4455 End
			    
end Inter2d;

