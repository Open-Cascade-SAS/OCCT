-- Created on: 1993-05-06
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



deferred class Polygo from IntPatch

	---Purpose: 

inherits Polygon2d from Intf

uses Pnt2d from gp,
     Box2d from Bnd

raises OutOfRange from Standard

is

    Initialize (theError : Real from Standard = 0.0)
        returns Polygo from IntPatch;

    Error (me) returns Real from Standard;
    ---C++: inline

    NbPoints (me) returns Integer is deferred;

    Point (me; Index : Integer) returns Pnt2d from gp is deferred;

    DeflectionOverEstimation (me)
    returns Real from Standard is redefined virtual;
    ---C++: inline
    ---Purpose: Returns the tolerance of the polygon.

    NbSegments (me)
    returns Integer from Standard is redefined virtual;
    ---C++: inline
    ---Purpose: Returns the number of Segments in the polyline.

    Segment (me; theIndex : in Integer from Standard;
                 theBegin, theEnd : in out Pnt2d from gp)
        raises OutOfRange from Standard is redefined virtual;
    ---C++: inline
    ---Purpose: Returns the points of the segment <Index> in the Polygon.

    Dump (me);

fields

    myError : Real from Standard is protected;

end Polygo;
