-- Created on: 1997-01-22
-- Created by: Prestataire Michael ALEONARD
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class SymmetricPresentation from DsgPrs
    	---Purpose: A framework to define display of symmetry between shapes.
uses
    Presentation from Prs3d,
    Pnt  from gp,
    Dir  from gp,
    Lin  from gp,
    Circ from gp,
    Drawer from Prs3d,
    ExtendedString from TCollection
    	
is  
    Add( myclass; aPresentation: Presentation from Prs3d;
    	    	  aDrawer: Drawer from Prs3d;
	       	  AttachmentPoint1: Pnt from gp;
		  AttachmentPoint2: Pnt from gp;
		  aDirection1: Dir from gp;  
		  aAxis: Lin from gp;
		  OffsetPoint: Pnt from gp);
	---Purpose: Adds the points OffsetPoint, AttachmentPoint1,
    	-- AttachmentPoint2, the direction aDirection1 and the
    	-- axis anAxis to the presentation object aPresentation.
    	-- The display attributes of the symmetry are defined by
    	-- the attribute manager aDrawer.
    	-- This syntax is used for display of symmetries between two segments.
		  
     
    Add( myclass; aPresentation: Presentation from Prs3d;
    	    	  aDrawer: Drawer from Prs3d;
	       	  AttachmentPoint1: Pnt from gp;
		  AttachmentPoint2: Pnt from gp; 
		  aCircle1: Circ from gp;
		  aAxis: Lin from gp;
		  OffsetPoint: Pnt from gp);
	---Purpose: Adds the points OffsetPoint, AttachmentPoint1,
    	-- AttachmentPoint2, the direction aDirection1 the circle
    	-- aCircle1 and the axis anAxis to the presentation
    	-- object aPresentation.
    	-- The display attributes of the symmetry are defined by
    	-- the attribute manager aDrawer.
    	-- This syntax is used for display of symmetries between two arcs.
	  
    Add( myclass; aPresentation: Presentation from Prs3d;
    	    	  aDrawer: Drawer from Prs3d;
	       	  AttachmentPoint1: Pnt from gp;
		  AttachmentPoint2: Pnt from gp; 
	          aAxis: Lin from gp;
	          OffsetPoint: Pnt from gp);
	---Purpose: Adds the points OffsetPoint, AttachmentPoint1,
    	-- AttachmentPoint2 and the axis anAxis to the
    	-- presentation object aPresentation.
    	-- The display attributes of the symmetry are defined by
    	-- the attribute manager aDrawer.
    	-- This syntax is used for display of symmetries between two vertices.
		  
end SymmetricPresentation;









