-- Created on: 1993-06-08
-- Created by: Laurent BOURESCHE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class Iterator from BRepSweep

	---Purpose: This class provides iteration services required by
	--          the Generating Line (TopoDS Shape) of a BRepSweep.
	--          This   tool is  used  to   iterate  on the  direct
	--          sub-shapes of a Shape.
	--          

uses

    Iterator from TopoDS,
    Shape from TopoDS,
    Orientation from TopAbs

raises

    NoMoreObject from Standard,
    NoSuchObject from Standard

is

    Create;

    Init(me : in out; aShape: Shape from TopoDS)
	---Purpose: Resest the Iterator on sub-shapes of <aShape>.
    is static;
    
    More(me) returns Boolean
	---Purpose: Returns True if there is a current sub-shape.
	--          
	---C++: inline
    is static;
    
    Next(me : in out)
	---Purpose: Moves to the next sub-shape.
    raises
    	NoMoreObject from Standard
    is static;
    
    Value(me) returns Shape from TopoDS
	---Purpose: Returns the current sub-shape.
    raises
    	NoSuchObject from Standard
	---C++: return const &
	---C++: inline
    is static;
    
    Orientation(me) returns Orientation from TopAbs
	---Purpose: Returns the orientation of the current sub-shape.
    raises
    	NoSuchObject from Standard
	---C++: inline
    is static;

fields

    myIterator : Iterator from TopoDS;

end Iterator from BRepSweep;
