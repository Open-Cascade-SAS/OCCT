-- Created on: 1993-01-26
-- Created by: Laurent PAINNOT
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




package AdvApprox
    
     ---Purpose: This package provides algorithms approximating a function
     --          that can be multidimensional creating in the end a 
     --          BSpline function with the required continuity
     --          
               
uses gp,
     math,
     GeomAbs,
     TColStd, 
     TColgp, 
     TCollection, 
     Standard,
     StdFail, 
     PLib

    
is
    

    class ApproxAFunction from AdvApprox ;
    ---Purpose:
    -- this approximate a given function
    class SimpleApprox; 
--  class ApproxAFunction;  

    imported EvaluatorFunction ;
    ---Purpose:
    --  typedef  void (*EvaluatorFunction)  (
    --  Standard_Integer *
    --  Standard_Real    *
    --  Standard_Real    *
    --  Standard_Integer *
    --  Standard_Real    *
    --  Standard_Integer *) ;
    

    deferred class Cutting;
    ---Purpose : 
    -- this class is used to choose the way of cutting if needed 

    class DichoCutting;
    ---Purpose :
    -- inherits class Cutting;
    -- if Cutting is necessary in [a,b], we cut at (a+b) / 2.
    -- 

    class PrefCutting;
    ---Purpose : 
    -- inherits class Cutting; contains a list of preferential points (di)i
    -- if Cutting is necessary in [a,b], we cut at the di nearest from (a+b)/2.
    
    class PrefAndRec;
    ---Purpose : 
    -- inherits class Cutting; contains two lists of preferential points to
    -- manage to level of preferential cutting.
    -- if Cutting is necessary in [a,b], we cut at the di nearest from (a+b)/2


end AdvApprox;
