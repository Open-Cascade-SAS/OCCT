-- Created on: 1993-01-09
-- Created by: CKY / Contract Toubro-Larsen ( Anand NATRAJAN )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ExternalReferenceFile from IGESBasic  inherits IGESEntity

        ---Purpose: defines ExternalReferenceFile, Type <406> Form <12>
        --          in package IGESBasic
        --          References definitions residing in another file

uses

        HAsciiString from TCollection,
        HArray1OfHAsciiString from Interface

raises OutOfRange

is

        Create returns mutable ExternalReferenceFile;

        -- Specific Methods pertaining to the class

        Init (me : mutable; aNameArray : HArray1OfHAsciiString);
        ---Purpose : This method is used to set the fields of the class
        --           ExternalReferenceFile
        --       - aNameArray : External Reference File Names

        NbListEntries (me) returns Integer;
        ---Purpose : returns number of External Reference File Names

        Name (me; Index : Integer) returns HAsciiString from TCollection
        raises OutOfRange;
        ---Purpose : returns External Reference File Name
        -- raises exception if Index <= 0 or Index > NbListEntries()

fields

--
-- Class    : IGESBasic_ExternalReferenceFile
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class ExternalReferenceFile.
--
-- Reminder : A ExternalReferenceFile instance is defined by :
--            - External Reference File Names

        theNames : HArray1OfHAsciiString;

end ExternalReferenceFile;
