-- File:        EdgeLoop.cdl
-- Created:     Fri Dec  1 11:11:19 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class EdgeLoop from StepShape 

inherits Loop from StepShape 
-- WARNING : Multiple EXPRESS inheritance
-- Not yet automaticly managed
-- inherits Path from StepShape 


-- Hand made changes : All the attributes theoricly inherited from the Path
-- entity are explicitly declared in the EdgeLoop entity.
-- The path is not directly referenced by any other entities. As far as
-- Path supertype, topological representation item, is also a 
-- supertype of Edge, this mapping is equivalent.

uses

    	HAsciiString          from TCollection,
	HArray1OfOrientedEdge from StepShape, 
	OrientedEdge          from StepShape

is

	Create returns mutable EdgeLoop;
	---Purpose: Returns a EdgeLoop

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aEdgeList : mutable HArray1OfOrientedEdge from StepShape);

	-- Specific Methods for Field Data Access --

	SetEdgeList(me : mutable; aEdgeList : mutable HArray1OfOrientedEdge);
	EdgeList (me) returns mutable HArray1OfOrientedEdge;
	EdgeListValue (me; num : Integer) returns mutable OrientedEdge;
	NbEdgeList (me) returns Integer;

fields

	edgeList : HArray1OfOrientedEdge from StepShape;

end EdgeLoop;
