-- File:	StepElement_SurfaceSectionFieldConstant.cdl
-- Created:	Thu Dec 12 17:29:04 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class SurfaceSectionFieldConstant from StepElement
inherits SurfaceSectionField from StepElement

    ---Purpose: Representation of STEP entity SurfaceSectionFieldConstant

uses
    SurfaceSection from StepElement

is
    Create returns SurfaceSectionFieldConstant from StepElement;
	---Purpose: Empty constructor

    Init (me: mutable; aDefinition: SurfaceSection from StepElement);
	---Purpose: Initialize all fields (own and inherited)

    Definition (me) returns SurfaceSection from StepElement;
	---Purpose: Returns field Definition
    SetDefinition (me: mutable; Definition: SurfaceSection from StepElement);
	---Purpose: Set field Definition

fields
    theDefinition: SurfaceSection from StepElement;

end SurfaceSectionFieldConstant;
