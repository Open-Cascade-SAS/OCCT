-- Created on: 1993-03-01
-- Created by: Philippe DAUTRY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class TrimmedCurve from PGeom inherits BoundedCurve from PGeom

        ---Purpose :
        --  Defines a portion of a curve limited by two values of 
        --  parameters inside the parametric domain of the curve.
        --  
	---See Also : TrimmedCurve from Geom.


uses Curve from PGeom

is


  Create returns mutable TrimmedCurve from PGeom;
	---Purpose: Creates a TrimmedCurve with default values.
    	---Level: Internal 


  Create (
    	aBasisCurve: Curve from PGeom;
    	aFirstU, aLastU: Real from Standard)
     returns mutable TrimmedCurve from PGeom;
        ---Purpose : Creates a TrimmedCurve with these field values.
    	---Level: Internal 


  FirstU(me : mutable; aFirstU: Real from Standard);
        ---Purpose : Set the value of the field firstU with <aFirstU>.
    	---Level: Internal 


  FirstU(me) returns Real from Standard;
        ---Purpose : Returns the value of the field firstU.
    	---Level: Internal 


  LastU(me : mutable; aLastU: Real from Standard);
        ---Purpose : Set the value of the field lastU with <aLastU>.
    	---Level: Internal 


  LastU(me) returns Real from Standard;
        ---Purpose : Returns the value of the field lastU.
    	---Level: Internal 


  BasisCurve (me: mutable; aBasisCurve: Curve from PGeom);
        ---Purpose : Set the value of the field basisCurve with <aBasisCurve>.
        --  This curve can be a trimmed curve.
    	---Level: Internal 


  BasisCurve (me) returns Curve from PGeom;
        ---Purpose : Returns the value of the field basisCurve. 
        --  This curve can be a trimmed curve.
    	---Level: Internal 


fields

    basisCurve : Curve from PGeom;
    firstU     : Real from Standard;
    lastU      : Real from Standard;

end;
