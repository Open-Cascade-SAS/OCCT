-- Created on: 1992-02-07
-- Created by: Laurent PAINNOT
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



generic class DoubleTab from math (Item as any)
uses Address from Standard
is

    Create(LowerRow, UpperRow, LowerCol, UpperCol: Integer)
    	returns DoubleTab;

    Create(Tab : Item; LowerRow, UpperRow, LowerCol, UpperCol: Integer)
    	returns DoubleTab;

    Init(me : in out; InitValue: Item) is static;

    Create(Other: DoubleTab)
    	returns DoubleTab;

    Allocate(me : in out) is private;
    
    Copy(me; Other: in out DoubleTab)
    	---C++: inline
    is static;

    
    SetLowerRow(me: in out; LowerRow: Integer)
    is static;


    SetLowerCol(me: in out; LowerCol: Integer)
    is static;

        
    Value(me; RowIndex, ColIndex: Integer)
    	---C++: alias operator()
    	---C++: return &
    	---C++: inline
      returns Item
      is static;		
	
	
    Free(me: in out)
        ---C++: alias ~

    is static;
    
    
fields

Addr        : Address;
isAllocated : Boolean;
LowR        : Integer;
UppR        : Integer;
LowC        : Integer;
UppC        : Integer;

end DoubleTab;	
