-- Created on: 1993-03-10
-- Created by: JCV
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class VectorWithMagnitude from Geom inherits Vector from Geom

        ---Purpose :
        --  Defines a vector with magnitude.
        --  A vector with magnitude can have a zero length.

uses Pnt       from gp,
     Trsf      from gp,
     Vec       from gp,
     Geometry  from Geom

raises ConstructionError from Standard

is

  Create (V : Vec) returns mutable VectorWithMagnitude;
        ---Purpose : Creates a transient copy of V.


  Create (X, Y, Z : Real)   returns mutable VectorWithMagnitude;
        ---Purpose : Creates a vector with three cartesian coordinates. 


  Create (P1, P2 : Pnt)   returns mutable VectorWithMagnitude;
        ---Purpose :
        --  Creates a vector from the point P1 to the point P2.
        --  The magnitude of the vector is the distance between P1 and P2




  SetCoord (me : mutable; X, Y, Z : Real);
        ---Purpose :  Assigns the values X, Y and Z to the coordinates of this vector.


  SetVec (me : mutable; V : Vec);
    	--- Purpose :  Converts the gp_Vec vector V into this vector.

  SetX (me : mutable; X : Real);
        ---Purpose : Changes the X coordinate of <me>.


  SetY (me : mutable; Y : Real);
        ---Purpose :  Changes the Y coordinate of <me>


  SetZ (me : mutable; Z : Real);
        ---Purpose : Changes the Z coordinate of <me>.


  Magnitude (me)  returns Real;
        ---Purpose : Returns the magnitude of <me>.


  SquareMagnitude (me)  returns Real;
        ---Purpose : Returns the square magnitude of <me>.


  Add (me : mutable; Other : Vector);
        ---Purpose :
        --  Adds the Vector Other to <me>.


  Added (me; Other : Vector)  returns mutable VectorWithMagnitude
        ---Purpose :
        --  Adds the vector Other to <me>.

     is static;


  Cross (me : mutable; Other : Vector);
        ---Purpose :
        --  Computes the cross product  between <me> and Other
        --  <me> ^ Other.


  Crossed (me; Other : Vector)  returns mutable like me
        ---Purpose :
        --  Computes the cross product  between <me> and Other 
        --  <me> ^ Other. A new vector is returned.
     is static;


  CrossCross (me : mutable; V1, V2 : Vector);
        ---Purpose : 
        --  Computes the triple vector product  <me> ^ (V1 ^ V2).


  CrossCrossed (me; V1, V2 : Vector)   returns mutable like me
        ---Purpose :
        --  Computes the triple vector product  <me> ^ (V1 ^ V2).
        --  A new vector is returned.
     is static;


  Divide (me : mutable; Scalar : Real);
        ---Purpose : Divides <me> by a scalar.


  Divided (me; Scalar : Real)  returns mutable VectorWithMagnitude
        ---Purpose :
        --  Divides <me> by a scalar. A new vector is returned.
     is static;


  Multiplied (me; Scalar : Real)  returns mutable VectorWithMagnitude
        ---Purpose :
        --  Computes the product of the vector <me> by a scalar.
        --  A new vector is returned.

     is static;


  Multiply (me : mutable; Scalar : Real);
        ---Purpose : 
        --  Computes the product of the vector <me> by a scalar.

  Normalize (me : mutable)
        ---Purpose : Normalizes <me>.
     raises ConstructionError;
        ---Purpose : 
        --  Raised if the magnitude of the vector is lower or equal to
        --  Resolution from package gp.


  Normalized (me)  returns mutable VectorWithMagnitude
        ---Purpose : Returns a copy of <me> Normalized.
     raises ConstructionError
        ---Purpose :
        --  Raised if the magnitude of the vector is lower or equal to
        --  Resolution from package gp.
     is static;


  Subtract (me : mutable; Other : Vector);
        ---Purpose : Subtracts the Vector Other to <me>.


  Subtracted (me; Other : Vector)  returns mutable VectorWithMagnitude
        ---Purpose :
        --  Subtracts the vector Other to <me>. A new vector is returned.

     is static;



  Transform (me: mutable; T : Trsf);

    	---Purpose: Applies the transformation T to this vector.


  Copy (me)  returns mutable like me;
    	---Purpose: Creates a new object which is a copy of this vector.

end;
