-- Created on: 2002-11-19
-- Created by: Vladimir ANIKIN
-- Copyright (c) 2002-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class ApplicationDelta from TDocStd inherits TShared from MMgt

uses

	SequenceOfDocument from TDocStd,
	ExtendedString from TCollection,
	OStream from Standard

is

	Create returns ApplicationDelta from TDocStd;

	GetDocuments(me : mutable)
	returns SequenceOfDocument from TDocStd;
	---C++: return &
	---C++: inline

	GetName(me)
	returns ExtendedString from TCollection;
	---C++: return const &
	---C++: inline

    	SetName(me : mutable;
	    	theName : ExtendedString from TCollection);
	---C++: inline

	Dump(me;
	     anOS : in out OStream from Standard);

fields

	myDocuments : SequenceOfDocument from TDocStd;
	myName      : ExtendedString from TCollection;

end ApplicationDelta;
