-- Created on: 1993-04-06
-- Created by: Philippe DAUTRY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Circle from PGeom2d inherits Conic from PGeom2d

        ---Purpose : Defines a circle in 3D space.
        --         
	---See Also : Circle from Geom2d.

uses Ax22d from gp

is


  Create returns Circle from PGeom2d;
	---Purpose : Creates a circle with default values.
	---Level: Internal 


  Create (aPosition : Ax22d from gp; aRadius : Real from Standard)
    returns Circle from PGeom2d;
        ---Purpose : Creates a Circle with <aPosition> and <aRadius> as field
        --         values.
	---Level: Internal 


  Radius (me : mutable; aRadius : Real from Standard);
	---Purpose: Set the value of the field radius with <aRadius>.
	---Level: Internal 


  Radius (me) returns Real from Standard;
	---Purpose: Returns the value of the field radius.
	---Level: Internal 


fields

  radius : Real from Standard;

end;

