-- Created on: 1998-11-10
-- Created by: Igor FEOKTISTOV
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ElementsOfRefMatrix from FEmTool inherits  FunctionSet  from  math

	---Purpose: this  class  describes  the  functions  needed  for   
    	--          calculating  matrix  elements  of  RefMatrix  for  linear   
	--          criteriums  (Tension,  Flexsion  and  Jerk).
	--          Each  function  from  set  gives  value  Pi(u)'*Pj(u)'  or 
	--          Pi(u)''*Pj(u)''  or  Pi(u)'''*Pj(u)'''  for  each  i  and  j,  
    	--          where  Pi(u)  is  i-th  basis  function  of  expansion  and 
	--          (')  means  derivative.
uses 
    Vector  from  math, 
    Base  from  PLib

raises 
    ConstructionError  from  Standard

is 
    Create(TheBase  :  Base  from  PLib;  DerOrder  :  Integer  from  Standard)
    
     	--  DerOrder  is  order  of  derivative  (1,  2,  3)  
	 
    returns ElementsOfRefMatrix  from  FEmTool 
    raises  ConstructionError  from  Standard; 
    --  if  DerOrder  is  not  valid
     
    NbVariables(me)
    	---Purpose: returns the number of variables of the function. 
	--  It  is  supposed  that  NbVariables  =  1.

    returns Integer;

    
    
    NbEquations(me)
    	---Purpose: returns the number of equations of the function.

    returns Integer;
    
    
    Value(me: in out; X: Vector; F: out Vector)
    	---Purpose: computes the values <F> of the functions for the 
    	--          variable <X>.
    	--          returns True if the computation was done successfully, 
    	--          False otherwise. 
	--          F  contains  results  only  for  i<=j  in  following  order: 
	--          P0*P0,  P0*P1,  P0*P2...  P1*P1,  P1*P2,...  (upper  triangle of 
	--          matrix  {PiPj})

    returns Boolean;

fields 
    myBase  :  Base  from  PLib; 
    myDerOrder  :  Integer; 
    myNbEquations  :  Integer;

end ElementsOfRefMatrix;
