-- Created on: 1993-06-21
-- Created by: Martine LANGLOIS
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MakeBoundedCurve from GeomToStep inherits Root from GeomToStep

    ---Purpose: This class implements the mapping between classes 
    --          BoundedCurve from Geom, Geom2d and the class BoundedCurve from 
    --          StepGeom which describes a BoundedCurve from prostep.
    --          As BoundedCurve is an abstract BoundedCurve this class 
    --          is an access to the sub-class required.
  
uses BoundedCurve from Geom,
     BoundedCurve from Geom2d,
     BoundedCurve from StepGeom
     
raises NotDone from StdFail
     
is 

Create ( C : BoundedCurve from Geom ) returns MakeBoundedCurve;

Create ( C : BoundedCurve from Geom2d ) returns MakeBoundedCurve;

Value (me) returns BoundedCurve from StepGeom
    raises NotDone
    is static;
    ---C++: return const&
 
fields

    theBoundedCurve : BoundedCurve from StepGeom;
    	-- The solution from StepGeom
    	
end MakeBoundedCurve;



