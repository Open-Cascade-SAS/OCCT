-- File:        Parabola.cdl
-- Created:     Mon Dec  4 12:02:28 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWParabola from RWStepGeom

	---Purpose : Read & Write Module for Parabola

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     Parabola from StepGeom,
     EntityIterator from Interface

is

	Create returns RWParabola;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable Parabola from StepGeom);

	WriteStep (me; SW : in out StepWriter; ent : Parabola from StepGeom);

	Share(me; ent : Parabola from StepGeom; iter : in out EntityIterator);

end RWParabola;
