deferred class ExternShareable from ObjMgt 

inherits Persistent from Standard

uses HAsciiString from PCollection

is
fields

    myEntry: HAsciiString ;

end ExternShareable;
