-- Created on: 1991-05-16
-- Created by: Isabelle GRIGNON
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Int3Pln from IntAna 

	---Purpose: Intersection between 3 planes. The algorithm searches
	--          for an intersection point. If two of the planes are
	--          parallel or identical, IsEmpty returns TRUE.

uses Pln from gp,
     Pnt from gp

raises NotDone     from StdFail,
       DomainError from Standard

is

    Create
    
    	returns Int3Pln from IntAna;


    Create(P1,P2,P3 : Pln from gp)
    
    	---Purpose: Determination of the intersection point between
    	--          3 planes.

    	returns Int3Pln from IntAna;


    Perform(me: in out; P1,P2,P3 : Pln from gp)
    
    	---Purpose: Determination of the intersection point between
    	--          3 planes.

    	is static;


    IsDone(me)
    
	---Purpose: Returns True if the computation was successful.

    	returns Boolean from Standard
	---C++: inline
	is static;


    IsEmpty(me)
    
    	---Purpose: Returns TRUE if there is no intersection POINT.
    	--          If 2 planes are identical or parallel, IsEmpty
    	--          will return TRUE.

    	returns Boolean from Standard
	---C++: inline

	raises NotDone from StdFail
	--- The exception NotDone is raised when IsDone() returns False.
	is static;


    Value(me)
    
    	---Purpose: Returns the intersection point.

    	returns Pnt from gp
	---C++: inline
	---C++: return const&

   	raises NotDone     from StdFail,
               DomainError from Standard
	--- The exception NotDone is raised when IsDone() returns False.
	--- The exception Domain is raised when IsEmpty() returns False.
	
	is static;


fields

    done: Boolean from Standard;
    empt: Boolean from Standard;
    pnt : Pnt     from gp;

end Int3Pln;
