-- Created on: 1997-01-15
-- Created by: Joelle CHAUVET
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class Criterion from AdvApp2Var

uses
    Patch,Context from AdvApp2Var,
    CriterionType,CriterionRepartition from AdvApp2Var

is

    Delete(me:out) is virtual;
    ---C++: alias "Standard_EXPORT virtual ~AdvApp2Var_Criterion(){Delete() ; }"
    
    Value(me; P : in out Patch; C : Context )
     is deferred; 

    IsSatisfied(me; P : Patch ) returns Boolean
     is deferred; 

    MaxValue(me) returns Real; 

    Type(me) returns CriterionType; 

    Repartition(me) returns CriterionRepartition; 

   
fields
    myMaxValue : Real is protected;
    myType : CriterionType is protected;
    myRepartition : CriterionRepartition is protected;
    
end Criterion;
