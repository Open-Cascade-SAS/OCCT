-- Created on: 1997-11-21
-- Created by: ZOV
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

--		ZOV - Mars 30 1998


deferred class PositionLight from V3d


inherits Light from V3d  

	---Purpose: Base class for Positional, Spot and Directional Light classes

uses 

	Viewer from V3d,
	Coordinate from V3d,
	View from V3d,
	TypeOfRepresentation from V3d,
	TypeOfPickLight from V3d,
	NameOfColor from Quantity,
	Coefficient from Quantity,
	Parameter from Quantity,
	Structure from Graphic3d,
	Vertex from Graphic3d,
	Group from Graphic3d

raises BadValue from V3d

is

	Initialize( VM : mutable Viewer )  ;

        --------------------------------------------------------
        ---Category: Methods to modify the Attributes of the Light
        --------------------------------------------------------

    	SetPosition ( me : mutable; X,Y,Z : Coordinate ) is deferred;
	---Level: Public
	---Purpose: Defines the position of the light source. Should be redefined!

        SetTarget (me : mutable; X,Y,Z : Coordinate);
	---Level: Public
	---Purpose: Defines the target of the light (the center 
	--          of the sphere)

        SetRadius ( me : mutable; Radius : Parameter) raises BadValue from V3d is static;
	---Level: Public
	---Purpose: Define the radius.
	---Warning: raises BadValue from V3d if the radius is <= 0	or if the light is directional
	
        OnHideFace (me : mutable; aView : View from V3d);
	---Level: Public
	---Purpose: Calculate the position of the light, on the hide face
	--          of the picking sphere.

        OnSeeFace (me : mutable; aView : View from V3d);
	---Level: Public
	---Purpose: Calculate the position of the light, on the seen face
	--          of the picking sphere.      
	
    	  Tracking (me : mutable;  aView : View from V3d;
	    	    	    	 WathPick : TypeOfPickLight from V3d; 
    	    	    	    	 Xpix,Ypix : Integer from Standard) is static;
	---Level: Public
	---Purpose: Tracking the light position, or the light space,
	--          or the radius of the light space, that depends of
	--          initial picking "WhatPick" (see the pick method).
	--          If WhatPick is SPACELIGHT, then the parameters
	--          Xpix, Ypix are the coordinates of a translation vector.

     	---------------------------------------------------
      ---Category: Displaying methods 
      ---------------------------------------------------

        Display(me: mutable; aView: View from V3d;  Representation : TypeOfRepresentation = V3d_SIMPLE)
	is virtual;
	---Level: Public
	---Purpose: Display the graphic structure of light source
	--          in the choosen view. We have three type of representation
	--          - SIMPLE   : Only the light source is displayed.
	--          - PARTIAL  : The light source and the light space are
	--                       displayed.
	--          - COMPLETE : The light source, the light space and the
	--                       radius of light space are displayed.
	--          We can choose the "SAMELAST" as parameter of representation
	--          In this case the graphic structure representation will be 
	--          the last displayed.

        Erase(me: mutable) is static;
	---Level: Public
	---Purpose: Erase the graphic structure of light source.
	
        ---------------------------------------------------
        ---Category: Inquire methods
        ---------------------------------------------------

        Radius (me ) returns Parameter is static;
	---Level: Public
	---Purpose: Returns the radius of the picking sphere.

        SeeOrHide (me; aView: View from V3d) returns Boolean is static;
	---Level: Public
	---Purpose: Returns the visibility status
	--          If True the source is visible.
	--          If False it's hidden.

	    	Position ( me; X,Y,Z : out Coordinate ) is deferred;
	---Level: Public
	---Purpose : Returns the position of the light source.

        Target ( me; X,Y,Z : out Coordinate) is static;
	---Level: Public
	---Purpose: Returns the position of the target of the light source.

        -----------------------------------------
        ---Category: Private or Protected methods
        -----------------------------------------

        Symbol ( me ; gsymbol : mutable Group from Graphic3d ;
                      aView   : View from V3d ) is deferred private;
	---Level: Internal
	---Purpose: Defines representation of the light source.



fields

        MyTarget:               Vertex from Graphic3d  is protected;
        MyTypeOfRepresentation: TypeOfRepresentation from V3d  is protected;	

end PositionalLight;


