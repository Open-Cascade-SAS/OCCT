-- Created on: 1999-03-11
-- Created by: data exchange team
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ExtrudedFaceSolid from StepShape 
inherits SweptFaceSolid from StepShape

uses

    	Direction from StepGeom, 
	Real from Standard, 
	HAsciiString from TCollection, 
	FaceSurface from StepShape

is

	Create returns ExtrudedFaceSolid;
	---Purpose: Returns a ExtrudedFaceSolid


	Init (me : mutable;
	      aName : HAsciiString from TCollection;
	      aSweptArea : FaceSurface from StepShape) is redefined;

	Init (me : mutable;
	      aName : HAsciiString from TCollection;
	      aSweptArea : FaceSurface from StepShape;
	      aExtrudedDirection : Direction from StepGeom;
	      aDepth : Real from Standard) ;

	-- Specific Methods for Field Data Access --

	SetExtrudedDirection(me : mutable; aExtrudedDirection : Direction);
	ExtrudedDirection (me) returns Direction;
	SetDepth(me : mutable; aDepth : Real);
	Depth (me) returns Real;


fields

	extrudedDirection : Direction from StepGeom;
	depth : Real from Standard;

end ExtrudedFaceSolid;
