-- Created on: 1997-04-23
-- Created by: Alexander BRIVIN
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class LineAspect from VrmlConverter inherits TShared from MMgt

	---Purpose: qualifies the aspect properties for  
	--          the VRML conversation of a Curve and  a  DeflectionCurve . 

uses 

    Material    from   Vrml

is

    Create
    returns mutable LineAspect from VrmlConverter;

    ---Purpose: create a default LineAspect. 
    --  Default value: HasMaterial  =  False  - a  line  hasn't  own  material (color) 

    Create  (aMaterial: Material from Vrml; 
    	    	 OnOff: Boolean from Standard)
    returns mutable LineAspect from VrmlConverter;
 
    SetMaterial(me: mutable; aMaterial: Material from Vrml)
    is static;
 
    Material(me) returns mutable Material from Vrml 
    is  static; 

    SetHasMaterial(me: mutable; OnOff: Boolean from Standard)
    ---Purpose: defines the necessary of writing  own  Material from Vrml into  output  OStream. 
    --          By default False  -  the material is not writing into OStream, 
    --          True  -  the material is writing. 
    is  static; 

    HasMaterial(me) returns Boolean from Standard 
    ---Purpose: returns True if the  materials is  writing into OStream.
    is static;
 
--    Copy (me)  returns mutable like me;
    
fields
     
    myMaterial		:	Material    from   Vrml;    
    myHasMaterial       :       Boolean  from  Standard;
    
end LineAspect;
