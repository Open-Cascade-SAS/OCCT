-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SiUnit from StepBasic 

inherits NamedUnit from StepBasic 

uses

	SiPrefix from StepBasic, 
	SiUnitName from StepBasic, 
	DimensionalExponents from StepBasic, 
	Boolean from Standard
is

	Create returns mutable SiUnit;
	---Purpose: Returns a SiUnit


	Init (me : mutable;
	      aDimensions : mutable DimensionalExponents from StepBasic) is redefined;

	Init (me : mutable;
	      hasAprefix : Boolean from Standard;
	      aPrefix : SiPrefix from StepBasic;
	      aName : SiUnitName from StepBasic) is virtual;

	-- Specific Methods for Field Data Access --

	SetPrefix(me : mutable; aPrefix : SiPrefix);
	UnSetPrefix (me:mutable);
	Prefix (me) returns SiPrefix;
	HasPrefix (me) returns Boolean;
	SetName(me : mutable; aName : SiUnitName);
	Name (me) returns SiUnitName;
	SetDimensions(me : mutable; aDimensions : mutable DimensionalExponents) is redefined;
	Dimensions (me) returns mutable DimensionalExponents is redefined;

fields

	prefix : SiPrefix from StepBasic; -- an Enumeration   -- OPTIONAL can be NULL
	name : SiUnitName from StepBasic; -- an Enumeration
	hasPrefix : Boolean from Standard;

 -- 
 -- NB : field <dimensions> inherited from classe <named_unit> is redeclared.
 --      it shall appears in a physical file as a *.
 --

end SiUnit;
