-- Created on: 1992-01-21
-- Created by: GG
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class OrthographicView from V3d

        ---Version:

	---Purpose: Define an orthographic view.
        --          See the methods of the Class View

        ---Keywords: View,Orthographic

        ---Warning:

        ---References:


inherits View from V3d

uses

	Viewer from V3d,
	PerspectiveView from V3d

is

    	Create ( VM : mutable Viewer ) returns mutable OrthographicView; 
	---Level : Public
	---Purpose: Define an orthographic view in the viewer VM.

    	Create ( VM : mutable Viewer ; V : PerspectiveView ) 
					returns mutable OrthographicView; 
	---Level : Public
	---Purpose: Defines an orthographic view from a Perspective view.
	--	    The parameters of the original view are duplicated
	--	    in the resulting view (Projection,Mapping,Context) .
	--	    The view thus created must be activated in a new
	--	    window.

    	Create ( VM : mutable Viewer ; V : OrthographicView ) 
					returns mutable OrthographicView; 
	---Level : Public
	---Purpose: Defines one orthographic view from another.
	--	    The parameters of the original view are duplicated 
	--	    in the resulting view. (Projection,Mapping,Context) .
	--	    The view thus created must be activated in a new window.

        Copy ( me ) returns mutable OrthographicView from V3d is static;
	---Level : Public
end OrthographicView;
