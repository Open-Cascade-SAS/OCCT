-- Created on: 1993-11-19
-- Created by: Yves FRICAUD
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class BiInt from MAT2d 

	---Purpose: BiInt is a set of two integers.
is

    Create ( I1,I2 : Integer) returns BiInt from MAT2d;
    
    FirstIndex(me) returns Integer
    is static;
    
    SecondIndex(me) returns Integer
    is static;
    
    FirstIndex(me : in out ; I1 : Integer)
    is static;
    
    SecondIndex(me : in out ; I2 : Integer)
    is static;
    
    IsEqual (me ;B : BiInt from MAT2d) returns Boolean
    	---C++: alias operator ==
    is static;
    
fields

    i1 : Integer;
    i2 : Integer;
    
end BiInt;
