-- Created on: 2012-12-06
-- Created by: Sergey KHROMOV
-- Copyright (c) 2004-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class POnSurfParams from Extrema inherits POnSurf from Extrema
    ---Purpose: Data container for point on surface parameters. These parameters
    --          are required to compute an initial approximation for extrema
    --          computation.
    
uses
    
    POnSurf     from Extrema,
    ElementType from Extrema,
    Pnt         from gp
    
is
    Create returns POnSurfParams;
	    ---Purpose: empty constructor
    	---C++: inline

    Create (theU, theV: Real from Standard; thePnt: Pnt from gp)
    	---Purpose: Creation of a point on surface with parameter 
    	--          values on the surface and a Pnt from gp.
    	---C++: inline
    returns POnSurfParams;

    SetSqrDistance(me: in out; theSqrDistance: Real from Standard);
	    ---Purpose: Sets the square distance from this point to another one
	    --          (e.g. to the point to be projected).
    	---C++: inline

    GetSqrDistance(me)
	    ---Purpose: Query the square distance from this point to another one.
    	---C++: inline
    returns Real from Standard;

    SetElementType(me: in out; theElementType: ElementType from Extrema);
	    ---Purpose: Sets the element type on which this point is situated.
    	---C++: inline

    GetElementType(me)
	    ---Purpose: Query the element type on which this point is situated.
    	---C++: inline
    returns ElementType from Extrema;
    
    SetIndices(me: in out; theIndexU: Integer from Standard;
                           theIndexV: Integer from Standard);
	    ---Purpose: Sets the U and V indices of an element that contains
	    --          this point.
    	---C++: inline

    GetIndices(me; theIndexU: out Integer from Standard;
                   theIndexV: out Integer from Standard);
	    ---Purpose: Query the U and V indices of an element that contains
	    --          this point.
    	---C++: inline

fields

    mySqrDistance : Real        from Standard;
    myElementType : ElementType from Extrema;
    myIndexU      : Integer     from Standard;
    myIndexV      : Integer     from Standard;
    
end POnSurfParams;
