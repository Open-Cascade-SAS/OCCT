-- Created on: 1993-08-18
-- Created by: Laurent BUCHARD
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



generic class QuadricCurveExactInter from IntCurveSurface (
    TheSurface        as any;
    TheSurfaceTool    as any;
    TheCurve          as any;
    TheCurveTool      as any)

    
    ---Purpose: ---------------------------------------------------------
    --                                                                 --
    --  find a root (u,v,w) from a starting point (w0) of the problem :--
    --        Q(X(w),Y(w),Z(w)) = 0                                    --
    --                                                                 --
    --  where Q(X,Y,Z) = 0    is the implicit expression of a quadric  -- 
    --  and (X(w),Y(w),Z(w)) the point of parameter w on a parametric  --
    --  curve.                                                         --
    ----------------------------------------------------------------------


uses 
    Quadric        from IntSurf,
    SequenceOfReal from TColStd

------------------------------------------------------------
class  TheQuadCurvFunc  instantiates QuadricCurveFunc from IntCurveSurface (
    Quadric        from IntSurf,
    TheCurve,
    TheCurveTool);
    
    ---Purpose: Provides the signed distance function : Q(w) 
    --          and its first derivative dQ(w)/dw
------------------------------------------------------------

is 

    Create(S: TheSurface;   C: TheCurve)
    	---Purpose: 
    returns QuadricCurveExactInter  from IntCurveSurface;


    IsDone(me)  
    	---Purpose:
    returns Boolean from Standard
    is static;
    

    NbRoots(me)
    	---Purpose: 
    returns Integer from Standard
    is static;


    Root(me; Index: Integer from Standard) 
    	---Purpose:
    returns Real from Standard
    is static; 
    
    
    NbIntervals(me)
    	---Purpose: 
    returns Integer from Standard
    is static;
    
    
    Intervals(me; Index: Integer from Standard;
                  U1,U2: out Real from Standard) 
    	---Purpose: U1 and U2 are the parameters of
    	--          a segment on the curve.
    is static;
    
    
    	
fields

    nbpnts :  Integer        from Standard;
    pnts   :  SequenceOfReal from TColStd;
    nbintv :  Integer        from Standard;
    intv   :  SequenceOfReal from TColStd;    
    
end QuadricCurveExactInter; 
