-- Created on: 1994-08-31
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class FaceInfo from Draft

	---Purpose: 

uses Surface  from Geom,
     Curve    from Geom,
     Face     from TopoDS


raises DomainError from Standard

is

    Create
    
    	returns FaceInfo from Draft;


    Create(S: Surface from Geom; HasNewGeometry: Boolean from Standard)
    
    	returns FaceInfo from Draft;


    RootFace(me: in out; F: Face from TopoDS)
    
    	is static;


    NewGeometry(me)
    
    	returns Boolean from Standard
	is static;
	

    Add(me: in out; F: Face from TopoDS)
    
    	is static;

    FirstFace(me)
    
    	returns Face from TopoDS
	---C++: return const&
	is static;


    SecondFace(me)
    
    	returns Face from TopoDS
	---C++: return const&
	is static;


    Geometry(me)
    
    	returns Surface from Geom
	is static;
	---C++: return const&

    ChangeGeometry(me: in out)
    
    	returns Surface from Geom
	is static;
	---C++: return &

    RootFace(me)
    
	---C++: return const&
    	returns Face from TopoDS
	is static;

    ChangeCurve(me: in out)
    
    	returns Curve from Geom
	---C++: return &
	is static;

    Curve(me)
    
    	returns Curve from Geom
	---C++: return const&
	is static;




fields

    myNewGeom : Boolean from Standard;
    myGeom    : Surface from Geom;
    myRootFace: Face    from TopoDS;
    myF1      : Face    from TopoDS;
    myF2      : Face    from TopoDS;
    myCurv    : Curve   from Geom;

end FaceInfo;
