-- Created on: 1993-04-06
-- Created by: Philippe DAUTRY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class CartesianPoint from PGeom2d inherits Point from PGeom2d

        ---Purpose : Point defined  in  3D space with its 3  cartesian
        --         coordinates X, Y, Z.
        --         
    	---See Also : CartesianPoint from Geom2d.

uses Pnt2d from gp

is


  Create returns CartesianPoint from PGeom2d;
        ---Purpose : Returns a CartesianPoint with default values..
	---Level: Internal 


  Create (aPnt2d : Pnt2d from gp) returns CartesianPoint from PGeom2d;
        ---Purpose : Returns a CartesianPoint built with <aPnt2d>.
	---Level: Internal 


  Pnt (me : mutable; aPnt2d : Pnt2d from gp);
        ---Purpose : Set the field Pnt2d.
	---Level: Internal 


  Pnt (me)  returns Pnt2d;
        ---Purpose : Returns the value of the field Pnt2d.
	---Level: Internal 


fields

    pnt : Pnt2d from gp;

end;
