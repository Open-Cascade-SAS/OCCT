-- File:	MeshDS_Link.cdl
-- Created:	Thu Apr 29 11:23:38 1993
-- Author:	Didier PIFFAULT
--		<dpf@phylox>
---Copyright:	 Matra Datavision 1993


deferred generic class Link from MeshDS (dummyarg as any)

	---Purpose: Describes the necessary services of  a Link  for a
	--          mesh data structure.


uses    Integer from Standard,
    	Boolean from Standard,
    	DegreeOfFreedom from MeshDS


is      Initialize     (node1, node2 : Integer from Standard;
    	    	    	canMove      : DegreeOfFreedom from MeshDS);
        ---Purpose: Contructs a Link beetween to vertices.



    	FirstNode     (me)
        ---Purpose: Give the index of first node of the Link.
    	    	    returns Integer from Standard;

    	LastNode      (me)
        ---Purpose: Give the index of Last node of the Link.
    	    	    returns Integer from Standard;

	Movability     (me)
    	    returns DegreeOfFreedom from MeshDS;

	SetMovability     (me      : in out;
    	    	    	   canMove : DegreeOfFreedom from MeshDS);

	SameOrientation(me; Other : Link from MeshDS)
	    returns Boolean from Standard;


---Purpose: For maping the Links.
--          Same Link -> Same HashCode
--          Different Links -> Not IsEqual but can have same HashCode 

    	HashCode      (me;
    	    	       Upper : Integer from Standard)
	    ---C++: function call
    	        returns Integer from Standard;
		    
    	IsEqual       (me; Other: Link from MeshDS)
	    ---C++: alias operator ==
    	    	    returns Boolean from Standard;
		    
end Link;
