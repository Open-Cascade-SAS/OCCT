-- Created on: 1995-04-24
-- Created by: Modelistation
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ChamfSpine from ChFiDS inherits Spine from ChFiDS 

	---Purpose:  Provides  data specific to chamfers 
	--         distances on  each  of faces.
uses
  ChamfMethod from ChFiDS           
 
is
    Create  returns  mutable ChamfSpine from ChFiDS;
    Create (Tol : Real from Standard) returns  mutable ChamfSpine from ChFiDS;
    
    SetDist (me : mutable; Dis : Real from Standard) is static;

    GetDist (me; Dis : in out Real from Standard) is static;    
    
    SetDists (me : mutable; Dis1, Dis2 : Real from Standard) is static;

    Dists (me; Dis1, Dis2 : in out Real from Standard) is static;

    GetDistAngle (me; 
                  Dis, Angle : in out Real from Standard;
                  DisOnF1    : in out Boolean from Standard) is static;
    
    SetDistAngle(me : mutable;
               	 Dis, Angle : Real from Standard;
                 DisOnF1    : Boolean from Standard) is static;

              
    IsChamfer(me) returns ChamfMethod from ChFiDS is static;
    	---Purpose: Return the method of chamfers used 


fields
    d1     : Real        from Standard;
    d2     : Real        from Standard;
    dison1 : Boolean     from Standard;
    angle  : Real        from Standard;
    mChamf : ChamfMethod from ChFiDS;
end ChamfSpine;



