-- Created on: 1995-02-27
-- Created by: Christian CAILLET
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class BinderOfTransientInteger  from Transfer  inherits SimpleBinderOfTransient

    ---Purpose : This type of Binder allows to attach as result, besides a
    --           Transient Object, an Integer Value, which can be an Index
    --           in the Object if it defines a List, for instance
    --           
    --           This Binder is otherwise a kind of SimpleBinderOfTransient,
    --           i.e. its basic result (for iterators, etc) is the Transient

uses Integer

is

    Create returns mutable BinderOfTransientInteger;
    ---Purpose : Creates an empty BinderOfTransientInteger; Default value for
    --           the integer part is zero

    SetInteger (me : mutable; value : Integer);
    ---Purpose : Sets a value for the integer part

    Integer (me) returns Integer;
    ---Purpose : Returns the value set for the integer part

fields

    theintval : Integer;

end BinderOfTransientInteger;
