-- Created on: 1992-11-18
-- Created by: Christian CAILLET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SelectEntityNumber  from IFSelect  inherits SelectBase

    ---Purpose : A SelectEntityNumber gets in an InterfaceModel (through a
    --           Graph), the Entity which has a specified Number (its rank of
    --           adding into the Model) : there can be zero (if none) or one.
    --           The Number is not directly defined as an Integer, but as a
    --           Parameter, which can be externally controled

uses AsciiString from TCollection, EntityIterator, Graph, IntParam

is

    Create  returns SelectEntityNumber;
    ---Purpose : Creates a SelectEntityNumber, initially with no specified Number

    SetNumber (me : mutable; num : IntParam);
    ---Purpose : Sets Entity Number to be taken (initially, none is set : 0)

    Number (me) returns IntParam;
    ---Purpose : Returns specified Number (as a Parameter)

    RootResult (me; G : Graph) returns EntityIterator;
    ---Purpose : Returns the list of selected entities : the Entity having the
    --           specified Number (this result assures naturally uniqueness)

    Label (me) returns AsciiString from TCollection;
    ---Purpose : Returns a text defining the criterium : "Entity Number ..."

fields

    thenum : IntParam;

end SelectEntityNumber;
