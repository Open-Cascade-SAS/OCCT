-- Created on: 2000-05-25
-- Created by: Peter KURNEV
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DrawableShape from BOPTest inherits DrawableShape from DBRep

    ---Purpose: 

uses  

    Shape           from TopoDS,
    Color           from Draw,
    Display         from Draw,
    Text3D          from Draw,
    Marker3D        from Draw,
    CString         from Standard,
    Pnt             from gp

is

    Create (S         : Shape from TopoDS;
    	    FreeCol   : Color from Draw;    -- color for free edges
    	    ConnCol   : Color from Draw;    -- color for shared edges
	    EdgeCol   : Color from Draw;    -- color for other edges
	    IsosCol   : Color from Draw;    -- color for Isos
	    size      : Real;               -- size for infinite isos
	    nbisos    : Integer;            -- # of isos on each face
	    discret   : Integer;            -- # of points on curves
    	    Text      : CString from Standard; 
    	    TextColor : Color from Draw
    	    )
    	returns mutable DrawableShape from BOPTest;

    Create (S         : Shape from TopoDS;
    	    Text      : CString from Standard; 
    	    TextColor : Color from Draw
    	    )
    	returns mutable DrawableShape from BOPTest; 
	
    Pnt(me) returns Pnt from gp  is private;
  
    DrawOn(me; dis : in out Display from Draw)
    is redefined;
    
fields

    myText : Text3D from Draw;
    myTextColor : Color from Draw;

end DrawableShape;
