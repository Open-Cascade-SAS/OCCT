-- Created on: 1998-06-03
-- Created by: data exchange team
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class ShellSewing from ShapeUpgrade 

    ---Purpose: This class provides a tool for applying sewing algorithm from
    --          BRepAlgo: it takes a shape, calls sewing for each shell, 
    --          and then replaces sewed shells with use of ShapeBuild_ReShape

uses 
    Shape from TopoDS,
    IndexedMapOfShape from TopTools,
    ReShape from ShapeBuild

is

    Create returns ShellSewing;
    ---Purpose: Creates a ShellSewing, empty

    ApplySewing (me: in out; shape: Shape from TopoDS; tol: Real = 0.0)
    	returns Shape from TopoDS;
    ---Purpose: Builds a new shape from a former one, by calling Sewing from
    --          BRepOffsetAPI. Rebuilt solids are oriented to be "not infinite"
    --           
    --          If <tol> is not given (i.e. value 0. by default), it is
    --          computed as the mean tolerance recorded in <shape>
    --           
    --          If no shell has been sewed, this method returns the input
    --          shape

    Init (me: in out; shape: Shape from TopoDS) is private;

    Prepare (me: in out; tol: Real) returns Integer is private;
    
    Apply (me: in out; shape: Shape from TopoDS; tol: Real) 
    returns Shape from TopoDS is private;
    
fields

    myShells: IndexedMapOfShape from TopTools;
    myReShape: ReShape from ShapeBuild;

end ShellSewing;
