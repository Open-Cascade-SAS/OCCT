-- Created on: 1993-01-09
-- Created by: CKY / Contract Toubro-Larsen ( Anand NATRAJAN )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class ExternalRefFile from IGESBasic  inherits IGESEntity

        ---Purpose: defines ExternalRefFile, Type <416> Form <1>
        --          in package IGESBasic
        --          Used when entire reference file is to be instanced

uses

        HAsciiString from TCollection

is

        Create returns mutable ExternalRefFile;

        -- Specific Methods pertaining to the class

        Init (me : mutable; aFileIdent : HAsciiString);
        ---Purpose : This method is used to set the field of the class
        --           ExternalRefFile
        --       - aFileIdent : External Reference File Identifier

        FileId (me) returns HAsciiString from TCollection;
        ---Purpose : returns External Reference File Identifier

fields

--
-- Class    : IGESBasic_ExternalRefFile
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class ExternalRefFile.
--
-- Reminder : A ExternalRefFile instance is defined by :
--            - an External Reference File Identifier

        theExtRefFileIdentifier : HAsciiString from TCollection;

end ExternalRefFile;
