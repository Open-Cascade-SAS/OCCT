-- Created on: 1995-12-15
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Face from BRepCheck inherits Result from BRepCheck

	---Purpose: 

uses Shape  from TopoDS,
     Face   from TopoDS,
     Status from BRepCheck,
     DataMapOfShapeListOfShape from TopTools

is

    Create(F: Face from TopoDS)
    
    	returns mutable Face from BRepCheck;


    InContext(me: mutable; ContextShape: Shape from TopoDS);
    


    Minimum(me: mutable);
    

    
    Blind(me: mutable);
    
    
    
    IntersectWires(me: mutable; Update: Boolean from Standard = Standard_False)
    
    	returns Status from BRepCheck
	is static;


    ClassifyWires(me: mutable; Update: Boolean from Standard = Standard_False)
    
    	returns Status from BRepCheck
	is static;



    OrientationOfWires(me: mutable; 
    	    	    	Update: Boolean from Standard = Standard_False)
    
    	returns Status from BRepCheck
	is static;


    SetUnorientable(me: mutable)
    
    	is static;


    IsUnorientable(me)
    
    	returns Boolean from Standard
	is static;

    GeometricControls(me)
    
    	returns Boolean from Standard
	is static;


    GeometricControls(me: mutable; B: Boolean from Standard)
    
	is static;



fields

    myIntdone : Boolean                   from Standard;
    myIntres  : Status                    from BRepCheck;
    myImbdone : Boolean                   from Standard;
    myImbres  : Status                    from BRepCheck;
    myOridone : Boolean                   from Standard;
    myOrires  : Status                    from BRepCheck;
    myMapImb  : DataMapOfShapeListOfShape from TopTools;
    myGctrl   : Boolean from Standard;

end Face;
