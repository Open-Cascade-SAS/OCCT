-- File:	StepFEA_SymmetricTensor43d.cdl
-- Created:	Thu Dec 12 17:51:05 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class SymmetricTensor43d from StepFEA
inherits SelectType from StepData

    ---Purpose: Representation of STEP SELECT type SymmetricTensor43d

uses
    SelectMember from StepData,
    HArray1OfReal from TColStd
    

is
    Create returns SymmetricTensor43d from StepFEA;
	---Purpose: Empty constructor

    CaseNum (me; ent: Transient) returns Integer;
	---Purpose: return 0
    
    CaseMem (me; ent: SelectMember from StepData) returns Integer is redefined;
    	---Purpose: Recognizes a items of select member CurveElementFreedomMember
	--          1 -> AnisotropicSymmetricTensor43d
	--          2 -> FeaIsotropicSymmetricTensor43d
	--          3 -> FeaIsoOrthotropicSymmetricTensor43d
	--          4 -> FeaTransverseIsotropicSymmetricTensor43d
	--          5 -> FeaColumnNormalisedOrthotropicSymmetricTensor43d
	--          6 -> FeaColumnNormalisedMonoclinicSymmetricTensor43d
	--          0 else
    
    NewMember(me) returns SelectMember from StepData is redefined;

    AnisotropicSymmetricTensor43d (me) returns HArray1OfReal from TColStd;
	---Purpose: Returns Value as AnisotropicSymmetricTensor43d (or Null if another type)
	
    SetFeaIsotropicSymmetricTensor43d(me: in out; val: HArray1OfReal from TColStd);

    FeaIsotropicSymmetricTensor43d (me) returns HArray1OfReal from TColStd;
	---Purpose: Returns Value as FeaIsotropicSymmetricTensor43d (or Null if another type)

    FeaIsoOrthotropicSymmetricTensor43d (me) returns HArray1OfReal from TColStd;
	---Purpose: Returns Value as FeaIsoOrthotropicSymmetricTensor43d (or Null if another type)

    FeaTransverseIsotropicSymmetricTensor43d (me) returns HArray1OfReal from TColStd;
	---Purpose: Returns Value as FeaTransverseIsotropicSymmetricTensor43d (or Null if another type)

    FeaColumnNormalisedOrthotropicSymmetricTensor43d (me) returns HArray1OfReal from TColStd;
	---Purpose: Returns Value as FeaColumnNormalisedOrthotropicSymmetricTensor43d (or Null if another type)

    FeaColumnNormalisedMonoclinicSymmetricTensor43d (me) returns HArray1OfReal from TColStd;
	---Purpose: Returns Value as FeaColumnNormalisedMonoclinicSymmetricTensor43d (or Null if another type)

end SymmetricTensor43d;
