-- Created on: 1992-03-09
-- Created by: Isabelle GRIGNON
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred generic class LoopPointTool from IntWalk 
    (LoopPoint as any)

	---Purpose: template class to describe the necessary ressources 
	--          for a point usedas a starting point for a marching 
	--          algorithm.
	--          The 'marching algorithm' determines the intersection 
	--          between an implicit surface and a parametrized surface.
	--          these point are inside the surface not on the boundaries.

uses Pnt from gp,
     Vec from gp,
     Dir2d from gp

is

    Value3d(myclass; PStart: LoopPoint)
    
      	---Purpose: Returns the 3d coordinates of the starting point.

    	returns Pnt from gp;


    Value2d(myclass; PStart: LoopPoint; U, V: out Real from Standard);
    
	---Purpose: Returns the <U,V> parameters which are associated 
	--          with <P>
	--          it's the parameters which start the marching algorithm


    Direction3d(myclass; PStart: LoopPoint)
    
        ---Purpose: returns the tangent at the intersectin in 3d space
        --          associated to <P>

    	returns Vec from gp;


    Direction2d(myclass; PStart: LoopPoint)
    
        ---Purpose: returns the tangent at the intersectin in the
        --          parametric space of the parametrized surface.This tangent
        --          is associated to the value2d

    	returns Dir2d from gp;


end LoopPointTool;
