-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class CartesianPoint from StepGeom 

inherits Point from StepGeom 

uses

	HArray1OfReal from TColStd, 
	Real from Standard, 
	HAsciiString from TCollection
is

	Create returns CartesianPoint;
	---Purpose: Returns a CartesianPoint


	Init (me : mutable;
	      aName : HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      aName : HAsciiString from TCollection;
	      aCoordinates : HArray1OfReal from TColStd) is virtual;

    	Init2D (me : mutable;
	      aName : HAsciiString from TCollection;
	      X,Y : Real);

    	Init3D (me : mutable;
	      aName : HAsciiString from TCollection;
	      X,Y,Z : Real);

	-- Specific Methods for Field Data Access --

	SetCoordinates(me : mutable; aCoordinates : HArray1OfReal);
	Coordinates (me) returns HArray1OfReal;
	CoordinatesValue (me; num : Integer) returns Real;
	NbCoordinates (me) returns Integer;

fields

    nbcoord : Integer; -- optimised formula
    coords  : Real[3];
--	coordinates : HArray1OfReal from TColStd;

end CartesianPoint;
