-- File:	StepFEA_ParametricCurve3dElementCoordinateDirection.cdl
-- Created:	Thu Dec 12 17:51:07 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class ParametricCurve3dElementCoordinateDirection from StepFEA
inherits FeaRepresentationItem from StepFEA

    ---Purpose: Representation of STEP entity ParametricCurve3dElementCoordinateDirection

uses
    HAsciiString from TCollection,
    Direction from StepGeom

is
    Create returns ParametricCurve3dElementCoordinateDirection from StepFEA;
	---Purpose: Empty constructor

    Init (me: mutable; aRepresentationItem_Name: HAsciiString from TCollection;
                       aOrientation: Direction from StepGeom);
	---Purpose: Initialize all fields (own and inherited)

    Orientation (me) returns Direction from StepGeom;
	---Purpose: Returns field Orientation
    SetOrientation (me: mutable; Orientation: Direction from StepGeom);
	---Purpose: Set field Orientation

fields
    theOrientation: Direction from StepGeom;

end ParametricCurve3dElementCoordinateDirection;
