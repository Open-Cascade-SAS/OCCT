-- File:	RWStepRepr_RWPropertyDefinitionRelationship.cdl
-- Created:	Thu Dec 12 17:15:59 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWPropertyDefinitionRelationship from RWStepRepr

    ---Purpose: Read & Write tool for PropertyDefinitionRelationship

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    PropertyDefinitionRelationship from StepRepr

is
    Create returns RWPropertyDefinitionRelationship from RWStepRepr;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : PropertyDefinitionRelationship from StepRepr);
	---Purpose: Reads PropertyDefinitionRelationship

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: PropertyDefinitionRelationship from StepRepr);
	---Purpose: Writes PropertyDefinitionRelationship

    Share (me; ent : PropertyDefinitionRelationship from StepRepr;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWPropertyDefinitionRelationship;
