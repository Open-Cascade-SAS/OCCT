-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package XmlMDataStd 

        ---Purpose: Storage and Retrieval drivers for modelling attributes.
        --          Transient attributes are defined in package TDataStd.

uses XmlMDF,
     XmlObjMgt,
     TDF,
     CDM

is
        ---Purpose: Storage/Retrieval drivers for TDataStd attributes
        --          =======================================

        class NameDriver;

        class IntegerDriver;
        
        class RealDriver;
        
        class IntegerArrayDriver;
        
        class RealArrayDriver;
        
        class ExtStringArrayDriver;
        
        class UAttributeDriver;
        
        class DirectoryDriver;
        
        class CommentDriver;
        
        class VariableDriver;
        
        class ExpressionDriver;
        
        class RelationDriver;
        
        class NoteBookDriver;
        
        class TreeNodeDriver;  
	
	-- Extension	 
        class TickDriver;

        -- Lists:
       class IntegerListDriver; 
       class RealListDriver;
       class ExtStringListDriver;
       class BooleanListDriver;
       class ReferenceListDriver;
    
       -- Arrays:
       class BooleanArrayDriver;
       class ReferenceArrayDriver;
       class ByteArrayDriver;


       class NamedDataDriver;  
       class AsciiStringDriver;
       class IntPackedMapDriver; 

    AddDrivers (aDriverTable : ADriverTable  from XmlMDF;
                anMsgDrv     : MessageDriver from CDM);
        ---Purpose: Adds the attribute drivers to <aDriverTable>.  
	
    SetDocumentVersion (DocVersion  : Integer from Standard); 
    
    DocumentVersion returns Integer from Standard; 	

end XmlMDataStd;
