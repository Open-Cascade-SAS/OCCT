-- Created on: 1992-01-22
-- Created by: GG
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Update:	FDA Oct 15 1994
--		ZOV - Mars 30 1998


class PositionalLight from V3d

        ---Version:

	---Purpose: Creation and modification of an isolated
	--          light source.

        ---Keywords: Light,Positional 

        ---Warning:

        ---References:


inherits PositionLight from V3d

uses 

	Viewer from V3d,
	Coordinate from V3d,
	View from V3d,
	TypeOfRepresentation from V3d,
	NameOfColor from Quantity,
	Coefficient from Quantity,
	Parameter from Quantity,
	Structure from Graphic3d,
	Vertex from Graphic3d,
	Group from Graphic3d
	
raises BadValue from V3d

is

    	Create ( VM : mutable Viewer ; X,Y,Z : Coordinate ;
		 Color : NameOfColor = Quantity_NOC_WHITE ;
		 Attenuation1 : Coefficient = 1.0 ; 
                 Attenuation2 : Coefficient = 0.0 ) 
				returns mutable PositionalLight 
        ---Level: Public
       	---Purpose: Creates an isolated light source X,Y,Z in the viewer.
    	--          It is also defined by the color Color and
    	--          two attenuation factors Attenuation1, Attenuation2.
	--	    The resulting attenuation factor determining the
	--	    illumination of a surface depends on the following
	--	    formula :
	--	    F = 1/(A1 + A2*Length)
	--		A1,A2 being the two factors of attenuation
	--	 	Length is the distance of the isolated source
	--	    from the surface.
	raises BadValue from V3d;
	---Purpose:  Warning!  raises BadValue from V3d
	--          if one of the attenuation coefficients is not between 0 et 1.

    	Create ( VM : mutable Viewer ; Xt,Yt,Zt : Coordinate;
	         Xp,Yp,Zp : Coordinate;
		 Color : NameOfColor = Quantity_NOC_WHITE ;
		 Attenuation1 : Coefficient = 1.0 ; 
                 Attenuation2 : Coefficient = 0.0 ) 
		       returns mutable PositionalLight 
	---Level: Public
	---Purpose: Creates a light source of the Positional type 
	--          in the viewer.
	--          Xt,Yt,Zt : Coordinate of Target light source.
	--          Xp,Yp,Zp : Coordinate of Position light source.
	--          The light source is also defined by the color Color
    	--          and two attenuation factors Attenuation1,
    	--          Attenuation2 that determine the illumination of a
    	--          surface using the following formula :
    	--          F = 1/(A1 + A2*Length) where:
    	--          -   A1,A2 are the two attenuation factors, and
    	--          -   Length is the distance from the isolated source.
	raises BadValue from V3d;
	---Purpose:  Warning! raises BadValue from V3d
	--          if one of the attenuation coefficients is not between 0 et 1.


        --------------------------------------------------------
        ---Category: Methods to modify the Attributes of the Light
        --------------------------------------------------------

    	SetPosition ( me : mutable; X,Y,Z : Coordinate ) is redefined;
	---Level: Public
	---Purpose: Defines the position of the light source.

	    SetAttenuation( me : mutable; A1,A2 : Coefficient ) raises BadValue from V3d is static;
	---Level: Public
	---Purpose: Defines the attenuation factors.
	--  Warning: raises BadValue from V3d
	--          if one of the attenuation coefficients is not between 0 et 1.

     	---------------------------------------------------
        ---Category: Displaying methods 
        ---------------------------------------------------

        Display(me: mutable; aView: View from V3d;
	        Representation : TypeOfRepresentation)
	is redefined static;
	---Level: Public
	---Purpose: Display the graphic structure of light source
	--          in the choosen view. We have three type of representation
	--          - SIMPLE   : Only the light source is displayed.
	--          - PARTIAL  : The light source and the light space are
	--                       displayed.
	--          - COMPLETE : The light source, the light space and the
	--                       radius of light space are displayed.
	--          We can choose the "SAMELAST" as parameter of representation
	--          In this case the graphic structure representation will be 
	--          the last displayed.
	
        ---------------------------------------------------
        ---Category: Inquire methods
        ---------------------------------------------------

    	Position ( me; X,Y,Z : out Coordinate ) is redefined static;
	---Level: Public
	---Purpose : Returns the position of the light source.

    	Attenuation ( me; A1,A2 : out Coefficient ) is static;
	---Level: Public
	---Purpose : Returns the attenuation factors A1,A2 of the light
    	-- source used at construction time.

        -----------------------------------------
        ---Category: Private or Protected methods
        -----------------------------------------

        Symbol ( me ; gsymbol : mutable Group from Graphic3d ;
                      aView   : View from V3d ) is redefined static private;
	---Level: Internal
	---Purpose: Defined the representation of the positional light source.

end PositionalLight;


