-- Created on: 2003-03-05
-- Created by: Sergey KUUL
-- Copyright (c) 2003-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Material from XCAFDoc inherits Attribute from TDF
uses
    Label from TDF,
    RelocationTable from TDF,
    HAsciiString from TCollection

is
    Create returns Material from XCAFDoc;
    
    ---Category: class methods
    --           =============

    GetID (myclass)   
    	---C++: return const &  
    returns GUID from Standard;
    
    Set (myclass; label : Label from TDF;
    	    	  aName : HAsciiString from TCollection;
    	    	  aDescription : HAsciiString from TCollection;
    	    	  aDensity : Real from Standard;
    	    	  aDensName : HAsciiString from TCollection;
    	    	  aDensValType : HAsciiString from TCollection)
    returns Material from XCAFDoc;

    Set (me : mutable; aName : HAsciiString from TCollection;
    	    	       aDescription : HAsciiString from TCollection;
    	    	       aDensity : Real from Standard;
    	    	       aDensName : HAsciiString from TCollection;
    	    	       aDensValType : HAsciiString from TCollection);
	     
    GetName (me) returns HAsciiString from TCollection;

    GetDescription (me) returns HAsciiString from TCollection;

    GetDensity (me) returns Real from Standard;

    GetDensName (me) returns HAsciiString from TCollection;

    GetDensValType (me) returns HAsciiString from TCollection;

    ID (me)
    	---C++: return const & 
    returns GUID from Standard;

    Restore (me: mutable; With : Attribute from TDF);

    NewEmpty (me)
    returns mutable Attribute from TDF;

    Paste (me; Into : mutable Attribute from TDF;
	       RT   : mutable RelocationTable from TDF);    

fields
    myName        : HAsciiString from TCollection;
    myDescription : HAsciiString from TCollection;
    myDensity     : Real from Standard;
    myDensName    : HAsciiString from TCollection;
    myDensValType : HAsciiString from TCollection;

end Material;
