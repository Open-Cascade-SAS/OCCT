-- Created on: 1994-02-03
-- Created by: Jean Marc LACHAUME
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package Geom2dHatch

uses
    Geom2dAdaptor ,
    Geom2dInt ,
    gp ,
    HatchGen

is
    
    class Intersector ;
    
    class Hatcher instantiates Hatcher from HatchGen
    	(Curve       from Geom2dAdaptor,
	 Curve       from Geom2dAdaptor,
	 Intersector from Geom2dHatch) ;

end Geom2dHatch ;
