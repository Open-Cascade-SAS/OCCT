-- Created on: 1995-12-05
-- Created by: Laurent BOURESCHE
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DegeneratedBound from GeomFill inherits Boundary from GeomFill 

	---Purpose: Description of a degenerated boundary (a point).

uses
    Pnt            from gp,
    Vec            from gp

is

    Create(Point       : Pnt from gp;
    	   First, Last : Real from Standard;
           Tol3d       : Real from Standard;
    	   Tolang      : Real from Standard)
    returns DegeneratedBound from GeomFill;

    Value(me; 
          U : Real from Standard) 
    returns Pnt from gp;

    D1(me; 
       U : Real from Standard; 
       P : out Pnt from gp; 
       V : out Vec from gp) ;

    Reparametrize(me           : mutable;
    	    	  First, Last  : Real from Standard;
                  HasDF, HasDL : Boolean from Standard;
                  DF, DL       : Real from Standard;
                  Rev          : Boolean from Standard);
		  
    Bounds(me; First, Last : out Real from Standard);

    IsDegenerated(me) returns Boolean from Standard;

fields

    myPoint : Pnt from gp;
    myFirst : Real from Standard;
    myLast  : Real from Standard;

end DegeneratedBound;
