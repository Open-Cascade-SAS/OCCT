-- Created on: 1994-03-25
-- Created by: model
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class HVertex from Adaptor3d 

	---Purpose: 


inherits TShared from MMgt

uses Pnt2d       from gp,
     Orientation from TopAbs,
     HCurve2d    from Adaptor2d

is

    Create
    
    	returns mutable HVertex from Adaptor3d;


    Create(P: Pnt2d from gp; Ori: Orientation from TopAbs;
           Resolution: Real from Standard)

    	returns mutable HVertex from Adaptor3d;


    Value(me: mutable)
    
    	returns Pnt2d from gp
    is virtual;


    Parameter(me: mutable; C: HCurve2d from Adaptor2d)
    
    	returns Real from Standard
    is virtual;


    Resolution(me: mutable; C: HCurve2d from Adaptor2d)
    
	---Purpose: Parametric resolution (2d).

    	returns Real from Standard
    is virtual;


    Orientation(me: mutable)
    
    	returns Orientation from TopAbs
    is virtual;


    IsSame(me: mutable; Other: mutable like me)
    
    	returns Boolean from Standard
    is virtual;


fields

    myPnt : Pnt2d       from gp;
    myTol : Real        from Standard;
    myOri : Orientation from TopAbs;

end HVertex;
