-- Created on: 1998-10-20
-- Created by: DCB
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class GIFAlienImage from AlienImage inherits AlienUserImage from AlienImage

uses
  GIFAlienData            from AlienImage,
  File                    from OSD,
  AsciiString             from TCollection,
  Image                   from Image

is
  Create
  returns mutable GIFAlienImage from AlienImage;

  Clear( me : in out mutable) ;
  ---Level: Public
  ---Purpose: Frees memory allocated by GIFAlienImage
  ---C++: alias ~

  SetName( me : in out mutable;
           aName : in AsciiString from TCollection) ;
  ---Level: Public
  ---Purpose: Set Image name .

  Name( me : in immutable ) returns AsciiString from TCollection ;
  ---C++: return const &
  ---Level: Public
  ---Purpose: get Image name .

  ToImage( me : in immutable ) 
  returns mutable Image from Image ;
  ---Level: Public
  ---Purpose : convert a GIFAlienImage object to a Image object.

  FromImage( me : in out mutable ; anImage : in Image from Image ) ;
  ---Level: Public
  ---Purpose : convert a Image object to a GIFAlienImage object.

  Read ( me : in out mutable; afile : in out File from OSD )
    returns Boolean from Standard ;
  ---Level: Public
  ---Purpose: Read content of a  GIFAlienImage object from a file .
  --          Returns True if file is a GIF file .

  Write( me : in immutable; afile : in out File from OSD )
  returns Boolean from Standard ;
  ---Level: Public
  ---Purpose: Write content of a  GIFAlienImage object to a file .

fields
  myData : GIFAlienData  from  AlienImage;

end;
 
