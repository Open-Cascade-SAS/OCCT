-- File:	RWStepBasic_RWGroupRelationship.cdl
-- Created:	Wed May 10 15:09:08 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class RWGroupRelationship from RWStepBasic

    ---Purpose: Read & Write tool for GroupRelationship

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    GroupRelationship from StepBasic

is
    Create returns RWGroupRelationship from RWStepBasic;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : GroupRelationship from StepBasic);
	---Purpose: Reads GroupRelationship

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: GroupRelationship from StepBasic);
	---Purpose: Writes GroupRelationship

    Share (me; ent : GroupRelationship from StepBasic;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWGroupRelationship;
