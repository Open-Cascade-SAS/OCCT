-- Created on: 2005-12-21
-- Created by: Sergey KHROMOV
-- Copyright (c) 2005-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class TFunction from BRepGProp inherits Function from math

    ---Purpose: This class represents the integrand function for the outer 
    --          integral computation. The returned value represents the 
    --          integral of UFunction. It depends on the value type and the 
    --          flag IsByPoint. 

uses

    Pnt       from gp,
    Address   from Standard,
    Boolean   from Standard,
    Integer   from Standard,
    Real      from Standard,
    ValueType from GProp,
    UFunction from BRepGProp,
    Face      from BRepGProp

is

    Create(theSurface  : Face    from BRepGProp; 
           theVertex   : Pnt     from gp; 
           IsByPoint   : Boolean from Standard; 
           theCoeffs   : Address from Standard; 
           theUMin     : Real    from Standard; 
           theTolerance: Real    from Standard) 
    ---Purpose: Constructor. Initializes the function with the face, the 
    --          location point, the flag IsByPoint, the coefficients 
    --          theCoeff that have different meaning depending on the value 
    --          of IsByPoint. The last two parameters are theUMin - the 
    --          lower bound of the inner integral. This value is fixed for 
    --          any integral. And the value of tolerance of inner integral 
    --          computation.
    --          If IsByPoint is equal to Standard_True, the number of the 
    --          coefficients is equal to 3 and they represent X, Y and Z 
    --          coordinates (theCoeff[0], theCoeff[1] and theCoeff[2] 
    --          correspondingly) of the shift if the inertia is computed 
    --          with respect to the point different then the location. 
    --          If IsByPoint is equal to Standard_False, the number of the 
    --          coefficients is 4 and they represent the compbination of 
    --          plane parameters and shift values.
    returns TFunction from BRepGProp;   

    Init(me: in out);

    SetNbKronrodPoints(me: in out; theNbPoints: Integer from Standard);
    ---Purpose: Setting the expected number of Kronrod points for the outer 
    --          integral computation. This number is required for 
    --          computation of a value of tolerance for inner integral 
    --          computation. After GetStateNumber method call, this number 
    --          is recomputed by the same law as in 
    --          math_KronrodSingleIntegration, i.e. next number of points 
    --          is equal to the current number plus a square root of the 
    --          current number. If the law in math_KronrodSingleIntegration
    --          is changed, the modification algo should be modified 
    --          accordingly.
    ---C++: inline 
 
    SetValueType(me: in out; aType: ValueType from GProp);
    ---Purpose: Setting the type of the value to be returned. This 
    --          parameter is directly passed to the UFunction. 
    ---C++: inline 

    SetTolerance(me: in out; aTol: Real from Standard);
    ---Purpose: Setting the tolerance  for  inner integration
    ---C++: inline 

    ErrorReached(me) 
    ---Purpose: Returns the relative reached error of all values computation since 
    --          the last call of GetStateNumber method.
    ---C++: inline 
    returns Real from Standard;

    AbsolutError(me) 
    ---Purpose: Returns the absolut reached error of all values computation since 
    --          the last call of GetStateNumber method.
    ---C++: inline 
    returns Real from Standard;
 
    Value(me: in out; X:     Real from Standard; 
                      F: out Real from Standard) 
    ---Purpose: Returns a value of the function. The value represents an 
    --          integral of UFunction. It is computed with the predefined 
    --          tolerance using the adaptive Gauss-Kronrod method.
    returns Boolean from Standard 
    is redefined; 
 
    GetStateNumber(me: in out) 
    ---Purpose:  Redefined  method. Remembers the error reached during 
    --           computation of integral values since the object creation 
    --           or the last call of GetStateNumber. It is invoked in each 
    --           algorithm from the package math. Particularly in the 
    --           algorithm math_KronrodSingleIntegration that is used to 
    --           compute the integral of TFunction.
    returns Integer
    is redefined;

fields

    mySurface   : Face from BRepGProp;
    myUFunction : UFunction from BRepGProp;
    myUMin      : Real      from Standard;
    myTolerance : Real      from Standard;
    myTolReached: Real      from Standard;
    myErrReached: Real      from Standard;
    myAbsError  : Real      from Standard;
    myValueType : ValueType from GProp;
    myIsByPoint : Boolean   from Standard;
    myNbPntOuter: Integer   from Standard;

end TFunction;
