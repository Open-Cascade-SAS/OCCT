-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Lin2d   from gp

        ---Purpose: Describes a line in 2D space.
        -- A line is positioned in the plane with an axis (a gp_Ax2d
        -- object) which gives the line its origin and unit vector. A
        -- line and an axis are similar objects, thus, we can convert
        -- one into the other.
        -- A line provides direct access to the majority of the edit
        -- and query functions available on its positioning axis. In
        -- addition, however, a line has specific functions for
        -- computing distances and positions.
        -- See Also
        -- GccAna and Geom2dGcc packages which provide
        -- functions for constructing lines defined by geometric
        -- constraints
        -- gce_MakeLin2d which provides functions for more
        -- complex line constructions
        -- Geom2d_Line which provides additional functions for
        -- constructing lines and works, in particular, with the
        -- parametric equations of lines


uses Ax2d   from gp,
     Dir2d  from gp, 
     Pnt2d  from gp,
     Trsf2d from gp,
     Vec2d  from gp

raises ConstructionError from Standard

is

  Create   returns Lin2d;
        ---C++:inline
        --- Purpose : Creates a Line corresponding to X axis of the
        --            reference coordinate system.

  Create (A : Ax2d)   returns Lin2d;
        ---C++:inline
        --- Purpose : Creates a line located with A.

  Create (P : Pnt2d; V : Dir2d)   returns Lin2d;
        ---C++:inline
        --- Purpose : 
        --  <P> is the location point (origin) of the line and
        --  <V> is the direction of the line.

  Create (A, B, C : Real)   returns Lin2d
        --- Purpose :
        --  Creates the line from the equation A*X + B*Y + C = 0.0 Raises ConstructionError if Sqrt(A*A + B*B) <= Resolution from gp.

     raises ConstructionError;
        --- Purpose : Raised if Sqrt(A*A + B*B) <= Resolution from gp.


  Reverse (me : in out)
        ---C++:inline
         is static;

  Reversed (me)  returns Lin2d  is static;
        ---C++:inline
        ---Purpose:
        -- Reverses the positioning axis of this line.
        -- Note:
        -- -   Reverse assigns the result to this line, while
        -- -   Reversed creates a new one.
   
  SetDirection (me : in out; V : Dir2d)
        ---C++:inline
        is static;
        --- Purpose :  Changes the direction of the line.

  SetLocation(me : in out; P : Pnt2d)
        ---C++:inline
     is static;
        --- Purpose : Changes the origin of the line.

  SetPosition (me : in out; A : Ax2d)   is static;
        ---C++:inline
        --- Purpose :
        --  Complete redefinition of the line.
        --  The "Location" point of <A> is the origin of the line.
        --  The "Direction" of <A> is  the direction of the line.

  Coefficients (me; A, B, C : out Real)   is static;
        ---C++:inline
        --- Purpose :
        --  Returns the normalized coefficients of the line :
        --  A * X + B * Y + C = 0.

  Direction (me)  returns Dir2d   is static;
        ---C++:inline
        --- Purpose : Returns the direction of the line.
    	---C++: return const&

  Location (me)   returns Pnt2d   is static;
        ---C++:inline
        --- Purpose : Returns the location point (origin) of the line.
    	---C++: return const&

  Position (me)   returns Ax2d    is static;
        --- Purpose :
        --  Returns the axis placement one axis whith the same
        --  location and direction as <me>.
        ---C++: inline
    	---C++: return const&

  Angle (me; Other : Lin2d)   returns Real   is static;
        ---C++: inline
        --- Purpose : Computes the angle between two lines in radians.

  Contains (me; P : Pnt2d; LinearTolerance : Real)   returns Boolean
     is static;
        ---C++: inline     
        --- Purpose :  Returns true if this line contains the point P, that is, if the
    	-- distance between point P and this line is less than or
    	-- equal to LinearTolerance.


  Distance (me; P : Pnt2d)   returns Real            is static;
        ---C++: inline
        --- Purpose : 
        --  Computes the distance between <me> and the point <P>.


  Distance (me; Other : Lin2d)   returns Real        is static;
        ---C++: inline
        --- Purpose : Computes the distance between two lines.


  SquareDistance (me; P : Pnt2d)   returns Real      is static;
        ---C++: inline
        --- Purpose : 
        --  Computes the square distance between <me> and the point 
        --  <P>.


  SquareDistance (me; Other : Lin2d)   returns Real  is static;
        ---C++: inline
        --- Purpose : Computes the square distance between two lines.



  Normal (me; P : Pnt2d)  returns Lin2d    is static;
        ---C++: inline
        --- Purpose :
        --  Computes the line normal to the direction of <me>,
        --  passing through the point <P>.

              

   
  Mirror (me : in out; P : Pnt2d) 
         is static;

  Mirrored (me; P : Pnt2d)  returns Lin2d  is static;

     --- Purpose :
        --  Performs the symmetrical transformation of a line 
        --  with respect to the point <P> which is the center 
        --  of the symmetry


  Mirror (me : in out; A : Ax2d) 
         is static;

  Mirrored (me; A : Ax2d)  returns Lin2d  is static;


        --- Purpose :
        --  Performs the symmetrical transformation of a line 
        --  with respect to an axis placement which is the axis 
        --  of the symmetry.


  Rotate(me : in out; P : Pnt2d; Ang : Real)
        ---C++:inline
           is static;

  Rotated (me; P : Pnt2d; Ang : Real)   returns Lin2d  is static;
        ---C++:inline

        --- Purpose :
        --  Rotates a line. P is the center of the rotation.
        --  Ang is the angular value of the rotation in radians.

  Scale (me : in out; P : Pnt2d; S : Real) 
         is static;

  Scaled (me; P : Pnt2d; S : Real)   returns Lin2d  is static;
        ---C++:inline
        --- Purpose : 
        --  Scales a line. S is the scaling value. Only the
        --  origin of the line is modified.



  Transform (me : in out; T : Trsf2d)
        ---C++:inline
             is static;

  Transformed (me; T : Trsf2d)   returns Lin2d    is static;
        ---C++:inline


        --- Purpose :
        --  Transforms a line with the transformation T from class Trsf2d.      

  Translate (me : in out; V : Vec2d)
        ---C++:inline
           is static;

  Translated (me; V : Vec2d)   returns Lin2d   is static;
        ---C++:inline



        --- Purpose :
        --  Translates a line in the direction of the vector V.
        --  The magnitude of the translation is the vector's magnitude.



  Translate (me : in out; P1, P2 : Pnt2d)           is static;
        ---C++:inline

  Translated (me; P1, P2 : Pnt2d)   returns Lin2d   is static;
        ---C++:inline


        --- Purpose :
        --  Translates a line from the point P1 to the point P2.


fields

   pos : Ax2d;

end;
