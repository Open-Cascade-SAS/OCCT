-- Created by: DAUTRY Philippe
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

--      	-------------------

---Version:	0.0
--Version	Date		Purpose
--		0.0	Sep  8 1998	Creation

class ClosureTool from TDF

	---Purpose: This class provides services to build the closure
	--          of an information set.
	--          
	--          You can set closure options by using IDFilter
	--          (to select or exclude specific attribute IDs) and
	--          CopyOption objects and by giving to Closure
	--          method.
	--          


uses

    Boolean             from Standard,
    Label               from TDF,
    Attribute           from TDF,
    DataSet             from TDF,
    RelocationTable     from TDF,
    AttributeMap        from TDF,
    LabelMap            from TDF,
    IDFilter            from TDF,
    ClosureMode         from TDF

-- raises

is

    Closure(myclass;
    	aDataSet : mutable DataSet from TDF);
	---Purpose: Builds the transitive closure of label and
	--          attribute sets into <aDataSet>.

    Closure(myclass;
    	aDataSet : mutable DataSet from TDF;
    	aFilter  : IDFilter from TDF;
    	aMode    : ClosureMode from TDF);
	---Purpose: Builds the transitive closure of label and
	--          attribute sets into <aDataSet>. Uses <aFilter> to
	--          determine if an attribute has to be taken in
	--          account or not. Uses <aMode> for various way of
	--          closing.


    -- ----------------------------------------------------------------------
    -- 
    -- Private methods
    -- 
    -- ----------------------------------------------------------------------

    Closure(myclass;
    	    aLabel   : Label        from TDF;
	    aLabMap  : in out LabelMap     from TDF;
	    anAttMap : in out AttributeMap from TDF;
    	    aFilter  : IDFilter     from TDF;
    	    aMode    : ClosureMode  from TDF);
	---Purpose: Builds the transitive closure of <aLabel>.


    LabelAttributes(myclass;
    	    	    aLabel   : Label        from TDF;
		    aLabMap  : in out LabelMap     from TDF;
		    anAttMap : in out AttributeMap from TDF;
    	    	    aFilter  : IDFilter     from TDF;
    	    	    aMode    : ClosureMode  from TDF)
    	is private;
	---Purpose: Adds label attributes and dependences.


end ClosureTool;
