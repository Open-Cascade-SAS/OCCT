-- Created on: 1992-09-22
-- Created by: Gilles DEBARBOUILLE
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Mat2d from MAT2d

	---Purpose: this class contains the generic algoritm of 
	--          computation of the bisecting locus.

uses
    Side                     from MAT,
    Bisector                 from MAT,
    ListOfEdge               from MAT,
    ListOfBisector           from MAT,
    DataMapOfIntegerBisector from MAT,
    DataMapOfIntegerInteger  from TColStd,
	Tool2d                   from MAT2d
    
is

    Create(IsOpenResult : Boolean from Standard = Standard_False)
    ---Purpose: Empty construtor.
    returns Mat2d from MAT2d;
    
--- Category : Computation.    
    
    CreateMat(me : in out ; aTool : in out Tool2d from MAT2d)
       ---Purpose: Algoritm of computation of the bisecting locus.
    is static;
    
    CreateMatOpen(me : in out ; aTool : in out Tool2d from MAT2d)
       ---Purpose: Algoritm of computation of the bisecting locus for
       --          open wire.
    is static;
    
    IsDone(me) returns Boolean from Standard
       ---Purpose:  Returns <TRUE> if CreateMat has succeeded. 
    is static;

    LoadBisectorsToRemove(me                    : in out ; 
    	    	    	  noofbisectorstoremove : in out Integer;
    	    	          distance1             :        Real;
			  distance2             :        Real;
			  bisector1             :        Bisector from MAT;
			  bisector2             :        Bisector from MAT;
			  bisector3             :        Bisector from MAT;
			  bisector4             :        Bisector from MAT)
    is static private;


    Intersect( me                   : in out                   ;
    	       atool                : in out  Tool2d from MAT2d;
    	       aside                :         Integer          ;
    	       noofbisectorstoremove: in out  Integer           ;
	       bisector1            : Bisector from MAT;
	       bisector2            : Bisector from MAT)
    is static private;	       
  			       

--- Category : Querying.    
    
    Init(me : in out)
	--- Purpose : Initialize an iterator on the set of the roots
	--            of the trees of bisectors.
    is static;
    
    More(me) returns Boolean
	--- Purpose : Return False if there is no more roots.
    is static;
    
    Next(me : in out)
	--- Purpose : Move to the next root.
    is static;
    
    Bisector(me) returns any Bisector from MAT
	--- Purpose : Returns the current root.
    is static;

    SemiInfinite(me) returns Boolean from Standard
	--- Purpose : Returns True if there are semi_infinite bisectors.
	--            So there is a tree for each semi_infinte bisector.
    is static;

    NumberOfBisectors(me) returns Integer from Standard
	--- Purpose : Returns the total number of bisectors.
    is static;

fields

    myIsOpenResult        : Boolean;
    thenumberofbisectors  : Integer;
    thenumberofedges      : Integer;
    semiInfinite          : Boolean;
    theedgelist           : ListOfEdge               from MAT;
    typeofbisectortoremove: DataMapOfIntegerInteger  from TColStd;
    bisectoronetoremove   : DataMapOfIntegerBisector from MAT;
    bisectortwotoremove   : DataMapOfIntegerBisector from MAT;
    bisectormap           : DataMapOfIntegerBisector from MAT;
    roots                 : ListOfBisector           from MAT;
    isDone                : Boolean;             
    
end Mat2d;
