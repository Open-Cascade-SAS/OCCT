-- Created on: 1994-02-18
-- Created by: Remi LEQUETTE
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




deferred class MakeSweep from BRepPrimAPI inherits MakeShape from BRepBuilderAPI

	---Purpose:  The abstract class MakeSweep is
    	-- the root class of swept primitives.
    	-- Sweeps are objects you obtain by sweeping a profile along a path.
    	-- The profile can be any topology and the path is usually a curve or
    	-- a wire. The profile generates objects according to the following rules:
    	--   -      Vertices generate Edges
    	--   -      Edges generate Faces.
    	--   -      Wires generate Shells.
    	--   -      Faces generate Solids.
    	--   -      Shells generate Composite  Solids.
    	--     You are not allowed to sweep Solids and Composite Solids.
    	-- Two kinds of sweeps are implemented in the BRepPrimAPI package:
    	--   -      The linear sweep called a   Prism
    	--   -      The rotational sweep    called a Revol
    	--   Swept constructions along complex profiles such as BSpline curves
    	-- are also available in the BRepOffsetAPI package..

uses Shape from TopoDS

is
    FirstShape (me : in out)
    	---Purpose: Returns the  TopoDS  Shape of the bottom of the sweep.
    returns Shape from TopoDS
    is deferred;

    LastShape (me : in out)
    	---Purpose: Returns the TopoDS Shape of the top of the sweep.
    returns Shape from TopoDS
    is deferred;

end MakeSweep;
