-- Created on: 2000-08-15
-- Created by: data exchange team
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class LocationStorageDriver from MXCAFDoc inherits ASDriver from MDF

	---Purpose: 

uses
    SRelocationTable from MDF,
    Attribute        from TDF,
    Attribute        from PDF,
    MessageDriver    from CDM

is

--    Create  -- Version 0
--    returns LocationStorageDriver from MXCAFDoc;
    Create (theMsgDriver : MessageDriver from CDM)
    returns LocationStorageDriver from MXCAFDoc;


    VersionNumber(me) returns Integer from Standard;
	---Purpose: Returns the version number from which the driver
	--          is available: 0.

    SourceType(me) returns Type from Standard;
	---Purpose: Returns the type: XCAFDoc_Location.

    NewEmpty (me) returns Attribute from PDF;


    Paste(me;
    	  Source     :         Attribute from TDF;
    	  Target     : Attribute from PDF;
    	  RelocTable : SRelocationTable from MDF);


end LocationStorageDriver;

    
