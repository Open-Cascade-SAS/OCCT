-- Created on: 1999-11-26
-- Created by: Andrey BETENEV
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0

class CertificationAssignment from StepBasic
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity CertificationAssignment

uses
    Certification from StepBasic

is
    Create returns CertificationAssignment from StepBasic;
	---Purpose: Empty constructor

    Init (me: mutable; aAssignedCertification: Certification from StepBasic);
	---Purpose: Initialize all fields (own and inherited)

    AssignedCertification (me) returns Certification from StepBasic;
	---Purpose: Returns field AssignedCertification
    SetAssignedCertification (me: mutable; AssignedCertification: Certification from StepBasic);
	---Purpose: Set field AssignedCertification

fields
    theAssignedCertification: Certification from StepBasic;

end CertificationAssignment;
