-- Created on: 1999-09-20
-- Created by: Peter KURNEV
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ShapeWithState from TopOpeBRepDS 

	---Purpose: 

uses
    Shape from TopoDS, 
    ListOfShape  from  TopTools,
    State from TopAbs 


is
    Create returns  ShapeWithState from TopOpeBRepDS ;
     
    Part  (me;  aState: State from TopAbs)  returns ListOfShape  from  TopTools ;  
    ---C++:  return  const& 
     
    AddPart (me:out;  aShape:Shape  from  TopoDS;  aState: State from TopAbs);  

    AddParts (me:out; aListOfShape:ListOfShape  from  TopTools;  aState: State from TopAbs);  
     
    SetState  (me:out;  aState: State from TopAbs);  
    
    State  (me)  returns  State from TopAbs; 
     
    SetIsSplitted  (me:out;  anIsSplitted:Boolean  from  Standard); 
     
    IsSplitted  (me)  returns  Boolean  from  Standard; 
    
fields
  
    myPartIn   :  ListOfShape  from  TopTools; 
    myPartOut  :  ListOfShape  from  TopTools; 
    myPartOn   :  ListOfShape  from  TopTools; 
    myState:  State from TopAbs ; 
    myIsSplitted:  Boolean  from  Standard; 
     
end ShapeWithState;
