-- File:        Colour.cdl
-- Created:     Mon Dec  4 12:02:24 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWColour from RWStepVisual

	---Purpose : Read & Write Module for Colour

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     Colour from StepVisual

is

	Create returns RWColour;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable Colour from StepVisual);

	WriteStep (me; SW : in out StepWriter; ent : Colour from StepVisual);

end RWColour;
