-- Created on: 1991-02-20
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class IntPoint from IntAna2d

    ---Purpose: Geometrical intersection between two 2d elements.


uses Pnt2d from gp

raises DomainError from Standard

is

    Create(X,Y: Real; U1,U2: Real)
    
    	---Purpose: Create an intersection point between 2 parametric 2d lines.
    	--          X,Y are the coordinate of the point. U1 is the parameter
    	--          on the first element, U2 the parameter on the second one.
    
    	returns IntPoint;


    Create(X,Y: Real; U1: Real)
    
    	---Purpose: Create an intersection point between a parametric 2d line,
    	--          and a line given by an implicit equation (ImplicitCurve).
    	--          X,Y are the coordinate of the point. U1 is the parameter
    	--          on the parametric element.
    
    	returns IntPoint;


    Create

	---Purpose: Empty constructor. It's necessary to use one of
	--          the SetValue method after this one.

    	returns IntPoint;


    SetValue(me : in out; X,Y: Real; U1,U2: Real)
    
	---Purpose: Set the values for a "non-implicit" point.
    is virtual;


    SetValue(me : in out; X,Y:Real; U1: Real)
    
	---Purpose: Set the values for an "implicit" point.
    is virtual;

    Value(me)
    
	---Purpose: Returns the geometric point.
    	---C++: inline
    	---C++: return const&
    	returns Pnt2d from gp

    is static;
    
    
    SecondIsImplicit(me)
    
    	---Purpose: Returns True if the second curve is implicit.
    	---C++: inline
    	returns Boolean from Standard
	
   is static;
	
    
    ParamOnFirst(me)
    
    	---Purpose: Returns the parameter on the first element.
    	---C++: inline
    	returns Real
	
    is static;

 
    ParamOnSecond(me)
    
    	---Purpose: Returns the parameter on the second element.
    	--          If the second element is an implicit curve, an exception
    	--          is raised.
    	---C++: inline
    	returns Real
	
	raises DomainError from Standard
    
    is static;



fields

    myu1        : Real  from Standard;
    myu2        : Real  from Standard;
    myp         : Pnt2d from gp;
    myimplicit  : Boolean from Standard;

end IntPoint;
