-- Created on: 1992-05-15
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

generic class SearchInside from IntStart (
       ThePSurface     as any;
       ThePSurfaceTool as any;
       TheTopolTool    as Transient; -- as SITopolTool from IntStart
       TheSITool       as any;
       TheFunction     as any)


	---Purpose: 

uses InteriorPoint           from IntSurf,
     SequenceOfInteriorPoint from IntSurf


raises NotDone    from StdFail,
       OutOfRange from Standard


is

    Create
    
    	returns SearchInside from IntStart;


    Create (F: in out TheFunction; Surf: ThePSurface; T: TheTopolTool;
            Epsilon : Real from Standard)
    
    	returns SearchInside from IntStart;


    Perform(me: in out; F: in out TheFunction; Surf: ThePSurface;
                        T: TheTopolTool;
                        Epsilon: Real from Standard)
    
    	is static;

    Perform(me: in out; F: in out TheFunction; Surf: ThePSurface;
                        UStart,VStart: Real from Standard)
    
    	is static;


    IsDone(me)
    
    	returns Boolean
	---C++: inline
	
	is static;


    NbPoints(me)
    
	---Purpose: Returns the number of points.
	--          The exception NotDone if raised if IsDone 
	--          returns False.
    
    	returns Integer
	---C++: inline
	
	raises NotDone from StdFail
	
	is static;


    Value(me; Index: Integer)
    
	---Purpose: Returns the point of range Index.
	--          The exception NotDone if raised if IsDone 
	--          returns False.
	--          The exception OutOfRange if raised if
	--          Index <= 0 or Index > NbPoints.

    	returns InteriorPoint from IntSurf
	---C++: return const&
	---C++: inline
	
	raises NotDone from StdFail,
	       OutOfRange from Standard

    	is static;


fields

    done : Boolean                 from Standard;
    list : SequenceOfInteriorPoint from IntSurf;

end SearchInside;
