-- File:        BoxedHalfSpace.cdl
-- Created:     Mon Dec  4 12:02:24 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWBoxedHalfSpace from RWStepShape

	---Purpose : Read & Write Module for BoxedHalfSpace

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     BoxedHalfSpace from StepShape,
     EntityIterator from Interface

is

	Create returns RWBoxedHalfSpace;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable BoxedHalfSpace from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : BoxedHalfSpace from StepShape);

	Share(me; ent : BoxedHalfSpace from StepShape; iter : in out EntityIterator);

end RWBoxedHalfSpace;
