-- File:	StepDimTol_CylindricityTolerance.cdl
-- Created:	Wed Jun  4 13:34:34 2003 
-- Author:	Galina KULIKOVA
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class CylindricityTolerance from StepDimTol
inherits GeometricTolerance from StepDimTol

    ---Purpose: Representation of STEP entity CylindricityTolerance

uses
    HAsciiString from TCollection,
    MeasureWithUnit from StepBasic,
    ShapeAspect from StepRepr

is
    Create returns CylindricityTolerance from StepDimTol;
	---Purpose: Empty constructor

end CylindricityTolerance;
