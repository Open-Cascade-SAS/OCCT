-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class GeometricSetSelect from StepShape inherits SelectType from StepData

	-- <GeometricSetSelect> is an EXPRESS Select Type construct translation.
	-- it gathers : Point, Curve, Surface

uses

	Point   from StepGeom,
	Curve   from StepGeom,
	Surface from StepGeom
is

	Create returns GeometricSetSelect;
	---Purpose : Returns a GeometricSetSelect SelectType

	CaseNum (me; ent : Transient) returns Integer;
	---Purpose: Recognizes a GeometricSetSelect Kind Entity that is :
	--        1 -> Point
	--        2 -> Curve
	--        3 -> Surface
	--        0 else

	Point (me) returns any Point;
	---Purpose : returns Value as a Point (Null if another type)

	Curve (me) returns any Curve;
	---Purpose : returns Value as a Curve (Null if another type)

	Surface (me) returns any Surface;
	---Purpose : returns Value as a Surface (Null if another type)


end GeometricSetSelect;

