-- Created on: 2002-12-12
-- Created by: data exchange team
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class AlignedCurve3dElementCoordinateSystem from StepFEA
inherits FeaRepresentationItem from StepFEA

    ---Purpose: Representation of STEP entity AlignedCurve3dElementCoordinateSystem

uses
    HAsciiString from TCollection,
    FeaAxis2Placement3d from StepFEA

is
    Create returns AlignedCurve3dElementCoordinateSystem from StepFEA;
	---Purpose: Empty constructor

    Init (me: mutable; aRepresentationItem_Name: HAsciiString from TCollection;
                       aCoordinateSystem: FeaAxis2Placement3d from StepFEA);
	---Purpose: Initialize all fields (own and inherited)

    CoordinateSystem (me) returns FeaAxis2Placement3d from StepFEA;
	---Purpose: Returns field CoordinateSystem
    SetCoordinateSystem (me: mutable; CoordinateSystem: FeaAxis2Placement3d from StepFEA);
	---Purpose: Set field CoordinateSystem

fields
    theCoordinateSystem: FeaAxis2Placement3d from StepFEA;

end AlignedCurve3dElementCoordinateSystem;
