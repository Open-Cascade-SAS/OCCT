-- File:	RWStepFEA_RWFeaShellMembraneStiffness.cdl
-- Created:	Thu Dec 12 17:51:06 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWFeaShellMembraneStiffness from RWStepFEA

    ---Purpose: Read & Write tool for FeaShellMembraneStiffness

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    FeaShellMembraneStiffness from StepFEA

is
    Create returns RWFeaShellMembraneStiffness from RWStepFEA;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : FeaShellMembraneStiffness from StepFEA);
	---Purpose: Reads FeaShellMembraneStiffness

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: FeaShellMembraneStiffness from StepFEA);
	---Purpose: Writes FeaShellMembraneStiffness

    Share (me; ent : FeaShellMembraneStiffness from StepFEA;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWFeaShellMembraneStiffness;
