-- Created on: 1993-05-05
-- Created by: Christian CAILLET
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class Protocol  from IGESData  inherits  Protocol from Interface

    ---Purpose : Description of basic Protocol for IGES
    --           This comprises treatement of IGESModel and Recognition of
    --           Undefined-FreeFormat-Entity

uses OStream, Type, InterfaceModel, Check

is

    Create returns mutable Protocol from IGESData;

    NbResources (me) returns Integer;
    ---Purpose : Gives the count of Resource Protocol. Here, none

    Resource (me; num : Integer) returns Protocol from Interface;
    ---Purpose : Returns a Resource, given a rank. Here, none

    TypeNumber (me; atype : any Type) returns Integer;
    ---Purpose : Returns a Case Number, specific of each recognized Type
    --         Here, Undefined and Free Format Entities have the Number 1.

    	-- --    General Services (defined at Norm level)    -- --

    NewModel (me) returns mutable InterfaceModel;
    ---Purpose : Creates an empty Model for IGES Norm

    IsSuitableModel (me; model : InterfaceModel) returns Boolean;
    ---Purpose : Returns True if <model> is a Model of IGES Norm

    UnknownEntity (me) returns mutable Transient;
    ---Purpose : Creates a new Unknown Entity for IGES (UndefinedEntity)

    IsUnknownEntity (me; ent : Transient) returns Boolean;
    ---Purpose : Returns True if <ent> is an Unknown Entity for the Norm, i.e.
    --           Type UndefinedEntity, status Unknown

end Protocol;
