-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class LocalTime from StepBasic 

inherits TShared from MMgt

uses

	Integer from Standard, 
	Real from Standard, 
	CoordinatedUniversalTimeOffset from StepBasic, 
	Boolean from Standard
is

	Create returns mutable LocalTime;
	---Purpose: Returns a LocalTime

	Init (me : mutable;
	      aHourComponent : Integer from Standard;
	      hasAminuteComponent : Boolean from Standard;
	      aMinuteComponent : Integer from Standard;
	      hasAsecondComponent : Boolean from Standard;
	      aSecondComponent : Real from Standard;
	      aZone : mutable CoordinatedUniversalTimeOffset from StepBasic) is virtual;

	-- Specific Methods for Field Data Access --

	SetHourComponent(me : mutable; aHourComponent : Integer);
	HourComponent (me) returns Integer;
	SetMinuteComponent(me : mutable; aMinuteComponent : Integer);
	UnSetMinuteComponent (me:mutable);
	MinuteComponent (me) returns Integer;
	HasMinuteComponent (me) returns Boolean;
	SetSecondComponent(me : mutable; aSecondComponent : Real);
	UnSetSecondComponent (me:mutable);
	SecondComponent (me) returns Real;
	HasSecondComponent (me) returns Boolean;
	SetZone(me : mutable; aZone : mutable CoordinatedUniversalTimeOffset);
	Zone (me) returns mutable CoordinatedUniversalTimeOffset;

fields

	hourComponent : Integer from Standard;
	minuteComponent : Integer from Standard;   -- OPTIONAL can be NULL
	secondComponent : Real from Standard;   -- OPTIONAL can be NULL
	zone : CoordinatedUniversalTimeOffset from StepBasic;
	hasMinuteComponent : Boolean from Standard;
	hasSecondComponent : Boolean from Standard;

end LocalTime;
