-- Created on: 1991-10-23
-- Created by: Denis PASCAL
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

generic class SortedStrgCmptsIterator from GraphTools
             (Graph      as any;
    	      Vertex     as any;
	      GIterator  as any;
	      SSCIterator as any)

--generic class SortedStrgCmptsIterator from GraphTools
--            (Graph     as any;
--    	       Vertex    as any;
--	       GIterator as GraphIterator  (Graph,Vertex))
--	       SSCIterator as  SortedStrgCmptsFromIterator

    ---Purposes: This     generic    class        implements       the
    --           SortedStrgCptsFromIterator  with all  vertices of <G>
    --           reached by the Tool GIterator.
     
raises NoMoreObject from Standard,
       NoSuchObject from Standard
    
is


    Create 
    returns SortedStrgCmptsIterator from GraphTools;
	---Purpose: Create an empty algorithm.
    
    Create (G : Graph) 	
    	---Purpose: Create the   algorithm setting each vertex  of <G>
	--          reached by  GIterator tool, as initial conditions.
	--          Use Perform   method before visting  the result of
	--          the algorithm.
    returns SortedStrgCmptsIterator from GraphTools;
    
    FromGraph (me : in out; G : Graph);	
    	---Purpose: Add each vertex of <G>  reached by GIterator  tool
	--          as   initial  conditions.   Use  Perform  method
	--          before   visiting the  result  of   the algorithm.
        ---Level: Public 
    
    FromVertex (me : in out; V : Vertex);	
    	---Purpose: Add  <V>  as  initial  condition.  This method  is
	--          cumulative.  Use Perform method before visting the
	--          result of the algorithm.  
	---Level: Public

    Reset (me : in out);	
    	---Purpose: Reset the algorithm.  It may   be reused with  new
    	--          initial conditions.  
        ---Level: Public

    Perform (me : in out; G : Graph);
       ---Purpose: Peform the  algorithm  in  <G> from initial  setted
       --          conditions.  
       ---Level: Public
    
    More(me) returns Boolean from Standard;
        ---Purpose: returns  True   if  there are   others  strong
        --          components.
       ---Level: Public

    Next(me : in out) 
        ---Purpose: Set the iterator to the next strong component.
       ---Level: Public
    raises NoMoreObject from Standard;

    NbVertices (me) returns Integer from Standard
	---Purpose: Returns number  of vertices of  the current Strong
	--          Components.
       ---Level: Public
    raises NoSuchObject from Standard;

    Value(me; I : Integer from Standard) 
    returns any Vertex
	---Purpose: returns  the vertex of  index <I> of  the  current
	--          Strong Component.
	---C++: return const &
       ---Level: Public
    raises NoSuchObject from Standard;

fields

    myIterator : SSCIterator;
    
end SortedStrgCmptsIterator;
















    
