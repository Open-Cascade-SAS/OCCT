-- Created on: 1997-07-28
-- Created by: Pierre CHALAMET
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Texture2Dmanual from Graphic3d

inherits Texture2D from Graphic3d

  ---Purpose: This class defined a manual texture 2D
  -- facets MUST define texture coordinate
  -- if you want to see somethings on.

uses

  NameOfTexture2D from Graphic3d,
  AsciiString     from TCollection,
  PixMap_Handle   from Image

is

  Create (theFileName : AsciiString from TCollection) returns mutable Texture2Dmanual from Graphic3d;
  ---Purpose: Creates a texture from a file

  Create (theNOT : NameOfTexture2D from Graphic3d) returns mutable Texture2Dmanual from Graphic3d;
  ---Purpose: Creates a texture from a predefined texture name set.

  Create (thePixMap : PixMap_Handle from Image) returns mutable Texture2Dmanual from Graphic3d;
  ---Purpose: Creates a texture from the pixmap.

end Texture2Dmanual;
