-- Created on: 1991-02-20
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package IntAna2d


    ---Purpose: This package defines the intersection between two elements of
    --          the geometric processor : Line, Circle, Ellipse, Parabola and
    --          Hyperbola; One of these elements is known with his real type,
    --          the other one is known by an implicit quadratic equation (see
    --          class Conic).
    --          A particular case has been made for the intersection between
    --          two Lin2d, two Circ2d, a Lin2d and a Circ2d.

uses

    Standard, TCollection, gp, StdFail

is

    class Conic;

    class AnaIntersection;

    class IntPoint;
     
end IntAna2d;
