-- Created on: 2003-10-21
-- Created by: Mikhail KLOKOV
-- Copyright (c) 2003-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class TrimShellCorner from BRepFill

uses
    Ax2    from  gp,
    Shape  from  TopoDS,
    Wire   from  TopoDS,
    Face   from  TopoDS,
    ListOfShape    from  TopTools,
    HArray2OfShape from  TopTools,
    DataMapOfShapeListOfShape  from  TopTools

is
    Create(theFaces         : HArray2OfShape from  TopTools;
    	   theAxeOfBisPlane : Ax2  from  gp;
    	   theSecPlane      : Face from TopoDS)
	 returns TrimShellCorner from BRepFill;

    Create(theFaces         : HArray2OfShape from  TopTools;
	   theAxeOfBisPlane :  Ax2  from  gp;
	   theSpine         :  Wire  from  TopoDS;
    	   theSecPlane      : Face from TopoDS)
	 returns TrimShellCorner from BRepFill;

    SetSpine(me: in out; theSpine:  Wire  from  TopoDS);

    AddBounds(me  :  in  out; Bounds : HArray2OfShape from  TopTools);

    AddUEdges(me  :  in  out; theUEdges : HArray2OfShape from  TopTools);

    Perform(me :  in  out);

    IsDone(me)  returns  Boolean from Standard; 
    
    HasSection(me)  returns  Boolean from Standard;

    Modified(me:in  out; S  :  Shape  from  TopoDS;
    	    	    	 theModified: out ListOfShape  from  TopTools);

fields
    myAxeOfBisPlane     : Ax2   from  gp;
    myShape1 : Shape from TopoDS;
    myShape2 : Shape from TopoDS;
    mySpine  : Wire from TopoDS;
    mySecPln : Face from TopoDS;
    myBounds : HArray2OfShape from  TopTools;
    myUEdges : HArray2OfShape from  TopTools;
    myFaces  : HArray2OfShape from  TopTools;
    myDone   : Boolean from Standard;
    myHasSection: Boolean from Standard;
    myHistMap:  DataMapOfShapeListOfShape  from  TopTools; 

end TrimShellCorner from BRepFill;
