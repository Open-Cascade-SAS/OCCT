--
-- File:	WNT_PixMap.cdl
-- Created:	27 October 1999
-- Author:	VKH
-- Updated:     SZV IMP100701 Add the "depth" field and method
--              to the pixmap object.
--
---Copyright:	MatraDatavision 1991,1992,1993

class PixMap from WNT

    ---Version:

    ---Purpose: This class defines a windows bitmap

    ---Keywords: Bitmap, Pixmap

inherits
    PixMap                from Aspect

uses
    Handle                from Aspect,
    Color                 from Quantity,
    Window                from Aspect

raises
    PixmapDefinitionError from Aspect,
    PixmapError           from Aspect

is

    Create ( aWindow          : Window from Aspect;
             aWidth, anHeight : Integer from Standard;
             aCDepth          : Integer from Standard = 0 )
    returns mutable PixMap from WNT
    raises PixmapDefinitionError from Aspect;
    ---Level: Public
    ---Purpose:  Warning! When <aDepth> is NULL , the pixmap is created
    -- with the SAME depth than the window <aWindow>

    ---------------------------------------------------
    -- Category: Methods to modify the class definition
    ---------------------------------------------------

    Destroy ( me : mutable )
    ---Level: Advanced
    ---Purpose: Destroies the Bitmap
    ---C++: alias ~
    --  Trigger: Raises if Bitmap is not defined properly
    raises PixmapError from Aspect is virtual;

    Dump ( me; aFilename : CString from Standard ;
           aGammaValue: Real from Standard = 1.0 )
    returns Boolean
    ---Level: Advanced
    ---Purpose:
    -- Dumps the Bitmap to an image file with
    -- an optional gamma correction value
    -- and returns TRUE if the dump occurs normaly.
    ---Category: Methods to modify the class definition
    raises PixmapError from Aspect is virtual;

    PixelColor ( me         : in;
                 theX, theY : in Integer from Standard )
    returns Color from Quantity
    is virtual;
    ---Purpose:
    -- Returns the pixel color.

    ----------------------------
    -- Category: Inquire methods
    ----------------------------

    PixmapID ( me ) returns Handle from Aspect is virtual;
    ---Level: Advanced
    ---Purpose: Returns the ID of the just created bitmap
    ---Category: Inquire methods

    ----------------------------
    -- Category: Private methods
    ----------------------------

    PreferedDepth( me ; aWindow: Window from Aspect;
                   aDepth: Integer from Standard)
    returns Integer from Standard is private;

fields
    myDC       : Handle from Aspect is protected;
    myBitmap   : Handle from Aspect is protected;
    myWND      : Window from Aspect;
end PixMap;
