-- Created on: 1994-05-24
-- Created by: Christian CAILLET
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ActorDispatch  from Transfer  inherits ActorOfTransientProcess

    ---Purpose : This class allows to work with a TransferDispatch, i.e. to
    --          transfer entities from a data set to another one defined by
    --          the same interface norm, with the following features :
    --          - ActorDispatch itself acts as a default actor, i.e. it copies
    --            entities with the general service Copy, as CopyTool does
    --          - it allows to add other actors for specific ways of transfer,
    --            which may include data modifications, conversions ...
    --          - and other features from TransferDispatch (such as mapping
    --            other than one-one)

uses Transient,        InterfaceModel,   GeneralLib, Protocol from Interface,
     TransferDispatch, TransientProcess, Binder

raises InterfaceError

is

    Create (amodel : InterfaceModel; lib : GeneralLib)
    	 returns ActorDispatch;
    ---Purpose : Creates an ActorDispatch from a Model. Works with a General
    --           Service Library, given as an Argument
    --           This causes TransferDispatch and its TransientProcess to be
    --           created, with default actor <me>

    Create (amodel : InterfaceModel; protocol : Protocol from Interface)
    	returns ActorDispatch;
    ---Purpose : Same as above, but Library is defined through a Protocol

    Create (amodel : InterfaceModel) returns ActorDispatch
    ---Purpose : Same as above, but works with the Active Protocol
    	raises InterfaceError;
    --           Error if no Active Protocol is defined

    AddActor (me : mutable; actor : ActorOfTransientProcess from Transfer);
    ---Purpose : Utility which adds an actor to the default <me> (it calls
    --           SetActor from the TransientProcess)

    TransferDispatch (me : mutable) returns TransferDispatch;
    ---Purpose : Returns the TransferDispatch, which does the work, records
    --           the intermediate data, etc...
    --           See TransferDispatch & CopyTool, to see the available methods
    ---C++ : return &


    Transfer (me : mutable; start : Transient; TP : TransientProcess)
    	returns Binder  is redefined;
    ---Purpose : Specific action : it calls the method Transfer from CopyTool
    --           i.e. the general service Copy, then returns the Binder
    --           produced by the TransientProcess

fields

    thetool : TransferDispatch;

end ActorDispatch;
