-- Created on: 1997-02-13
-- Created by: Alexander BRIVIN
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class TextureCoordinate2 from Vrml inherits  TShared  from  MMgt

	---Purpose:  defines a TextureCoordinate2 node of VRML specifying properties of geometry
	--  and its appearance.
	--  This  node  defines  a  set  of  2D  coordinates  to  be  used  to  map  textures 
	--  to  the  vertices  of  subsequent  PointSet,  IndexedLineSet,  or  IndexedFaceSet 
	--  objects.  It  replaces  the  current  texture  coordinates  in  the  rendering 
	--  state  for  the  shapes  to  use. 
	--  Texture  coordinates  range  from  0  to  1  across  the  texture. 
	--  The  horizontal  coordinate,  called  S,  is  specified  first,  followed   
	--  by  vertical  coordinate,  T.
    	--  By  default  : 
	--    myPoint (0 0)

uses
 
    HArray1OfVec2d  from TColgp 

is
    Create returns  mutable TextureCoordinate2 from Vrml; 

    Create  ( aPoint  :  HArray1OfVec2d   from  TColgp ) 
    	returns  mutable TextureCoordinate2 from Vrml; 
	  
    SetPoint ( me : mutable;  aPoint : HArray1OfVec2d   from  TColgp );
    Point ( me )  returns  HArray1OfVec2d   from  TColgp;

    Print  ( me;  anOStream: in out OStream from Standard) returns OStream from Standard;
    ---C++:  return  & 

fields
 
    myPoint  :  HArray1OfVec2d   from  TColgp;

end TextureCoordinate2;
