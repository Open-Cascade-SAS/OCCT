-- Created on: 1991-03-14
-- Created by: Laurent PAINNOT
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class BissecNewton from math
    	---Purpose:
    	-- This class implements a combination of Newton-Raphson and bissection 
    	--  methods to find the root of the function between two bounds.
        -- Knowledge of the derivative is required.

uses Vector from math, 
     Matrix from math, 
     FunctionWithDerivative from math,
     Status from math,
     OStream from Standard

raises NotDone from StdFail

is


    Perform(me: in out; F: out FunctionWithDerivative;
    	    Bound1, Bound2: Real;
	    NbIterations: Integer)

    is static protected;
    

    Create(F: in out FunctionWithDerivative;
    	   Bound1, Bound2, TolX: Real;
    	   NbIterations: Integer = 100)
    	---Purpose:
    	-- A combination of Newton-Raphson and bissection methods is done to find
    	-- the root of the function F between the bounds Bound1 and Bound2.
    	-- on the function F.
    	-- The tolerance required on the root is given by TolX.
    	-- The solution is found when :
    	--    abs(Xi - Xi-1) <= TolX and F(Xi) * F(Xi-1) <= 0
    	-- The maximum number of iterations allowed is given by NbIterations.

    returns BissecNewton;
    
    
    IsSolutionReached(me: in out; F: out FunctionWithDerivative)
    	---Purpose:    
    	-- This method is called at the end of each iteration to check if the
    	-- solution has been found.
    	-- It can be redefined in a sub-class to implement a specific test to
    	-- stop the iterations.

    returns Boolean
    is virtual;

    
    IsDone(me)
    	---Purpose: Tests is the root has been successfully found.
    	---C++: inline
    returns Boolean
    is static;
    
    
    Root(me)
       ---Purpose: returns the value of the root.
       -- Exception NotDone is raised if the minimum was not found.
       ---C++: inline
    returns Real
    raises NotDone
    is static;

    Derivative(me)
    	---Purpose: returns the value of the derivative at the root.
        -- Exception NotDone is raised if the minimum was not found.
    	---C++: inline

    returns Real
    raises NotDone
    is static;
    

    Value(me)
        ---Purpose: returns the value of the function at the root.
        -- Exception NotDone is raised if the minimum was not found.
    	---C++: inline

    returns Real
    raises NotDone
    is static;

    
    Dump(me; o: in out OStream)
    	---Purpose: Prints on the stream o information on the current state 
    	--          of the object.
    	--          Is used to redifine the operator <<.

    is static;


fields

Done:         Boolean;
TheStatus:    Status is protected;
XTol:         Real is protected;
x:            Real is protected;
dx:           Real is protected;
f:            Real is protected;
df:           Real is protected;

end BissecNewton;
