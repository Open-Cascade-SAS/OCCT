-- Created on: 1997-08-22
-- Created by: Prestataire Mary FABIEN
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class EdgeConnector from BRepAlgo inherits TShared from MMgt

    ---Purpose: Used by DSAccess to reconstruct an EdgeSet of connected edges. The result produced by
    --           MakeBlock is a list of non-standard TopoDS_wire,
    --          which  can present connexions of edge  of  order > 2 
    --           in certain  vertex. The method  IsWire
    --            indicates standard/non-standard character of  all wire produced.

uses

    ListOfShape    from TopTools,
    MapOfShape from TopTools,
    Shape from TopoDS,
    Edge from TopoDS,
    HDataStructure from TopOpeBRepDS,
    ShapeSet from TopOpeBRepBuild,
    BlockBuilder from TopOpeBRepBuild,
    DataMapOfShapeBoolean from BRepAlgo
    
is

    Create returns EdgeConnector from BRepAlgo;
    
    Add(me : mutable; e : Edge from TopoDS);
    ---Purpose: 
    
    Add(me : mutable; LOEdge : in out ListOfShape from TopTools);
    ---Purpose: 
    
    AddStart(me : mutable; e : Shape from TopoDS);
    ---Purpose: 
    
    AddStart(me : mutable; LOEdge : in out ListOfShape from TopTools);
    ---Purpose: 

    ClearStartElement(me : mutable);
    
    MakeBlock(me : mutable)
    ---Purpose: returns a list of wire non standard
    ---C++: return &
    returns ListOfShape from TopTools;
    
    Done(me : mutable);

    IsDone(me)
    ---Purpose: NYI
    ---Purpose: returns true if proceeded  to MakeBlock()
    returns Boolean from Standard;

    IsWire(me : mutable; W : Shape from TopoDS) 
    ---Purpose: NYI
    ---Purpose: returns true if W is  a Wire standard.
    --          W must belong  to the list returned  by MakeBlock.
    returns Boolean from Standard;

fields

    myListeOfEdge : ListOfShape from TopTools;
    myListeOfStartEdge : ListOfShape from TopTools;
    myResultMap : DataMapOfShapeBoolean from BRepAlgo;
    myResultList : ListOfShape from TopTools;
    myBlockB : BlockBuilder from TopOpeBRepBuild;
    myIsDone : Boolean from Standard;
    
end EdgeConnector from BRepAlgo;
