-- Created on: 2001-01-06
-- Created by: OCC Team
-- Copyright (c) 2001-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class Printer from Message inherits TShared from MMgt

  ---Purpose: Abstract interface class defining printer as output context for text messages
  --
  --          The message, besides being text string, has associated gravity
  --          level, which can be used by printer to decide either to process a message or ignore it.

uses

  Gravity from Message,
  AsciiString from TCollection,
  ExtendedString from TCollection

is

  Initialize returns Printer from Message;
  ---Purpose: Empty constructor with Message_Info trace level

  GetTraceLevel (me) returns Gravity from Message;
  ---C++: inline
  ---Purpose: Return trace level used for filtering messages;
  --          messages with lover gravity will be ignored.

  SetTraceLevel (me : mutable;
                 theTraceLevel : Gravity from Message);
  ---C++: inline
  ---Purpose: Set trace level used for filtering messages.
  --          By default, trace level is Message_Info, so that all messages are output

  Send (me;
        theString   : ExtendedString from TCollection;
        theGravity  : Gravity from Message;
        theToPutEol : Boolean) is deferred;
  ---Purpose: Send a string message with specified trace level.
  --          The parameter theToPutEol specified whether end-of-line should be added to the end of the message.
  --          This method must be redefined in descentant.

  Send (me;
        theString   : CString;
        theGravity  : Gravity from Message;
        theToPutEol : Boolean) is virtual;
  ---Purpose: Send a string message with specified trace level.
  --          The parameter theToPutEol specified whether end-of-line should be added to the end of the message.
  --          Default implementation calls first method Send().

  Send (me;
        theString   : AsciiString from TCollection;
        theGravity  : Gravity from Message;
        theToPutEol : Boolean) is virtual;
  ---Purpose: Send a string message with specified trace level.
  --          The parameter theToPutEol specified whether end-of-line should be added to the end of the message.
  --          Default implementation calls first method Send().

fields

  myTraceLevel : Gravity from Message is protected;

end Printer;
