-- Created on: 1998-07-27
-- Created by: Philippe MANGIN
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class EdgeOnSurfLaw from BRepFill inherits LocationLaw  from  BRepFill 

	---Purpose: Build Location Law, with a Wire and a  Surface.

uses
  Wire  from  TopoDS, 
  Shape  from TopoDS   

is 
    Create (Path   :  Wire  from  TopoDS; 
            Surf   :  Shape  from TopoDS)  
    returns EdgeOnSurfLaw  from BRepFill; 
     
     
    HasResult(me)   
	---Purpose: returns <False> if one  Edge of <Path> do not have
	--           representation on  <Surf>.   In this  case  it is
	--          impossible to use this object.          
    returns  Boolean; 
     
fields 
    hasresult  :  Boolean; 
    
end EdgeOnSurfLaw;
