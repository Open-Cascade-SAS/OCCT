-- Created on: 1993-12-02
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




generic class Iterator from Blend (Item as any)

	---Purpose: Template class for an iterator.
	--          A Sequence from TCollection can implement this iterator.

is

    Create

	---Purpose: Creates an empty iterator.

    	returns Iterator;


    Clear(me: in out);

	---Purpose: Clears the content of the iterator.



    Append(me: in out; I: Item);

	---Purpose: Adds an element in the iterator.


    Length(me: in out)
    
	---Purpose: Returns the number of elements in the iterator.

    	returns Integer;


    Value(me: in out; Index: Integer from Standard)
    
	---Purpose: Returns the element of range Index.
    
    	returns any Item;
	---C++: return const&
	---C++: alias operator()


end Iterator;
