-- File:	PDataStd_Axis.cdl
-- Created:	Wed Apr  9 13:43:28 1997
-- Author:	VAUTHIER Jean-Claude 
-- modified     Sergey Zaritchny
---Copyright:	 Matra Datavision 1997


class Axis from PDataXtd inherits Attribute from PDF

	---Purpose: 

is

    Create returns mutable Axis from  PDataXtd;
    
end Axis;
