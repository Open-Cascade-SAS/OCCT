-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Mat2d   from gp   inherits Storable
        ---Purpose:
        -- Describes a two column, two row matrix. This sort of
        -- object is used in various vectorial or matrix computations.
    
uses XY  from gp, 
     XYZ from gp

raises ConstructionError from Standard,
       OutOfRange        from Standard

is





  Create  returns Mat2d;
    	---C++: inline
        --- Purpose : Creates  a matrix with null coefficients.


  Create (Col1, Col2 : XY)   returns Mat2d;
        --- Purpose : 
        --  Col1, Col2 are the 2 columns of the matrix.



 

  SetCol (me : in out; Col : Integer; Value : XY)
        --- Purpose :  Assigns the two coordinates of Value to the column of range
        --   Col of this matrix 
        -- Raises OutOfRange if Col < 1 or Col > 2.
     raises OutOfRange
     is static;


  SetCols (me : in out; Col1, Col2 : XY)
        --- Purpose : Assigns the number pairs Col1, Col2 to the two columns of   this matrix
     is static;


  SetDiagonal (me : in out; X1, X2 : Real)     is static;
       ---C++: inline
       --- Purpose : 
       --  Modifies the main diagonal of the matrix.
       --  <me>.Value (1, 1) = X1
       --  <me>.Value (2, 2) = X2
       --  The other coefficients of the matrix are not modified.


  SetIdentity (me : in out)      is static;
    	---C++: inline
        --- Purpose : Modifies this matrix, so that it represents the Identity matrix.


  SetRotation (me : in out; Ang : Real)   is static;
        --- Purpose :
        --  Modifies this matrix, so that it representso a rotation. Ang is the angular
        --  value in radian of the rotation.
    	---C++: inline

  SetRow (me : in out; Row : Integer; Value : XY)
        --- Purpose : Assigns the two coordinates of Value to the row of index Row of this matrix. 
        -- Raises OutOfRange if Row < 1 or Row > 2.
     raises OutOfRange
     is static;


  SetRows (me : in out; Row1, Row2 : XY)    is static;
        --- Purpose : Assigns the number pairs Row1, Row2 to the two rows of this matrix.


  SetScale (me : in out; S : Real)    is static;
       ---C++: inline
       --- Purpose :
       --  Modifies the matrix such that it
       -- represents a scaling transformation, where S is the scale   factor :
       --           | S    0.0 |
       --   <me> =  | 0.0   S  |


  SetValue (me : in out; Row, Col : Integer; Value : Real)
        --- Purpose : Assigns <Value> to the coefficient of row Row, column Col of this matrix.
	-- Raises OutOfRange if Row < 1 or Row > 2 or Col < 1 or Col > 2
    	---C++: inline
     raises OutOfRange
     is static;

  Column (me; Col : Integer)   returns XY
        --- Purpose : Returns the column of Col index.
        -- Raises OutOfRange if Col < 1 or Col > 2
     raises OutOfRange
     is static;


  Determinant (me)   returns Real    is static;
    	---C++: inline
        --- Purpose : Computes the determinant of the matrix.


  Diagonal (me)  returns XY    is static;
        --- Purpose : Returns the main diagonal of the matrix.


  Row (me; Row : Integer)  returns XY
        --- Purpose : Returns the row of index Row.
     raises OutOfRange
        --- Purpose : Raised if Row < 1 or Row > 2
     is static;


  Value (me; Row, Col : Integer)  returns Real
        --- Purpose : Returns the coefficient of range (Row, Col)
	-- Raises OutOfRange
        -- if Row < 1 or Row > 2 or Col < 1 or Col > 2
	---C++: inline
    	---C++: return const &
    	---C++: alias operator()
     raises OutOfRange
       
     is static;


  ChangeValue (me : in out; Row, Col : Integer)  returns Real
        --- Purpose : Returns the coefficient of range (Row, Col)
     	-- Raises OutOfRange
        -- if Row < 1 or Row > 2 or Col < 1 or Col > 2
	---C++: inline
    	---C++: return  &
    	---C++: alias operator()
     raises OutOfRange
      
     is static;


  IsSingular (me)  returns Boolean   is static;
        --- Purpose :
    	-- Returns true if this matrix is singular (and therefore, cannot be inverted).
    	--  The Gauss LU decomposition is used to invert the matrix 
    	--  so the matrix is considered as singular if the largest 
    	--  pivot found is lower or equal to Resolution from gp.
    	---C++: inline


  Add (me : in out; Other : Mat2d)    is static;
    	---C++: inline
        ---C++: alias operator +=

  Added (me; Other : Mat2d)  returns Mat2d   is static;
        ---C++: inline
        ---C++: alias operator +

        --- Purpose :
        --  Computes the sum of this matrix and the matrix
    	-- Other.for each coefficient of the matrix :
        --  <me>.Coef(i,j) + <Other>.Coef(i,j)
    	-- Note:
    	-- -   operator += assigns the result to this matrix, while
    	-- -   operator + creates a new one.
    	
    

  Divide (me : in out; Scalar : Real)    is static;
        ---C++: inline
        ---C++: alias operator /=

  Divided (me; Scalar : Real)  returns Mat2d   is static;
    	---C++: inline
        ---C++: alias operator /
	    --- Purpose : 
	    --  Divides all the coefficients of the matrix by a scalar.



  Invert (me : in out)  raises ConstructionError   is static;

  Inverted (me)  returns Mat2d   raises ConstructionError   is static;
        --- Purpose :
        --  Inverses the matrix and raises exception if the matrix
        --  is singular.
    	---C++: inline

     

  Multiplied (me; Other : Mat2d)   returns Mat2d   is static;
    	  ---C++: inline
          ---C++: alias operator *

  Multiply (me : in out; Other : Mat2d)            is static;
       --- Purpose :
       --  Computes the product of two matrices <me> * <Other>
       ---C++: inline
       -- C++: alias operator *=

  PreMultiply(me : in out; Other : Mat2d)          is static;
       --- Purpose : Modifies this matrix by premultiplying it by the matrix Other
       -- <me> = Other * <me>.
       ---C++: inline

          
    
  Multiplied (me; Scalar : Real)   returns Mat2d   is static;
    	---C++: inline
        ---C++: alias operator *

  Multiply (me : in out; Scalar : Real)    is static;
        --- Purpose :
        --  Multiplies all the coefficients of the matrix by a scalar.
    	---C++: inline
        ---C++: alias operator *=


  Power (me : in out; N : Integer)  raises ConstructionError is static;

  Powered (me; N : Integer)  returns Mat2d  raises ConstructionError is static;
    	--- Purpose :
        --  computes <me> = <me> * <me> * .......* <me>, N time.
        --  if N = 0 <me> = Identity
        --  if N < 0 <me> = <me>.Invert() *...........* <me>.Invert().
        --  If N < 0 an exception can be raised if the matrix is not
        --  inversible
    	---C++: inline

  
  Subtract (me : in out; Other : Mat2d)           is static;
    	---C++: inline
        ---C++: alias operator -=

  Subtracted (me; Other : Mat2d)  returns Mat2d   is static;
    	---C++: inline
        ---C++: alias operator -
        --- Purpose :
        --  Computes for each coefficient of the matrix :
        --  <me>.Coef(i,j) - <Other>.Coef(i,j)


  Transpose (me : in out)        is static;
    	---C++: inline  

  Transposed (me)  returns Mat2d is static;
        --- Purpose : 
        --  Transposes the matrix. A(j, i) -> A (i, j)
        ---C++: inline
fields

  matrix : Real[2, 2];

friends

  class Trsf2d   from gp,
  class GTrsf2d  from gp,
  class XY       from gp

end;
