-- Created on: 1993-06-16
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class ShapeSet from BOP

    ---Purpose:  
    
    -- Auxiliary class providing an exploration of a set
    -- of shapes to build faces or solids. 
    
    -- To build faces  : shapes are wires, elements are edges.
    -- To build solids : shapes are shells, elements are faces. 
    
    -- The ShapeSet stores a list of shapes, a list of elements
    -- to start reconstructions, and a map to search neighbours.
    -- The map stores the connection  between elements through 
    -- subshapes of type <SubShapeType> given in constructor.  
    
    -- <SubShapeType> is :
    --  - TopAbs_VERTEX to connect edges
    --  - TopAbs_EDGE to connect faces
    --
 	
uses

    ShapeEnum     from TopAbs, 
    
    Orientation   from TopAbs,
    Shape         from TopoDS,
     
    ListOfShape                      from TopTools,
    ListIteratorOfListOfShape        from TopTools,
    IndexedDataMapOfShapeListOfShape from TopTools,
    IndexedMapOfOrientedShape        from TopTools,
     
    Explorer from TopExp

is

    Create (SubShapeType  :  ShapeEnum from TopAbs)
    	 returns ShapeSet from BOP;
    	---Purpose:  
    	--- Creates a ShapeSet  in order to build shapes connected
    	--- by <SubShapeType>  shapes. 
    	---

    Delete(me:out)  
    	is virtual;
    	---C++: alias "Standard_EXPORT virtual ~BOP_ShapeSet(){Delete() ; }"
    	---Purpose:  
    	--- Destructor 
    	---
    AddShape(me:out; 
    	    S:Shape from TopoDS)  
    	is virtual;
    	---Purpose:  
    	--- Adds <S> to the list of shapes. (wires or shells).
    	---
    AddStartElement(me:out; 
    	    S:Shape from TopoDS)  
    	is virtual;
    	---Purpose:  
    	--- Add S to the list of starting shapes used for reconstructions.
    	--- apply AddElement(S).
    	---
    AddElement(me:out; 
    	    S:Shape from TopoDS)  
    	is virtual;
    	---Purpose: 
    	--- For each subshape SE of S of type mySubShapeType
    	--- Add subshapes of S to the map of subshapes (mySubShapeMap)
    	--- Add S to the list of shape incident to subshapes of S.
    	---
    ProcessAddShape(me:out; 
    	    S:Shape from TopoDS)  
    	is static protected;
    	---Purpose: 
    	--- Internal  purpose
    	---
    ProcessAddStartElement(me:out; 
    	    S:Shape from TopoDS)  
    	is static protected;
    	---Purpose: 
    	--- Internal  purpose
    	---
    ProcessAddElement(me:out; 
    	    S:Shape from TopoDS)  
    	is static protected;
    	---Purpose: 
    	--- Internal  purpose
    	---
    StartElements(me)  
    	returns ListOfShape from TopTools;
	---C++: return const & 
    	---Purpose:  
    	--- Selector. 
	---
    --
    --
    -- Iteration on the shapes of AddShape()
    -- 
    InitShapes(me:out); 
    	---Purpose: 
    	--- Internal  purpose
    	---
    MoreShapes(me)  
    	returns Boolean from Standard; 
    	---Purpose: 
    	--- Internal  purpose
    	---
    NextShape(me:in out); 
    	---Purpose: 
    	--- Internal  purpose
    	---
    Shape(me)  
    	returns Shape from TopoDS;
    	---C++: return const &

    --
    -- Iteration on the start elements of AddStartElement()
    -- 
    InitStartElements(me:out); 
    	
    MoreStartElements(me)  
    	returns Boolean from Standard; 
    	---Purpose: 
    	--- Internal  purpose
    	---
    NextStartElement(me:out);
    	---Purpose: 
    	--- Internal  purpose
    	---
    StartElement(me)  
    	returns Shape;
    	---C++: return const &
    	---Purpose: 
    	--- Iteration on the neighbours of a shape of type myShapeType
    	--- through its subshapes of type mySubShapeType. 
    	---
    InitNeighbours(me:out; 
    	    S:Shape from TopoDS)  
    	is virtual;
     
    MoreNeighbours(me:out)  
    	returns Boolean from Standard;
    	---Purpose: 
    	--- Internal  purpose
    	---
    NextNeighbour(me: out);
    	---Purpose: 
    	--- Internal  purpose
    	---
    Neighbour(me)  
    	returns Shape from TopoDS;
    	---C++: return const & 
    	---Purpose: 
    	--- Internal  purpose
    	---
    ChangeStartShapes(me:out)  
    	returns ListOfShape from TopTools;
    	---C++: return &
    	---Purpose: 
    	--- Modifier 
    	---

    FindNeighbours(me:in out)  
    	is virtual;
    	---Purpose: 
    	--- Build the list of neighbour shapes of myCurrentShape
    	--- (neighbour shapes and myCurrentShapes are of type t)
    	--- Initialize myIncidentShapesIter on neighbour shapes.
	---
   
    MakeNeighboursList(me:in out;E,V:Shape)  
    	returns ListOfShape from TopTools  
    	is virtual;
    	---C++: return const &
    
    MaxNumberSubShape(me:in out;Shape:Shape)  
    	returns Integer; 


    ClearContents(me:out);
    	---Purpose:  
    	--- Clears myStartShapes,mySubShapeMap,myShapes   
    	---
fields

    myShapeType : ShapeEnum from TopAbs is protected;  
    -- shape type : edge

    mySubShapeType : ShapeEnum from TopAbs is protected;
    -- subshape type : vertex
    
    --mySubShapeExplorer : ShapeExplorer from BOP is protected;
    mySubShapeExplorer : Explorer from TopExp is protected;
    -- explorer of edge vertices

    myStartShapes : ListOfShape from TopTools is protected;
    -- list of starting edges

    myStartShapesIter : ListIteratorOfListOfShape from TopTools is protected; 
    -- myStartShapes iterator

    mySubShapeMap : IndexedDataMapOfShapeListOfShape from TopTools is protected;
    -- map of vertices
    -- mySubShapeMap(vertex) = list of incident edges to a vertex

    myIncidentShapesIter : ListIteratorOfListOfShape from TopTools is protected;
    -- iter on list L of edges incident to a vertex, L = mySubShapeMap(vertex)

    myShapes : ListOfShape from TopTools is protected;
    -- list of wires which are not to be reconstructed
	
    myShapesIter : ListIteratorOfListOfShape from TopTools is protected;
    -- myShapes iterator

    myCurrentShape : Shape from TopoDS is protected;
    -- current edge which neighbours are searched, using FindNeighbours()
	
    myCurrentShapeNeighbours : ListOfShape from TopTools is protected;
    -- list of edges neighbour of the edge myCurrentShape

end ShapeSet;
