-- Created on: 1997-02-11
-- Created by: Alexander BRIVIN and Dmitry TARASOV
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class ShapeHints from Vrml 

	---Purpose: defines a ShapeHints node of VRML specifying properties of geometry and its appearance.
    	--  The ShapeHints node indicates that IndexedFaceSets are solid, contain ordered vertices, or
	--  contain convex faces. 
	--  These hints allow VRML implementations to optimize certain rendering features.
       	--  Optimizations that may be performed include enabling back-face culling and disabling
       	--  two-sided lighting. For example, if an object is solid and has ordered vertices, an
       	--  implementation may turn on backface culling and turn off two-sided lighting. To ensure
       	--  that an IndexedFaceSet can be viewed from either direction, set shapeType to be
       	--  UNKNOWN_SHAPE_TYPE. 
	--  If you know that your shapes are closed and will alwsys be viewed from the outside, set
       	--  vertexOrdering to be either CLOCKWISE or COUNTERCLOCKWISE (depending on
       	--  how you built your object), and set shapeType to be SOLID. Placing this near the top of
       	--  your VRML file will allow the scene to be rendered much faster.  
       	--  The ShapeHints node also affects how default normals are generated. When an
       	--  IndexedFaceSet has to generate default normals, it uses the creaseAngle field to determine
       	--  which edges should be smoothly shaded and which ones should have a sharp crease. The
       	--  crease angle is the angle between surface normals on adjacent polygons. For example, a
       	--  crease angle of .5 radians (the default value) means that an edge between two adjacent
       	--  polygonal faces will be smooth shaded if the normals to the two faces form an angle that is
       	--  less than .5 radians (about 30 degrees). Otherwise, it will be faceted. 
uses
 
    VertexOrdering from  Vrml, 
    ShapeType      from  Vrml, 
    FaceType       from  Vrml

is
    Create  ( aVertexOrdering : VertexOrdering from  Vrml = Vrml_UNKNOWN_ORDERING; 
    	      aShapeType      : ShapeType      from  Vrml = Vrml_UNKNOWN_SHAPE_TYPE;
    	      aFaceType       : FaceType       from  Vrml = Vrml_CONVEX; 
	      aAngle          : Real           from  Standard  =  0.5  ) 
	  returns ShapeHints from Vrml;
	     
    SetVertexOrdering ( me : in out;  
           aVertexOrdering : VertexOrdering from Vrml ); 
    VertexOrdering ( me )  returns  VertexOrdering from Vrml; 

    SetShapeType ( me : in out; aShapeType  :  ShapeType  from  Vrml  );
    ShapeType ( me ) returns  ShapeType  from  Vrml;

    SetFaceType ( me : in out; aFaceType  : FaceType  from  Vrml ); 
    FaceType ( me ) returns  FaceType  from  Vrml; 

    SetAngle  ( me : in out; aAngle  :  Real from Standard );
    Angle  ( me ) returns  Real from Standard;

    Print  ( me;  anOStream: in out OStream from Standard) returns OStream from Standard;
    ---C++:  return  & 
 
fields
 
    myVertexOrdering  :  VertexOrdering  from  Vrml;     -- Ordering of face vertices
    myShapeType       :  ShapeType       from  Vrml;     -- Info about shape geometry
    myFaceType        :  FaceType        from  Vrml;     -- Info about face geometry
    myAngle           :  Real            from  Standard; -- Smallest angle for sharp edge
    
end ShapeHints;
