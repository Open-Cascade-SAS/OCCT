-- Created on: 1998-02-23
-- Created by: Christian CAILLET
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class TypedValue  from Interface    inherits TypedValue  from MoniTool

    ---Purpose : Now strictly equivalent to TypedValue from MoniTool,
    --           except for ParamType which remains for compatibility reasons
    --           
    --           This class allows to dynamically manage .. typed values, i.e.
    --           values which have an alphanumeric expression, but with
    --           controls. Such as "must be an Integer" or "Enumerative Text"
    --           etc
    --           
    --           Hence, a TypedValue brings a specification (type + constraints
    --           if any) and a value. Its basic form is a string, it can be
    --           specified as integer or real or enumerative string, then
    --           queried as such.
    --           Its string content, which is a Handle(HAsciiString) can be
    --           shared by other data structures, hence gives a direct on line
    --           access to its value.

uses CString, Type from Standard,
     AsciiString from TCollection, HAsciiString from TCollection,
     HSequenceOfAsciiString  from TColStd, HArray1OfAsciiString  from TColStd,
     HSequenceOfHAsciiString from TColStd,
     DictionaryOfInteger from Dico,
     ParamType from Interface , ValueType from MoniTool,
     ValueSatisfies from Interface, ValueInterpret from Interface

raises InterfaceError

is

    Create (name : CString;
    	    type : ParamType from Interface = Interface_ParamText;
	    init : CString = "")  returns mutable TypedValue;
    ---Purpose : Creates a TypedValue, with a name
    --           
    --           type gives the type of the parameter, default is free text
    --           Also available : Integer, Real, Enum, Entity (i.e. Object)
    --           More precise specifications, titles, can be given to the
    --           TypedValue once created
    --           
    --           init gives an initial value. If it is not given, the
    --           TypedValue begins as "not set", its value is empty

    Type   (me) returns ParamType from Interface;
    ---Purpose : Returns the type
    --           I.E. calls ValueType then makes correspondance between
    --             ParamType from Interface (which remains for compatibility
    --              reasons) and ValueType from MoniTool

    ParamTypeToValueType (myclass; typ : ParamType from Interface)
    	returns ValueType from MoniTool;
    ---Purpose : Correspondance ParamType from Interface  to
    --               ValueType from MoniTool

    ValueTypeToParamType (myclass; typ : ValueType from MoniTool)
    	returns ParamType from Interface;
    ---Purpose : Correspondance ParamType from Interface  to
    --               ValueType from MoniTool

fields

    thename   : AsciiString;
    thedef    : AsciiString;
    thelabel  : AsciiString;
    thetype   : ParamType from Interface;
    theotyp   : Type from Standard;  -- for object

    thelims   : Integer;  -- status for integer/enum/real limits
    themaxlen : Integer;
    theintlow : Integer;
    theintup  : Integer;
    therealow : Real;
    therealup : Real;
    theunidef : AsciiString;

    theenums  : HArray1OfAsciiString    from TColStd;
    theeadds  : DictionaryOfInteger;

    theinterp : ValueInterpret;
    thesatisf : ValueSatisfies;
    thesatisn : AsciiString;

    theival   : Integer;
    thehval   : HAsciiString from TCollection;
    theoval   : Transient;

end Static;
