-- Created on: 1993-01-09
-- Created by: CKY / Contract Toubro-Larsen ( TCD )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class HighLight from IGESGraph  inherits IGESEntity

        ---Purpose: defines IGESHighLight, Type <406> Form <20>
        --          in package IGESGraph
        --
        --          Attaches information that an entity is to be
        --          displayed in some system dependent manner

uses  Integer  -- no one specific type


is

        Create returns mutable HighLight;

        -- Specific Methods pertaining to the class

        Init (me               : mutable;
              nbProps          : Integer;
              aHighLightStatus : Integer);
        ---Purpose : This method is used to set the fields of the class
        --           HighLight
        --      - nbProps          : Number of property values (NP = 1)
        --      - aHighLightStatus : HighLight Flag

        NbPropertyValues(me) returns Integer;
        ---Purpose : returns the number of property values in <me>

        HighLightStatus(me) returns Integer;
        ---Purpose : returns 0 if <me> is not highlighted(default),
        --         1 if <me> is highlighted

        IsHighLighted(me) returns Boolean;
        ---Purpose : returns True if entity is highlighted

fields

--
-- Class    : IGESGraph_HighLight
--
-- Purpose  : Declaration of the variables specific to a
--            HighLight property.
--
-- Reminder : A HighLight property is defined by :
--                  - Number of property values (NP=1)
--                  - Flag
--

        theNbPropertyValues : Integer;

        theHighLight        : Integer;

end HighLight;
