-- Created on: 2000-12-25
-- Created by: Igor FEOKTISTOV <ifv@nnov.matra-dtv.fr>
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Intersection from QANewModTopOpe   
    inherits BooleanOperation from BRepAlgoAPI 
 
---Purpose: provides  intersection  of  two  shapes;
 
uses

    Shape from TopoDS, 
    DataMapOfShapeListOfShape from TopTools,
    ListOfShape from TopTools
     
is 
  
    Create(theObject1,  theObject2 : Shape from TopoDS )
    ---Purpose: 
    
    returns Intersection  from QANewModTopOpe;   

    Generated (me: in out; theS : Shape from TopoDS)
    	---Purpose: Returns the list  of shapes generated from the shape <S>. 
        ---C++: return const & 
        ---Level: Public
    returns ListOfShape from TopTools
    is redefined; 

    HasGenerated (me)
    	returns Boolean from Standard
	is redefined;
    	---Purpose: Returns true if there is at least one generated shape.
    	---         For use in BRepNaming.

    IsDeleted (me: in out;  
    	    aS : Shape from TopoDS)
    	returns Boolean
    	is redefined;


    HasDeleted (me)
    	returns Boolean from Standard
	is redefined;
    	---Purpose: Returns true if there is at least one deleted shape.
    	---         For use in BRepNaming.

fields
    
    myMapGener: DataMapOfShapeListOfShape from TopTools;

end  Intersection;
