-- Created on: 1993-01-09
-- Created by: CKY / Contract Toubro-Larsen ( SIVA )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class SelectedComponent from IGESSolid  inherits IGESEntity

        ---Purpose: defines SelectedComponent, Type <182> Form Number <0>
        --          in package IGESSolid
        --          The Selected Component entity provides a means of
        --          selecting one component of a disjoint CSG solid

uses

        BooleanTree     from IGESSolid,
        XYZ             from gp,
        Pnt             from gp

is

        Create returns mutable SelectedComponent;

        -- Specific Methods pertaining to the class

        Init (me        : mutable;
              anEntity  : BooleanTree;
              selectPnt : XYZ);
        ---Purpose : This method is used to set the fields of the class
        --           SelectedComponent
        --       - anEntity  : the Boolean tree entity
        --       - selectPnt : Point in or on the desired component

        Component(me) returns BooleanTree;
        ---Purpose : returns the Boolean tree entity

        SelectPoint(me) returns Pnt;
        ---Purpose : returns the point on/in the selected component

        TransformedSelectPoint(me) returns Pnt;
        ---Purpose : returns the point on/in the selected component
        -- after applying TransformationMatrix

fields

--
-- Class    : IGESSolid_SelectedComponent
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class SelectedComponent.
--
-- Reminder : A SelectedComponent instance is defined by :
--            a pointer to the Boolean Tree entity(Entity) and the X, Y
--            and Z components (X,Y,Z) of a selected point.

        theEntity      : BooleanTree;
            -- the desired boolean tree entity

        theSelectPoint : XYZ;
            -- the X, Y and Z coordinates of the point

end SelectedComponent;
