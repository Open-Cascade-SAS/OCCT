-- Created on: 1994-11-14
-- Created by: Jean Claude VAUTHIER 
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package StlTransfer 

	---Purpose: The  package   Algorithm  for Meshing   implements
	--          facilities to compute  the Mesh data-structure, as
	--          defined in package StlMesh, from a shape of package
	--          TopoDS.  The triangulation  is  computed  with the
	--          Delaunay      algorithm   implemented in   package
	--          BRepMesh.  The  result   is  stored  in  the  mesh
	--          data-structure Mesh from package StlMesh.
	--          

uses  

    StlMesh,
    TopoDS

is
    BuildIncrementalMesh (Shape      : in      Shape from TopoDS; 
    	       	    	  Deflection : in      Real  from Standard;
    	       	    	  InParallel : in      Boolean from Standard;
    	       	          Mesh       : Mesh  from StlMesh)
     raises ConstructionError;
end StlTransfer;






