-- File:	PTopoDS_Compound.cdl
-- Created:	Wed May  5 16:57:51 1993
-- Author:	Remi LEQUETTE
--		<rle@sdsun1>
---Copyright:	 Matra Datavision 1993



class Compound from PTopoDS inherits HShape from PTopoDS

is
    Create returns mutable Compound from PTopoDS;
	---Level: Internal 

end Compound;
