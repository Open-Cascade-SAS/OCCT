-- File:	BRepFeat_MakePipe.cdl
-- Created:	Tue Sep  3 11:13:22 1996
-- Author:	Olga PILLOT
--		<jag@mobilox.lyon.matra-dtv.fr>
---Copyright:	 Matra Datavision 1996




class MakeDPrism from BRepFeat inherits Form from BRepFeat

	---Purpose: Describes functions to build draft
    	-- prism topologies from basis shape surfaces. These can be depressions or protrusions.
    	-- The semantics of draft prism feature creation is based on the
    	-- construction of shapes:
    	-- -          along a length
    	-- -          up to a limiting face
    	-- -          from a limiting face to a height.
    	-- The shape defining construction of the draft prism feature can be
    	-- either the supporting edge or the concerned area of a face.
    	-- In case of the supporting edge, this contour can be attached to a
    	-- face of the basis shape by binding. When the contour is bound to this
    	-- face, the information that the contour will slide on the face
    	-- becomes available to the relevant class methods.
    	-- In case of the concerned area of a face, you could, for example, cut
    	-- it out and move it to a different height which will define the
    	-- limiting face of a protrusion or depression.

uses Shape                     from TopoDS,
     Face                      from TopoDS,
     Wire                      from TopoDS,
     Edge                      from TopoDS,
     DataMapOfShapeListOfShape from TopTools,
     DataMapOfShapeShape       from TopTools,
     SequenceOfCurve           from TColGeom,
     Curve                     from Geom,
     ListOfShape               from TopTools,
     StatusError               from BRepFeat

raises ConstructionError from Standard

is


    Create(Sbase     : Shape   from TopoDS;
           Pbase     : Face    from TopoDS;
           Skface    : Face    from TopoDS;
           Angle     : Real    from Standard;
           Fuse      : Integer from Standard;
           Modify    : Boolean from Standard)

	   
	---Purpose: A face Pbase is selected in the shape
    	--   Sbase to serve as the basis for the draft prism. The
    	--   draft will be defined by the angle Angle and Fuse offers a choice between:
    	-- - removing matter with a Boolean cut using the setting 0
    	-- - adding matter with Boolean fusion using the setting 1.
    	--    The sketch face Skface serves to determine the type of
    	-- operation. If it is inside the basis shape, a local
    	-- operation such as glueing can be performed.
    		---C++: inline
    	    	returns MakeDPrism from BRepFeat;

    Create
	---Purpose: Initializes the draft prism class
    		---C++: inline
    	    	returns MakeDPrism from BRepFeat;




    Init(me: in out; Sbase     : Shape   from TopoDS;
 		     Pbase     : Face    from TopoDS;
                     Skface    : Face    from TopoDS;
                     Angle     : Real    from Standard;
                     Fuse      : Integer from Standard;
                     Modify    : Boolean from Standard)
    	is static;
    	---Purpose: Initializes this algorithm for building draft prisms along surfaces.
    	-- A face Pbase is selected in the basis shape Sbase to
    	-- serve as the basis from the draft prism. The draft will be
    	-- defined by the angle Angle and Fuse offers a choice between:
    	-- -   removing matter with a Boolean cut using the setting 0
    	-- -   adding matter with Boolean fusion using the setting  1.
    	--   The sketch face Skface serves to determine the type of
    	-- operation. If it is inside the basis shape, a local
    	-- operation such as glueing can be performed.

    Add(me: in out; E: Edge from TopoDS; OnFace: Face from TopoDS)

	---Purpose: Indicates that the edge <E> will slide on the face
	--          <OnFace>. 
    	-- Raises ConstructionError if the  face does not belong to the
	-- basis shape, or the edge to the prismed shape.
    	raises ConstructionError from Standard
	
	is static;


    Perform(me: in out; Height: Real from Standard)
     
    	is static;


    Perform(me: in out; Until: Shape from TopoDS)
    
    	is static;


    Perform(me: in out; From : Shape from TopoDS;
                        Until: Shape from TopoDS)
    
    	is static;
    	---Purpose: Assigns one of the following semantics
    	-- -   to a height Height
    	-- -   to a face Until
    	-- -   from a face From to a height Until.
    	-- Reconstructs the feature topologically according to the semantic option chosen.
    
    PerformUntilEnd(me: in out)
    	---Purpose: Realizes a semi-infinite prism, limited by the position of the prism base.   
    	is static;

    PerformFromEnd(me: in out; FUntil: Shape from TopoDS)
    	---Purpose: Realizes a semi-infinite prism, limited by the face Funtil. 
    	is static;

    PerformThruAll(me: in out)
    	---Purpose: Builds an infinite prism. The infinite descendants will not be kept in the result.    
    	is static;

    PerformUntilHeight(me: in out; Until :  Shape from TopoDS;
                        Height:  Real  from Standard)
    	---Purpose: Assigns both a limiting shape, Until from
    	-- TopoDS_Shape, and a height, Height at which to stop
    	-- generation of the prism feature.    
    	is static;


    Curves(me: in out; S : in out SequenceOfCurve from TColGeom);
    

    BarycCurve(me: in out)    
    	returns Curve from Geom;
	
	
    BossEdges(me: in out; sig: Integer from Standard)
        ---Purpose: Determination of TopEdges and LatEdges.
        --          sig = 1 -> TopEdges = FirstShape of the DPrism
        --          sig = 2 -> TOpEdges = LastShape of the DPrism
	is static;

	
    TopEdges(me: in out)
        ---Purpose: Returns the list of TopoDS Edges of the top of the boss.
    returns ListOfShape from TopTools
	---C++: return const&
    	is static;


    LatEdges(me: in out)
        ---Purpose: Returns the list of TopoDS Edges of the bottom of the boss.
    returns ListOfShape from TopTools
	---C++: return const&
    	is static;


fields

    myPbase  : Face                      from TopoDS;
    mySlface : DataMapOfShapeListOfShape from TopTools;
    myAngle  : Real                      from Standard;
    myCurves : SequenceOfCurve           from TColGeom;
    myBCurve : Curve                     from Geom;    
    myTopEdges    : ListOfShape          from TopTools;
    myLatEdges    : ListOfShape          from TopTools; 
    myStatusError : StatusError          from BRepFeat;

end MakeDPrism;




