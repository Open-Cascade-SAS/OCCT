-- Created on: 1999-04-08
-- Created by: Fabrice SERVANT
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Couple from IntPolyh
 

uses
    
    Pnt from gp


is


    Create;
    
    Create(i1,i2: Integer from Standard) ; 
    
    FirstValue(me) 
    returns Integer from Standard
    is static;

    SecondValue(me) 
    returns Integer from Standard
    is static;
    
    AnalyseFlagValue(me)
    returns Integer from Standard
    is static;

    AngleValue(me)
    returns Real from Standard
    is static;

    SetCoupleValue(me: in out; v,w: Integer from Standard) 
    is static;
	
    SetAnalyseFlag(me: in out; v: Integer from Standard) 
    is static;
    
    SetAngleValue(me: in out; ang: Real from Standard) 
    is static;
	
    Dump(me; v: Integer from Standard) 
    is static;
     	
fields

    t1,t2,ia : Integer from Standard;
    angle : Real from Standard;
    
end Couple from IntPolyh;
