-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class AreaInSet from StepVisual 

inherits TShared from MMgt

uses

	PresentationArea from StepVisual, 
	PresentationSet from StepVisual
is

	Create returns mutable AreaInSet;
	---Purpose: Returns a AreaInSet

	Init (me : mutable;
	      aArea : mutable PresentationArea from StepVisual;
	      aInSet : mutable PresentationSet from StepVisual) is virtual;

	-- Specific Methods for Field Data Access --

	SetArea(me : mutable; aArea : mutable PresentationArea);
	Area (me) returns mutable PresentationArea;
	SetInSet(me : mutable; aInSet : mutable PresentationSet);
	InSet (me) returns mutable PresentationSet;

fields

	area : PresentationArea from StepVisual;
	inSet : PresentationSet from StepVisual;

end AreaInSet;
