-- Created on: 1996-08-30
-- Created by: Xavier BENVENISTE
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class Interpolate from GeomLib

	---Purpose: this class is used to construct a BSpline curve by
	--          interpolation  of points  at given parameters  The
	--          continuity   of the curve   is degree -  1 and the
	--          method used when boundary  condition are not given
	--          is to use odd degrees  and null the derivatives on
	--          both sides from degree -1 down to (degree+1) / 2
	--          When even degree is given the returned curve is of
	--          degree - 1 so that the degree of the curve is odd 
    	

uses
    Array1OfPnt         from TColgp,
    Array1OfReal        from TColStd,
    InterpolationErrors from GeomLib,
    BSplineCurve        from Geom

raises

    NotDone    from StdFail,
    OutOfRange from Standard
    
is

    Create( Degree     : Integer from Standard ;
    	    NumPoints  : Integer from Standard ;
	    Points     : Array1OfPnt from TColgp ;
	    Parameters : Array1OfReal from TColStd) 
	     
    returns Interpolate from GeomLib ;
    
    IsDone(me) returns Boolean from Standard
    	---Purpose: 
    	-- returns if everything went OK
	---C++: inline
    is static;


    Error(me) returns InterpolationErrors from GeomLib 
    ---Purpose: returns the error type if any 
    ---C++: inline	      
    --          
    is static ;

    Curve(me) 
    ---Purpose:  returns the interpolated curve of the requested degree 

    returns BSplineCurve from Geom
    raises
    	OutOfRange from Standard,
	NotDone    from StdFail
    is static;
 
    
    
fields

    myCurve : BSplineCurve from Geom ;
    myIsDone : Boolean from Standard ;
    myError  : InterpolationErrors  from GeomLib  ;
    
end Interpolate ;

