-- Created on: 2018-03-15
-- Created by: Stephan GARNAUD (ARM)
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.





class Printer from OSD 

 ---Purpose: Selects a printer.

uses Error, AsciiString from TCollection
raises ConstructionError, NullObject, OSDError

is
  Create (Name : AsciiString) returns Printer
   ---Purpose: Initializes printer to use with its name.
   --          The string must contain only ASCII characters
   --          between ' ' and '~'; this means no control character 
   --          and no extended ASCII code. If it is not the case the
   --          exception ConstructionError is raised.
   ---Level: Advanced
  raises ConstructionError;

  SetName (me : in out; Name : AsciiString)
  ---Purpose: Changes name of printer to use.
  ---Level: Advanced
  raises ConstructionError, NullObject is static;

  Name (me ;Name : out AsciiString) is static;
  ---Purpose: Returns name of current printer
  ---Level: Advanced

 Failed (me) returns Boolean is static;
  ---Purpose: Returns TRUE if an error occurs
  ---Level: Advanced

 Reset (me : in out) is static;
  ---Purpose: Resets error counter to zero
  ---Level: Advanced
      
 Perror (me : in out) 
  ---Level: Advanced
  ---Purpose: Raises OSD_Error
   raises OSDError is static;

 Error (me) returns Integer is static;
  ---Purpose: Returns error number if 'Failed' is TRUE.
  ---Level: Advanced

fields

  myName  : AsciiString;
  myError : Error;
end Printer from OSD;


