-- Created on: 1992-11-05
-- Created by: Remi LEQUETTE
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Cone from BRepPrim inherits Revolution from BRepPrim

	---Purpose: Implement the cone primitive.

uses
    Face from TopoDS,

    Pnt from gp,
    Ax2 from gp    

raises
    DomainError

is

    Create(Angle : Real; Position : Ax2 from gp; Height : Real;
    	       Radius : Real = 0)
    returns Cone from BRepPrim
	   ---Purpose: the STEP definition
	   --          Angle = semi-angle of the cone
	   --          Position : the coordinate system
	   --          Height : height of the cone.
	   --          Radius : radius of truncated face at z = 0
	   --          
	   --          The apex is on z < 0
	   --          
	   --          Errors : Height < Resolution
	   --                    Angle < Resolution / Height
	   --                    Angle > PI/2 - Resolution / Height
    raises DomainError;

    Create(Angle : Real)
    returns Cone from BRepPrim
	---Purpose: infinite cone at origin on Z negative
    raises DomainError;
    
    Create(Angle : Real; Apex : Pnt from gp)
    returns Cone from BRepPrim
	---Purpose: infinite cone at Apex on Z negative
    raises DomainError;
    
    Create(Angle : Real; Axes : Ax2 from gp)
    returns Cone from BRepPrim
	---Purpose: infinite cone with Axes
    raises DomainError;
    
    Create(R1,R2,H : Real)
    returns Cone from BRepPrim
	---Purpose: create a  Cone at origin  on Z axis, of height  H,
	--          radius R1 at Z = 0, R2 at  Z = H, X is  the origin
	--          of angles.  If R1 or  R2 is 0   there is  an apex.
	--          Otherwise, it is a truncated cone.
	--          
	--          Error  : R1 and R2  < Resolution
	--                   R1 or R2 negative
	--                   Abs(R1-R2) < Resolution
	--                   H < Resolution
	--                   H negative
    raises DomainError;
    
    Create(Center : Pnt from gp; R1,R2,H : Real)
    returns Cone from BRepPrim
	---Purpose: same as above but at a given point
    raises DomainError;
    
    Create(Axes : Ax2 from gp; R1,R2,H : Real)
    returns Cone from BRepPrim
	---Purpose: same as above with given axes system.
    raises DomainError;
    
    MakeEmptyLateralFace(me) returns Face from TopoDS
	---Purpose: The surface normal should be directed  towards the
	--          outside.
    is redefined;
    
    SetMeridian(me : in out)
    is static private;
    
    SetParameters(me : in out; R1, R2, H : Real)
    is static private;
    
fields
    myHalfAngle : Real;
    myRadius    : Real;

end Cone;
