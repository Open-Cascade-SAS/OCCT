-- Created on: 1994-04-05
-- Created by: Yves FRICAUD
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

private class FunctionH from Bisector 

inherits FunctionWithDerivative from math
     
             --                                  2           2 
	---Purpose: H(v) = (T1  .P2(v) - P1) * ||T(v)||  -
	--                                  2         2
	--                 (T(v).P2(v) - P1) * ||T1|| 
	
uses 
    Curve from Geom2d,
    Pnt2d from gp, 
    Vec2d from gp  

is

    Create (C2 : Curve from Geom2d ;
            P1 : Pnt2d from gp     ;
            T1   : Vec2d from gp   ) 
    returns FunctionH from Bisector;
    
    Value(me : in out; X : Real; F : out Real) 
    	---Purpose: Computes the values of the Functions for the variable <X>.
    returns Boolean;
    
    Derivative(me : in out; X : Real; D : out Real) 
    returns Boolean;

    Values(me : in out ; X  : Real; F  : out Real; D  : out Real)    
    	---Purpose: Returns the values of the functions and the derivatives
    	--          for the variable <X>.
    returns Boolean;

fields
    
    curve2 : Curve from Geom2d;
    p1     : Pnt2d from gp;
    t1     : Vec2d from gp;
    
end FunctionH;
