-- Created on: 1997-07-28
-- Created by: Pierre CHALAMET
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

class Texture1Dsegment from Graphic3d

inherits Texture1D from Graphic3d

  ---Purpose:  This class provides the implementation
  -- of a 1D texture applyable along a segment.
  -- You might use the SetSegment() method
  -- to set the way the texture is "streched" on facets.

uses

  NameOfTexture1D from Graphic3d,
  AsciiString     from TCollection

is

  Create (theFileName : AsciiString from TCollection) returns mutable Texture1Dsegment from Graphic3d;
  ---Purpose: Creates a texture from a file

  Create (theNOT : NameOfTexture1D from Graphic3d) returns mutable Texture1Dsegment from Graphic3d;
  ---Purpose: Creates a texture from a predefined texture name set.

  SetSegment (me : mutable;
              theX1, theY1, theZ1 : ShortReal from Standard;
              theX2, theY2, theZ2 : ShortReal from Standard);
  ---Purpose: Sets the texture application bounds. Defines the way
  -- the texture is stretched across facets.
  -- Default values are <0.0, 0.0, 0.0> , <0.0, 0.0, 1.0>

  --
  -- inquire methods
  --
  Segment (me;
           theX1, theY1, theZ1 : out ShortReal from Standard;
           theX2, theY2, theZ2 : out ShortReal from Standard);
  ---Purpose: Returns the values of the current segment X1, Y1, Z1 , X2, Y2, Z2.

fields

  myX1, myY1, myZ1 : ShortReal from Standard;
  myX2, myY2, myZ2 : ShortReal from Standard;
      
end  Texture1Dsegment;
