-- Created on: 1992-11-04
-- Created by: Gilles DEBARBOUILLE
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




private class ShiftedUnit from Units  

inherits

    Unit from Units

	---Purpose: This class is useful   to describe  units  with  a
	--          shifted origin in relation to another unit. A well
	--          known example  is the  Celsius degrees in relation
	--          to Kelvin degrees. The shift of the Celsius origin
	--          is 273.15 Kelvin degrees.


uses

    Quantity from Units,
    Token from Units

is

    Create(aname , asymbol : CString ;
           avalue , amove : Real ;
           aquantity : Quantity from Units)
    
    ---Level: Internal 
    
    ---Purpose: Creates  and  returns a  shifted unit.   <aname> is the
    --          name of the unit,  <asymbol> is the usual abbreviation
    --          of the unit, <avalue> is the  value in relation to the
    --          International System of Units, and <amove>  is the gap
    --          in relation to another unit.
    --          
    --          For  example Celcius   dregee   of temperature  is  an
    --          instance of ShiftedUnit  with <avalue> equal to 1. and
    --          <amove> equal to 273.15.
    
    returns mutable ShiftedUnit from Units;
    
    Create(aname , asymbol : CString)
    
    ---Level: Internal 
    
    ---Purpose: Creates  and returns a  unit.  <aname> is  the name of
    --          the  unit, <asymbol> is the  usual abbreviation of the
    --          unit.
    
    returns mutable ShiftedUnit from Units;
    
    Create(aname : CString)
    
    ---Level: Internal 
    
    ---Purpose: Creates  and returns a  unit.  <aname> is  the name of
    --          the  unit.
    
    returns mutable ShiftedUnit from Units;
    
    Move(me : mutable ; amove : Real)
    
    ---Level: Internal 
    
    ---Purpose: Sets the field <themove> to <amove>
    
    is static;
    
    Move(me) returns Real
    
    ---Level: Internal 
    
    ---Purpose: Returns the shifted value <themove>.
    
    is static;
    
    Token(me) returns mutable Token from Units
    
    ---Level: Internal 
    
    ---Purpose: This redefined method returns a ShiftedToken object.
    
    is redefined;
    
    Dump(me ; ashift , alevel : Integer)
    
    ---Level: Internal 
    
    is redefined;

fields

    themove : Real;

end ShiftedUnit;
