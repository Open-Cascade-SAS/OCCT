-- File:	RWStepShape_RWCompoundShapeRepresentation.cdl
-- Created:	Fri Dec 28 16:01:59 2001 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class RWCompoundShapeRepresentation from RWStepShape

    ---Purpose: Read & Write tool for CompoundShapeRepresentation

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    CompoundShapeRepresentation from StepShape

is
    Create returns RWCompoundShapeRepresentation from RWStepShape;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : CompoundShapeRepresentation from StepShape);
	---Purpose: Reads CompoundShapeRepresentation

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: CompoundShapeRepresentation from StepShape);
	---Purpose: Writes CompoundShapeRepresentation

    Share (me; ent : CompoundShapeRepresentation from StepShape;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWCompoundShapeRepresentation;
