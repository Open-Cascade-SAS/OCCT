-- File:	BOPTest_DrawableShape.cdl
-- Created:	Thu May 25 14:55:46 2000
-- Author:	Peter KURNEV
--		<pkv@irinox>
---Copyright:	 Matra Datavision 2000


class DrawableShape from BOPTest inherits DrawableShape from DBRep

    ---Purpose: 

uses  

    Shape           from TopoDS,
    Color           from Draw,
    Display         from Draw,
    Text3D          from Draw,
    Marker3D        from Draw,
    CString         from Standard,
    Pnt             from gp

is

    Create (S         : Shape from TopoDS;
    	    FreeCol   : Color from Draw;    -- color for free edges
    	    ConnCol   : Color from Draw;    -- color for shared edges
	    EdgeCol   : Color from Draw;    -- color for other edges
	    IsosCol   : Color from Draw;    -- color for Isos
	    size      : Real;               -- size for infinite isos
	    nbisos    : Integer;            -- # of isos on each face
	    discret   : Integer;            -- # of points on curves
    	    Text      : CString from Standard; 
    	    TextColor : Color from Draw
    	    )
    	returns mutable DrawableShape from BOPTest;

    Create (S         : Shape from TopoDS;
    	    Text      : CString from Standard; 
    	    TextColor : Color from Draw
    	    )
    	returns mutable DrawableShape from BOPTest; 
	
    Pnt(me) returns Pnt from gp  is private;
  
    DrawOn(me; dis : in out Display from Draw)
    is redefined;
    
fields

    myText : Text3D from Draw;
    myTextColor : Color from Draw;

end DrawableShape;
