-- Created on: 1996-12-16
-- Created by: Remi Lequette
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Iterator from TNaming 

	---Purpose: A tool to visit the contents of a named shape attribute.
    	-- Pairs of shapes in the attribute are iterated, one
    	-- being the pre-modification or the old shape, and
    	-- the other the post-modification or the new shape.
    	-- This allows you to have a full access to all
    	-- contents of an attribute. If, on the other hand, you
    	-- are only interested in topological entities stored
    	-- in the attribute, you can use the functions
    	-- GetShape and CurrentShape in TNaming_Tool.

uses

    Label       from TDF,
    Evolution   from TNaming,
    NamedShape  from TNaming,	
    PtrNode     from TNaming,
    Shape       from TopoDS

raises

    NoMoreObject from Standard,
    NoSuchObject from Standard 

is

    Create( anAtt  : NamedShape from TNaming) returns Iterator from TNaming;
	---Purpose: Iterates on all  the history records in
	--          <anAtt>.
    
    Create( aLabel : Label from TDF) returns Iterator from TNaming;
	---Purpose: Iterates on all  the history records in
	--          the current transaction

    Create( aLabel : Label from TDF; aTrans : Integer from Standard)
    returns Iterator from TNaming;
	---Purpose: Iterates on all  the history records in
	--          the transaction <aTrans>
	
    More(me) returns Boolean;
	---C++: inline
	---Purpose: Returns True if there is a current Item in
	--          the iteration.
     
    Next(me : in out)
    	---Purpose: Moves the iteration to the next Item 
    raises
	NoMoreObject from Standard;
   
    OldShape(me) returns Shape from TopoDS
    	---Purpose: Returns the old shape in this iterator object.
    	-- This shape can be a null one.
	---C++: return const&
    raises
	NoSuchObject from Standard;
	 
    NewShape(me) returns Shape from TopoDS
    	---Purpose: Returns the new shape in this iterator object.
 	---C++: return const&
   raises
	 NoSuchObject from Standard;
	 
    IsModification(me) returns Boolean;
	---Purpose: Returns true if the  new  shape is a modification  (split,
	--          fuse,etc...) of the old shape.
	--          
    
    Evolution(me) returns Evolution from TNaming;
    

fields

    myNode  : PtrNode from TNaming;
    myTrans : Integer from Standard;  -- is < 0 means in Current Transaction.

friends
    
    class NewShapeIterator from TNaming,
    class OldShapeIterator from TNaming    
    
end Iterator;
