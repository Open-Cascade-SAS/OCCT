-- Created on: 1993-07-06
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MakeEdge from BRepLib  inherits MakeShape from BRepLib

	---Purpose: Provides methods to build edges.
	--          
	--          The   methods have  the  following   syntax, where
	--          TheCurve is one of Lin, Circ, ...
	--          
	--          Create(C : TheCurve)
	--            
	--            Makes an edge on  the whole curve.  Add vertices
	--            on finite curves.
	--            
	--          Create(C : TheCurve; p1,p2 : Real)
	--          
	--            Make an edge  on the curve between parameters p1
	--            and p2. if p2 < p1 the edge will be REVERSED. If
	--            p1  or p2 is infinite the  curve will be open in
	--            that  direction. Vertices are created for finite
	--            values of p1 and p2.
	--            
	--          Create(C : TheCurve; P1, P2 : Pnt from gp)
	--          
	--            Make an edge on the curve  between the points P1
	--            and P2. The  points are projected on   the curve
	--            and the   previous method is  used. An  error is
	--            raised if the points are not on the curve.
	--            
	--          Create(C : TheCurve; V1, V2 : Vertex from TopoDS)
	--          
	--            Make an edge  on the curve  between the vertices
	--            V1 and V2. Same as the  previous but no vertices
	--            are created. If a vertex is  Null the curve will
	--            be open in this direction.

uses
    EdgeError from BRepLib,
    Edge   from TopoDS,
    Vertex from TopoDS,
    Pnt    from gp,
    Lin    from gp,
    Circ   from gp,
    Elips  from gp,
    Hypr   from gp,
    Parab  from gp,
    Curve  from Geom2d,
    Curve  from Geom,
    Surface from Geom
    
raises
    NotDone from StdFail
    
is

    Create returns MakeEdge from BRepLib;
    
    ----------------------------------------
    -- Points
    ----------------------------------------

    Create(V1, V2 : Vertex from TopoDS)                    
	---Level: Public
    returns MakeEdge from BRepLib;

    Create(P1, P2 : Pnt from gp)                           
	---Level: Public
    returns MakeEdge from BRepLib;


    ----------------------------------------
    -- Lin
    ----------------------------------------
	
    Create(L : Lin from gp)                                
	---Level: Public
    returns MakeEdge from BRepLib;

    Create(L : Lin from gp; p1,p2 : Real)                  
	---Level: Public
    returns MakeEdge from BRepLib;

    Create(L : Lin from gp; P1,P2 : Pnt from gp)           
	---Level: Public
    returns MakeEdge from BRepLib;

    Create(L : Lin from gp; V1, V2 : Vertex from TopoDS)   
	---Level: Public
    returns MakeEdge from BRepLib;

    ----------------------------------------
    -- Circ
    ----------------------------------------
	
    Create(L : Circ from gp)                               
	---Level: Public
    returns MakeEdge from BRepLib;

    Create(L : Circ from gp; p1,p2 : Real)                 
	---Level: Public
    returns MakeEdge from BRepLib;

    Create(L : Circ from gp; P1,P2 : Pnt from gp)          
	---Level: Public
    returns MakeEdge from BRepLib;

    Create(L : Circ from gp; V1, V2 : Vertex from TopoDS)  
	---Level: Public
    returns MakeEdge from BRepLib;

	
    ----------------------------------------
    -- Elips
    ----------------------------------------

    Create(L : Elips from gp)                               
	---Level: Public
    returns MakeEdge from BRepLib;

    Create(L : Elips from gp; p1,p2 : Real)                 
	---Level: Public
    returns MakeEdge from BRepLib;

    Create(L : Elips from gp; P1,P2 : Pnt from gp)          
	---Level: Public
    returns MakeEdge from BRepLib;

    Create(L : Elips from gp; V1, V2 : Vertex from TopoDS)  
	---Level: Public
    returns MakeEdge from BRepLib;

    ----------------------------------------
    -- Hypr
    ----------------------------------------

    Create(L : Hypr from gp)                               
	---Level: Public
    returns MakeEdge from BRepLib;

    Create(L : Hypr from gp; p1,p2 : Real)                 
	---Level: Public
    returns MakeEdge from BRepLib;

    Create(L : Hypr from gp; P1,P2 : Pnt from gp)          
	---Level: Public
    returns MakeEdge from BRepLib;

    Create(L : Hypr from gp; V1, V2 : Vertex from TopoDS)  
	---Level: Public
    returns MakeEdge from BRepLib;

    ----------------------------------------
    -- Parab
    ----------------------------------------

    Create(L : Parab from gp)                               
	---Level: Public
    returns MakeEdge from BRepLib;

    Create(L : Parab from gp; p1,p2 : Real)                 
	---Level: Public
    returns MakeEdge from BRepLib;

    Create(L : Parab from gp; P1,P2 : Pnt from gp)          
	---Level: Public
    returns MakeEdge from BRepLib;

    Create(L : Parab from gp; V1, V2 : Vertex from TopoDS)  
	---Level: Public
    returns MakeEdge from BRepLib;

    ----------------------------------------
    -- Curve
    ----------------------------------------

    Create(L : Curve from Geom)                               
	---Level: Public
    returns MakeEdge from BRepLib;

    Create(L : Curve from Geom; p1,p2 : Real)                 
	---Level: Public
    returns MakeEdge from BRepLib;

    Create(L : Curve from Geom; 
    P1,P2 : Pnt from gp)
	---Level: Public                        
    returns MakeEdge from BRepLib;

    Create(L : Curve from Geom; 
    V1, V2 : Vertex from TopoDS)
	---Level: Public
    returns MakeEdge from BRepLib;

    Create(L : Curve from Geom; 
    P1,P2 : Pnt from gp; p1,p2 : Real)                        
	---Level: Public
    returns MakeEdge from BRepLib;

    Create(L : Curve from Geom; 
    V1, V2 : Vertex from TopoDS;
    p1, p2 :Real)       
	---Level: Public                                      
    returns MakeEdge from BRepLib;

    ----------------------------------------
    -- Curve and surface
    ----------------------------------------

    Create(L : Curve from Geom2d; S : Surface from Geom)
    	---Level: Public
    returns MakeEdge from BRepLib;

    Create(L : Curve from Geom2d; S : Surface from Geom; p1,p2 : Real)
    	---Level: Public
    returns MakeEdge from BRepLib;

    Create(L : Curve from Geom2d; S : Surface from Geom; 
    P1,P2 : Pnt from gp)
	---Level: Public                        
    returns MakeEdge from BRepLib;

    Create(L : Curve from Geom2d; S : Surface from Geom; 
    V1, V2 : Vertex from TopoDS)
	---Level: Public
    returns MakeEdge from BRepLib;

    Create(L : Curve from Geom2d; S : Surface from Geom; 
    P1,P2 : Pnt from gp; p1,p2 : Real)                        
	---Level: Public
    returns MakeEdge from BRepLib;

    Create(L : Curve from Geom2d; S : Surface from Geom; 
    V1, V2 : Vertex from TopoDS;
    p1, p2 :Real)       
	---Level: Public                                      
    returns MakeEdge from BRepLib;

    ----------------------------------------
    --  Auxiliary methods
    ----------------------------------------

    Init(me : in out; C      : Curve from Geom)
	---Level: Public
    is static;
    
    Init(me : in out; C      : Curve from Geom;
		      p1, p2 : Real)
	---Level: Public
    is static;		      
	
    Init(me : in out; C      : Curve from Geom;
    	    	      P1, P2 : Pnt   from gp)
	---Level: Public
    is static;		      
	
    Init(me : in out; C      : Curve  from Geom;
    	              V1, V2 : Vertex from TopoDS)
	---Level: Public
    is static;
	
    Init(me : in out; C      : Curve from Geom;
    	    	      P1, P2 : Pnt   from gp;
		      p1, p2 : Real)
	---Level: Public
    is static;		      
	
    Init(me : in out; C      : Curve  from Geom;
    	              V1, V2 : Vertex from TopoDS;
		      p1, p2 : Real)
	---Level: Public
    is static;
	
    Init(me : in out; C      : Curve from Geom2d; S : Surface from Geom)
	---Level: Public
    is static;
    
    Init(me : in out; C      : Curve from Geom2d; S : Surface from Geom;
		      p1, p2 : Real)
	---Level: Public
    is static;		      
	
    Init(me : in out; C      : Curve from Geom2d; S : Surface from Geom;
    	    	      P1, P2 : Pnt   from gp)
	---Level: Public
    is static;		      
	
    Init(me : in out; C      : Curve  from Geom2d; S : Surface from Geom;
    	              V1, V2 : Vertex from TopoDS)
	---Level: Public
    is static;
	
    Init(me : in out; C      : Curve from Geom2d; S : Surface from Geom;
    	    	      P1, P2 : Pnt   from gp;
		      p1, p2 : Real)
	---Level: Public
    is static;		      
	
    Init(me : in out; C      : Curve  from Geom2d; S : Surface from Geom;
    	              V1, V2 : Vertex from TopoDS;
		      p1, p2 : Real)
	---Level: Public
    is static;
	

    ----------------------------------------
    --  Results
    ----------------------------------------

    Error(me) returns EdgeError from BRepLib
	---Purpose: Returns the error description when NotDone.
	---Level: Public
    is static;

    Edge(me) returns Edge from TopoDS
	---C++: return const &
	---C++: alias "Standard_EXPORT operator TopoDS_Edge() const;"
	---Level: Public
    raises
    	NotDone from StdFail
    is static;
    
    Vertex1(me) returns Vertex from TopoDS
	---Purpose: Returns the first vertex of the edge. May be Null.
	--          
	---C++: return const &
	---Level: Public
    is static;
    
    Vertex2(me) returns Vertex from TopoDS
	---Purpose: Returns the second vertex of the edge. May be Null.
	--          
	---C++: return const &
	---Level: Public
    is static; 
    
fields

    myError   : EdgeError from BRepLib;
    myVertex1 : Vertex    from TopoDS;
    myVertex2 : Vertex    from TopoDS;

end MakeEdge;
