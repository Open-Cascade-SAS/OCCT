-- Created on: 1994-11-04
-- Created by: Frederic MAUPAS
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MakeTrimmedCurve2d from StepToGeom

    ---Purpose: This class implements the mapping between classes 
    --          class TrimmedCurve from StepGeom which
    --          describes a Trimmed Curve from prostep and TrimmedCurve from 
    --          Geom. 
  
uses BSplineCurve from Geom2d,
     TrimmedCurve from StepGeom

is 

    Convert ( myclass; SC : TrimmedCurve from StepGeom;
                       CC : out BSplineCurve from Geom2d )
    returns Boolean from Standard;

end MakeTrimmedCurve2d;
