-- Created on: 1997-09-11
-- Created by: Philippe MANGIN
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class LinearCriteria from AppDef inherits SmoothCriterion from AppDef

	---Purpose: defined an Linear Criteria to used in variational
	--          Smoothing of points.


uses
   Vector  from  math, 
   Matrix  from  math, 
   Curve   from  FEmTool, 
   HAssemblyTable    from  FEmTool, 
   ElementaryCriterion  from  FEmTool,   
   HArray2OfInteger  from TColStd, 
   HArray1OfReal     from TColStd,
   Array1OfReal      from TColStd,
   MultiLine         from AppDef,
   MyLineTool        from AppDef
   
raises 
  NotImplemented,   
  DomainError 
   
 

is 
    Create(SSP: MultiLine from AppDef; 
    	   FirstPoint, LastPoint: Integer)  returns  LinearCriteria;

    SetParameters(me  :  mutable;  Parameters  : HArray1OfReal); 

    SetCurve(me  :  mutable;  C  :Curve from FEmTool) 
    is  static; 
     
    GetCurve(me;  C  :  out  Curve  from FEmTool) 
    is  static; 
     
    SetEstimation(me  :  mutable;  E1,  E2,  E3  :  Real)   
    is  static; 

    EstLength(me  :  mutable)   
    ---C++: return &
    returns  Real  is  static;      
      
    GetEstimation(me;  E1,  E2,  E3  : out Real)   
    is  static; 
     
    AssemblyTable(me)  
    returns HAssemblyTable  from  FEmTool   
    is  static; 
     
    DependenceTable(me)  
    returns  HArray2OfInteger  from TColStd   
    is  static;  
    
     
    QualityValues  (me : mutable; J1min,  J2min,  J3min  :  Real; 
    	    	    	    	  J1,  J2,  J3  :  out  Real) 
				 returns  Integer  is  static; 

    ErrorValues(me  :  mutable;   
                MaxError,  QuadraticError,  AverageError  :  out  Real) 
    is  static;
     
    Hessian(me  :  mutable ;  
            Element    :  Integer; 
	    Dimension1  :  Integer; 
	    Dimension2  :  Integer;
            H  :  out  Matrix  from  math)  
     raises  DomainError -- If DependenceTable(Dimension1,Dimension2) is False 
     is  static;  
   
    
    Gradient(me  :  mutable;  
             Element  :  Integer; 
	     Dimension  :  Integer;
             G  :  out  Vector  from  math) 
    is  static; 
    
    InputVector(me  :  mutable;  X : Vector from math;   
                                 AssTable : HAssemblyTable  from  FEmTool)  
    ---Purpose: Convert the assembly Vector in an Curve;
    --          
    raises  DomainError; 
     
    SetWeight(me:  mutable;  
              QuadraticWeight,  QualityWeight  :  Real; 
	      percentJ1,  percentJ2,  percentJ3  :  Real) 
    is  static; 
     
    GetWeight(me;  QuadraticWeight,  QualityWeight  :  out  Real)  
    is  static;  
    
    SetWeight(me:  mutable;  
              Weight  :  Array1OfReal)
    is  static; 
     
    BuildCache(me:  mutable;  E  :  Integer)  is  private;
          
fields
mySSP         :  MultiLine from AppDef; 
myParameters  :  HArray1OfReal; 
myCache     :    HArray1OfReal;
myCriteria  :  ElementaryCriterion  from  FEmTool[3]; 
myEstimation:  Real[3];  
myQuadraticWeight,  myQualityWeight  :  Real; 
myPercent   :  Real[3]; 
myPntWeight :  Array1OfReal;
myCurve     :  Curve  from  FEmTool; 
myLength    :  Real;  
myE         :  Integer; 
IF,  IL     :  Integer;
end LinearCriteria;


