-- Created on: 1997-05-06
-- Created by: Yves FRICAUD
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

private class IteratorOnShapesSet from TNaming 

	---Purpose: 

uses
    ShapesSet               from TNaming,
    Shape                   from TopoDS,
    MapIteratorOfMapOfShape from TopTools
    
raises
    NoMoreObject from Standard,
    NoSuchObject from Standard

is
    Create returns IteratorOnShapesSet;
         ---C++: inline

    Create (S : ShapesSet from TNaming) returns IteratorOnShapesSet;    	
    	 ---C++: inline
    
    Init (me : in out; S : ShapesSet from TNaming);
	---Purpose: Initialize the iteration
    	---C++: inline
    
    More (me) returns Boolean;
	---Purpose: Returns True if there is a current Item in
	--          the iteration.
    	---C++: inline
    
    Next (me : in out)
    	---Purpose: Move to the next Item 
    	---C++: inline
    raises
	NoMoreObject from Standard;
    
    Value(me) returns Shape from TopoDS
    	---C++: return const&
    raises
	NoSuchObject from Standard;


fields
    myIt    : MapIteratorOfMapOfShape from TopTools;

end IteratorOnShapesSet;
