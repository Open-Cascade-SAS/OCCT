-- Created on: 1995-01-25
-- Created by: Jean-Louis Frenkel
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Modified by Rob : 20-feb-1997
-- Modified by Rob : 16-dec-1997 : kind of presentation

deferred class Presentation from PrsMgr
inherits TShared  from MMgt

uses 

    PresentationManager from PrsMgr,
    KindOfPrs from PrsMgr

is

    Initialize(aPresentationManager: PresentationManager from PrsMgr)
    is protected;

    KindOfPresentation(me) returns KindOfPrs from PrsMgr is deferred;    
    ---Purpose: 2D or 3D
    
    Display(me: mutable) is deferred private;
    
    Erase(me: mutable) is deferred private;

    SetVisible (me: mutable; theValue: Boolean from Standard) is deferred private;

    Highlight(me: mutable) is deferred private;
    
    Unhighlight (me) is deferred private;
    
    IsHighlighted(me) returns Boolean from Standard
    is deferred private;

    IsDisplayed(me) returns Boolean from Standard
    is deferred private;

    Destroy ( me : mutable )
    is virtual; 
    ---Level: Public    
    ---Purpose: Destructor
    ---C++:     alias ~

    DisplayPriority(me) returns Integer from Standard
    is deferred private;
    
    SetDisplayPriority(me:mutable;aNewPrior:Integer from Standard)
    is deferred private;

    SetZLayer ( me : mutable;
                theLayerId : Integer from Standard )
      is deferred private;
    ---Purpose: Set Z layer ID for the presentation

    GetZLayer ( me )
      returns Integer from Standard is deferred private;
    ---Purpose: Get Z layer ID for the presentation

    Clear(me: mutable) 
    is deferred private;
    
---Category: Inquire Methods
--            
    PresentationManager(me) returns mutable PresentationManager
    ---Purpose: returns the PresentationManager in which the
    --          presentation has been created.
    is static;
    ---C++: inline
    ---C++: return const&


---Category: Internal Methods

    SetUpdateStatus(me:mutable; aStat : Boolean from Standard);
    ---C++: inline
    
    MustBeUpdated(me) returns Boolean from Standard;
    ---C++: inline


fields

    myPresentationManager: PresentationManager from PrsMgr is protected;
    myMustBeUpdated      : Boolean from Standard is protected;

friends
    class PresentationManager from PrsMgr
        
end Presentation from PrsMgr;
