-- Created on: 1997-08-07
-- Created by: Jean-Louis Frenkel
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Directory from CDF inherits Transient from Standard


---Purpose: A directory is a collection of documents. There is only one instance
--          of a given document in a directory.
--          put.

uses Document from CDM, ListOfDocument from CDM

raises  NoSuchObject
    
is
    Create 
    returns mutable Directory from CDF;
    ---Purpose: Creates an empty directory.
    
    
    Add(me:mutable; aDocument: Document from CDM);
    ---Purpose: adds a document into the directory.
    
    Remove(me: mutable; aDocument: Document from CDM);
    ---Purpose: removes the document.
    
    
---Category: Inquire Methods
--           

    Contains(me; aDocument: Document from CDM) 
    ---Purpose: Returns true if the document aDocument is in the directory
    returns Boolean from Standard
    is static;

    Last(me:mutable) returns Document from CDM
    ---Purpose: returns the last document (if any) which has been added
    --          in the directory.
    raises NoSuchObject from Standard
    ---Warning: if the directory is empty.
    is static;

    Length(me) returns Integer from Standard
    ---Purpose: returns the number of documents of the directory.
    is static;

    IsEmpty(me) returns Boolean from Standard
    ---Purpose: returns true if the directory is empty.
    is static;
    
---Category: Private methods
   
   List(me) returns ListOfDocument from CDM
   is static private;
   ---C++: return const &
   --      
   
fields

    myDocuments: ListOfDocument from CDM;

friends    
    class DirectoryIterator from CDF

end Directory from CDF;
