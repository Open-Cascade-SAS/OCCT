-- File:	IGESGeom_ToolRuledSurface.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolRuledSurface  from IGESGeom

    ---Purpose : Tool to work on a RuledSurface. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses RuledSurface from IGESGeom,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolRuledSurface;
    ---Purpose : Returns a ToolRuledSurface, ready to work


    ReadOwnParams (me; ent : mutable RuledSurface;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : RuledSurface;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : RuledSurface;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a RuledSurface <ent>, from
    --           its specific (own) parameters

    DirChecker (me; ent : RuledSurface) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : RuledSurface;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : RuledSurface; entto : mutable RuledSurface;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : RuledSurface;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolRuledSurface;
