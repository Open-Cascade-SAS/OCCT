-- File:	CircPnt2dBisec.cdl
-- Created:	Wed Apr  3 11:29:37 1991
-- Author:	Remi GILET
--		<reg@topsn2>
---Copyright:	 Matra Datavision 1991


class CircPnt2dBisec

from GccAna

	---Purpose: Describes functions for building a bisecting curve
    	-- between a 2D circle and a point.
    	-- A bisecting curve between a circle and a point is such a
    	-- curve that each of its points is at the same distance from
    	-- the circle and the point. It can be an ellipse, hyperbola,
    	-- circle or line, depending on the relative position of the
    	-- point and the circle. The algorithm computes all the
    	-- elementary curves which are solutions.
    	-- A CircPnt2dBisec object provides a framework for:
    	-- -   defining the construction of the bisecting curves,
    	-- -   implementing the construction algorithm, and
    	-- -   consulting the result.
  

uses Circ2d from gp,
     Pnt2d  from gp,
     Bisec  from GccInt
     
raises OutOfRange        from Standard,
       NotDone           from StdFail

is

Create(Circle1  : Circ2d from gp;
       Point2   : Pnt2d  from gp) returns CircPnt2dBisec;

    	---Purpose: Constructs bisecting curves between the circle Circle1 and the point Point2.
    
IsDone(me) returns Boolean from Standard
is static;
    	---Purpose: Returns true (this construction algorithm never fails).
    
NbSolutions(me) returns Integer from Standard
raises NotDone
is static;
    	---Purpose: Returns the number of curves, representing solutions computed by this algorithm.
    
ThisSolution(me                           ; 
    	     Index : Integer from Standard) returns Bisec from GccInt
raises OutOfRange, NotDone
is static;
    	---Purpose: Returns the solution number Index and raises OutOfRange 
    	--          exception if Index is greater than the number of solutions.
    	-- Exceptions
    	-- Standard_OutOfRange if Index is less than zero or
    	-- greater than the number of solutions computed by this algorithm.
fields

    WellDone : Boolean from Standard;
    	---Purpose: True if the algorithm succeeded.

    NbrSol   : Integer from Standard;
    	---Purpose: The number of possible solutions. We have to decide about the
    	--          status of the multiple solutions...

    circle   : Circ2d from gp;
    	---Purpose: The first argument used for ThisSolution.

    point   : Pnt2d from gp;
    	---Purpose: The second argument used for ThisSolution.

    theposition : Integer from Standard;
    	---Purpose: theposition = 1 when the point is outside the circle.
    	--          theposition = 0 when the point is on the circle.
    	--          theposition = -1 when the point is inside the circle.

end CircPnt2dBisec;
