-- Created on: 1992-09-24
-- Created by: Denis PASCAL
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

generic class DFSIterator from GraphTools 
	                 (Graph     as any;
                          Vertex    as any;
			  VHasher   as any;
                          VIterator as any)

    ---Purpose: This generic  class implement  the Depth  First Search
    --          algorithm from  a  Vertex with an iterator  to reached
    --          adjacent vertices of a  given  one.  The  interface of
    --          this algorithm is made as an iterator.

--generic class DFSIterator from GraphTools
--            (Graph     as any;
--    	       Vertex    as any;
--    	       VHasher   as MapHasher from TCollection (Vertex);
--	       VIterator as VertexIterator (Graph,Vertex))

raises NoMoreObject from Standard,
       NoSuchObject from Standard

    class DFSMap   instantiates IndexedMap from TCollection (Vertex,VHasher); 
    
is

    Create
    returns DFSIterator;
	---Purpose: Create an empty iterator.

    Perform (me : in out; G : Graph; V : Vertex);
	---Purpose: Initializes the research from <V> member vertex of
	--          <G>.
        ---Level: Public

    More (me) returns Boolean from Standard;
	---Purpose: Returns True if there are other vertices.
        ---Level: Public

    Next(me : in out) 
    	---Purpose: Set the iterator to the next vertex.
        ---Level: Public
    raises NoMoreObject from Standard;

    Value (me) returns any Vertex 
	---Purpose: returns the vertex  value for the current position
	--          of the iterator.
	---C++: return const &
        ---Level: Public
    raises NoSuchObject from Standard;


fields

    myVisited      : DFSMap from GraphTools;
    myCurrentIndex : Integer from Standard;

end DFSIterator;
    
    








