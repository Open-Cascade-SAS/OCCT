-- Created on: 1995-09-21
-- Created by: Philippe GIRODENGO
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class MeshTriangle from StlMesh inherits TShared from MMgt

	---Purpose: A  mesh triangle is defined with
	--          three geometric vertices and an orientation
	--          

raises 

    NegativeValue from Standard

is

    Create  returns mutable MeshTriangle;
    	---Purpose: empty constructor


    Create (V1, V2, V3 : Integer; Xn, Yn, Zn : Real)  returns mutable MeshTriangle
        ---Purpose: create a triangle defined with the indexes of its three vertices 
        --          and its orientation
    raises NegativeValue;
    	---Purpose: Raised if V1, V2 or V3 is lower than zero


    GetVertexAndOrientation (me; V1, V2, V3 : out Integer; Xn, Yn, Zn : out Real);
        ---Purpose: get indexes of the three vertices (V1,V2,V3) and the orientation

    SetVertexAndOrientation (me : mutable; V1, V2, V3 : in Integer; Xn, Yn, Zn : in Real)
        ---Purpose: set indexes of the three vertices (V1,V2,V3) and the orientation
    raises NegativeValue;
    	---Purpose: Raised if V1, V2 or V3 is lower than zero


    GetVertex  (me; V1, V2, V3 : out Integer);
        ---Purpose: get indexes of the three vertices (V1,V2,V3)

    SetVertex  (me : mutable; V1, V2, V3 : in Integer)
        ---Purpose: set indexes of the three vertices (V1,V2,V3)
    raises NegativeValue;
    	---Purpose: Raised if V1, V2 or V3 is lower than zero


fields 

    MyV1     : Integer;
    MyV2     : Integer;
    MyV3     : Integer;
    MyXn     : Real;
    MyYn     : Real;
    MyZn     : Real;

end MeshTriangle;


