-- Created on: 1992-10-02
-- Created by: Christian CAILLET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class AllConnected  from IFGraph  inherits GraphContent

    	---Purpose : this class gives content of the CONNECTED COMPONANT(S)
    	--           which include specific Entity(ies)

uses Transient, EntityIterator, Graph

is

    Create (agraph : Graph) returns AllConnected;
    ---Purpose : creates an AllConnected from a graph, empty ready to be filled

    Create (agraph : Graph; ent : any Transient)
    	returns AllConnected;
    ---Purpose : creates an AllConnected which memorizes Entities Connected to
    --           a given one, at any level : that is, itself, all Entities
    --           Shared by it and Sharing it, and so on.
    --           In other terms, this is the content of the CONNECTED COMPONANT
    --           which include a specific Entity

    GetFromEntity (me : in out; ent : any Transient);
    ---Purpose : adds an entity and its Connected ones to the list (allows to
    --           cumulate all Entities Connected by some ones)
    --           Note that if "ent" is in the already computed list,, no entity
    --           will be added, but if "ent" is not already in the list, a new
    --           Connected Componant will be cumulated 

    ResetData (me : in out);
    ---Purpose : Allows to restart on a new data set

    	-- --   Results   -- --
    	--   More-Next-Value give all entities noted in Connected Componant,
    	--   including the entities given for construction or to GetFromEntity

    Evaluate (me : in out) is redefined;
    ---Purpose : does the specific evaluation (Connected entities atall levels)

fields

    thegraph : Graph;

end AllConnected;
