-- Created on: 1993-06-22
-- Created by: Jean Louis FRENKEL, Gerard GRAS
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


-- Modified: TCL G002, 07-08-00, new inquire methods Center, Radius, FirstAngle, SecondAngle
--                               new methods SetRadius, SetCenter, SetAngles


class Circle from Graphic2d inherits Line from Graphic2d

	---Purpose: Constructs a primitive Circle

	
uses
	Drawer		from Graphic2d,
	GraphicObject	from Graphic2d,
	Length		from Quantity,
	PlaneAngle	from Quantity,
	FStream		from Aspect,
	IFStream	from Aspect

raises
	CircleDefinitionError	from Graphic2d

is
	-------------------------
	-- Category: Constructors
	-------------------------

	Create (aGraphicObject: GraphicObject from Graphic2d;
		X, Y: Length from Quantity;
		Radius: Length from Quantity)
	returns mutable Circle from Graphic2d
	---Level: Public
	---Purpose: Creates a complete circle.
	--	    The center is <X>, <Y>.
	--	    The radius is <Radius>.
	--  Warning: Raises CircleDefinitionError if the
	--          radius is null.
	raises CircleDefinitionError from Graphic2d;

	Create (aGraphicObject: GraphicObject from Graphic2d;
		X, Y: Length from Quantity;
		Radius: Length from Quantity;
		Alpha, Beta: PlaneAngle from Quantity)
	returns mutable Circle from Graphic2d
	---Level: Public
	---Purpose: Creates an arc.
	--	    The center is <X>, <Y>.
	--	    The radius is <Radius>.
	--	    Angles are measured counterclockwise with 0 radian
	--	    at 3 o'clock.
	--  Warning: Raises CircleDefinitionError if the
	--          radius is null.
	raises CircleDefinitionError from Graphic2d;

	----------------------------
	-- Category: Inquire methods
	----------------------------

	Center( me; X, Y: out Length from Quantity );  
	---Level: Public
	---Purpose: returns the coordinates of center of the circle
	
	Radius( me ) returns Length from Quantity;
	---Level: Public
	---Purpose: returns the radius of this circle
	
	FirstAngle( me ) returns PlaneAngle from Quantity;
	---Level: Public
	---Purpose: returns the first angle of the arc
	
	SecondAngle( me ) returns PlaneAngle from Quantity;
	---Level: Public
	---Purpose: returns the second angle of the arc
	

	--------------------------------------------------------
	-- Category: Methods for the definition of the circle's properties
	--------------------------------------------------------

	SetCenter( me: mutable; X, Y: Length from Quantity );  
	---Level: Public
	---Purpose: defines the coordinates of center of the circle
	
	SetRadius( me: mutable; theR: Length from Quantity );
	---Level: Public
	---Purpose: defines the radius of this circle
	
	SetAngles( me: mutable; Alpha, Beta: PlaneAngle from Quantity );
	---Level: Public
	---Purpose: defines the angles of the arc

	--------------------------
	-- Category: Draw and Pick
	--------------------------

	Draw (me : mutable; aDrawer: Drawer from Graphic2d)
	is static protected;
	---Level: Internal
	---Purpose: Draws the circle <me>.

	DrawElement( me : mutable; aDrawer: Drawer from Graphic2d;
		 anIndex: Integer from Standard)
	is redefined protected;
	---Level: Internal
	---Purpose: Draws element <anIndex> of the circle <me>.

	DrawVertex( me : mutable; aDrawer: Drawer from Graphic2d;
		anIndex: Integer from Standard)
	is redefined protected;
	---Level: Internal
	---Purpose: Draws vertex <anIndex> of the circle <me>.

	Pick (me : mutable; X, Y: ShortReal from Standard;
		aPrecision: ShortReal from Standard;
		aDrawer: Drawer from Graphic2d)
	returns Boolean from Standard is static protected;
	---Level: Internal
	---Purpose: Returns Standard_True if the circle <me> is picked,
	--	    Standard_False if not.

	DoMinMax( me: mutable ) is private;

	----------------------------------------------------------------------

	Save( me; aFStream: in out FStream from Aspect ) is virtual;
	Retrieve( myclass; anIFStream: in out IFStream from Aspect;
		aGraphicObject: GraphicObject from Graphic2d );

fields

	myX:		ShortReal from Standard;
	myY:		ShortReal from Standard;
	myRadius:	ShortReal from Standard;
	myFirstAngle:	ShortReal from Standard;
	mySecondAngle:	ShortReal from Standard;
	myisArc:	Boolean from Standard;

end Circle from Graphic2d;
