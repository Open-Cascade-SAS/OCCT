-- Created on: 1996-03-06
-- Created by: Laurent BOURESCHE
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class CircSection from ChFiDS 

	---Purpose: A Section of fillet.

uses
    Circ from gp,
    Lin  from gp
is
    Create;

    Set(me  : in out;
    	C   : Circ from gp;
	F,L : Real from Standard)
    is static;
    
    Set(me  : in out;
    	C   : Lin  from gp;
	F,L : Real from Standard)
    is static;

    Get(me;
    	C   : out Circ from gp;
	F,L : out Real from Standard)
    is static;
    
    Get(me;
    	C   : out Lin  from gp;
	F,L : out Real from Standard)
    is static;

fields
    myCirc : Circ from gp;
    myLin  : Lin  from gp;
    myF    : Real from Standard;
    myL    : Real from Standard;
end CircSection;
