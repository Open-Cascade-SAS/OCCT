-- File:	MXCAFDoc_AreaRetrievalDriver.cdl
-- Created:	Fri Sep  8 18:26:44 2000
-- Author:	data exchange team
--		<det@nordox.nnov.matra-dtv.fr>
---Copyright:	 Matra Datavision 2000


class AreaRetrievalDriver from MXCAFDoc inherits ARDriver from MDF

	---Purpose: 
uses
    RRelocationTable from MDF,
    Attribute        from PDF,
    Attribute        from TDF,
    MessageDriver    from CDM

is
--    Create  
--    returns mutable AreaRetrievalDriver from MXCAFDoc;
    Create (theMsgDriver : MessageDriver from CDM)
    returns mutable AreaRetrievalDriver from MXCAFDoc;

    VersionNumber(me) returns Integer from Standard;
	---Purpose: Returns the version number from which the driver
	--          is available: 0.

    SourceType(me) returns Type from Standard;
    ---Purpose: Returns the type: XCAFDoc_Area

    NewEmpty (me)  returns mutable Attribute from TDF;

    Paste(me;
    	  Source     :         Attribute from PDF;
    	  Target     : mutable Attribute from TDF;
    	  RelocTable : RRelocationTable from MDF);

end AreaRetrievalDriver from MXCAFDoc;
