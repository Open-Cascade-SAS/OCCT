-- Created on: 2008-01-20
-- Created by: Alexander A. BORODIN
-- Copyright (c) 2008-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SystemFont from Font inherits TShared from MMgt
---Purpose: Structure for store of Font System Information

uses FontAspect,
     HAsciiString from TCollection

is
  Create returns SystemFont;
  ---Purpose: Creates empty font object
  ---Level: Public

  Create (theFontName   : HAsciiString;
          theFontAspect : FontAspect;
          theFilePath   : HAsciiString ) returns SystemFont;
  ---Purpose: Creates Font object initialized with <FontName> as name
  ---         <FontAspect>.... TODO
  ---Level: Public

  Create (theXLFD     : HAsciiString;
          theFilePath : HAsciiString ) returns SystemFont;
  ---Purpose: Creates Font object and initialize class fields with
  ---         values taken from XLFD (X Logical Font Description)
  ---Level: Public
 
  FontName (me) returns HAsciiString;
  --- Purpose: Returns font family name
  ---Level: Public    
        
  FontPath (me) returns HAsciiString;
  --- Purpose: Returns font file path
  --- Level: Public

  FontAspect (me) returns FontAspect;
  --- Purpose: Returns font aspect
  --- Level: Public
    
  FontHeight (me) returns Integer from Standard;
  --- Purpose: Returns font height
  --- If returned value is equal -1 it means that font is resizable
  --- Level: Public

  IsValid (me) returns Boolean;
  
  IsEqual (me;
           theOtherFont: SystemFont) returns Boolean;
  --- Purpose: Return true if the FontName, FontAspect and FontSize are the same.
  --- Level: Public
  
fields
  MyFontName:           HAsciiString;  --Font family name
  MyFontAspect:         FontAspect;    
  MyFaceSize:           Integer;       --height of font
  MyFilePath:           HAsciiString;  --absolute path to font file
  MyVerification:       Boolean;       --indicator of font initialization errors. False if initialization is failed.

end SystemFont;
