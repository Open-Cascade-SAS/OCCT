-- Created on: 2002-03-04
-- Created by: Michael KLOKOV
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SectionAttribute from BOPAlgo
    ---Purpose: Class is a container of three flags used
    ---         by intersection algorithm
    ---

is

    Create(Aproximation : Boolean from Standard = Standard_True;
           PCurveOnS1   : Boolean from Standard = Standard_True;
           PCurveOnS2   : Boolean from Standard = Standard_True)
    returns SectionAttribute from BOPAlgo;
    ---Purpose:
    --- Initializes me by flags
    
    Approximation(me: in out; theFlag: Boolean from Standard);
    ---Purpose:
    --- Modifier
    ---
    
    PCurveOnS1(me: in out; theFlag: Boolean from Standard);
    ---Purpose:
    --- Modifier
    ---
    
    PCurveOnS2(me: in out; theFlag: Boolean from Standard);
    ---Purpose:
    --- Modifier
    ---

    Approximation(me)
    returns Boolean from Standard;
    ---C++: inline
    ---Purpose:
    --- Selector
    ---
    
    PCurveOnS1(me)
    returns Boolean from Standard;
    ---C++: inline
    ---Purpose:
    --- Selector
    ---
    
    PCurveOnS2(me)
    returns Boolean from Standard;
    ---C++: inline
    ---Purpose:
    --- Selector
    ---

fields
    myApproximation : Boolean from Standard;
    myPCurve1       : Boolean from Standard;
    myPCurve2       : Boolean from Standard;

end SectionAttribute from BOPAlgo;
