-- Created on: 1994-12-16
-- Created by: Frederic MAUPAS
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class TranslateVertexLoop from StepToTopoDS
    inherits Root from StepToTopoDS
    
    ---Purpose:
    --         

uses

    VertexLoop               from StepShape,
    TranslateVertexLoopError from StepToTopoDS,
    Tool                     from StepToTopoDS,
    Shape                    from TopoDS,
    NMTool                   from StepToTopoDS

raises NotDone from StdFail

is

    Create returns TranslateVertexLoop;
    
    Create (VL     : VertexLoop    from StepShape;
            T      : in out Tool   from StepToTopoDS;
            NMTool : in out NMTool from StepToTopoDS)
    	returns TranslateVertexLoop;
	    
    Init (me     : in out;
          VL     : VertexLoop    from StepShape;
          T      : in out Tool   from StepToTopoDS;
          NMTool : in out NMTool from StepToTopoDS);

    Value (me) returns Shape from TopoDS
    	raises NotDone
	is static;
	---C++: return const &

    Error (me) returns TranslateVertexLoopError from StepToTopoDS;
    
fields

    myError  : TranslateVertexLoopError from StepToTopoDS;
    
    myResult : Shape                    from TopoDS;
    
end TranslateVertexLoop;
