-- Created on: 1992-08-11
-- Created by: Remi LEQUETTE
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package TopCnx 

	---Purpose: This  algorithm  provides  algorithms  to computes
	--          transitions when many interferences occurs  at the
	--          same place on a shape.
	--          
	--          An interference is an intersection on a shape (i.e
	--          a vertex on an  edge  or an edge  on a  face) with
	--          data  about    the  transition (how  the  shape is
	--          crossing  the   boundary  where the   intersection
	--          occurs).
	--          
	--          There     are      three  algorithms   to  process
	--          interferences : 
	--          
	--          * EdgeFaceTransition : To process interferences on
	--          an adge crossing other edges  on the boundary of a
	--          face.
	--          
	--          * EdgeSolidTransition : To   process interferences
	--          on  an   edge  crossing  faces   and edges  on the
	--          boundary of a solid.
	--          
	--          *  FaceSolidTransition : To  process interferences
	--          on a face crossing other faces on  the boundary of
	--          a solid.
	--          
	--          This package  relies on the  TopTrans  package for
	--          the geometric computations.

uses
    Standard,
    gp,
    TopAbs,
    TopTrans

is
    class EdgeFaceTransition;
	---Purpose: Algorithm  to compute cumulated transitions  on an
	--          edge crossing the boundary of a face.

end TopCnx;
