-- Created on: 1999-11-26
-- Created by: Andrey BETENEV
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0

class ActionRequestSolution from StepBasic
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity ActionRequestSolution

uses
    ActionMethod from StepBasic,
    VersionedActionRequest from StepBasic

is
    Create returns ActionRequestSolution from StepBasic;
	---Purpose: Empty constructor

    Init (me: mutable; aMethod: ActionMethod from StepBasic;
                       aRequest: VersionedActionRequest from StepBasic);
	---Purpose: Initialize all fields (own and inherited)

    Method (me) returns ActionMethod from StepBasic;
	---Purpose: Returns field Method
    SetMethod (me: mutable; Method: ActionMethod from StepBasic);
	---Purpose: Set field Method

    Request (me) returns VersionedActionRequest from StepBasic;
	---Purpose: Returns field Request
    SetRequest (me: mutable; Request: VersionedActionRequest from StepBasic);
	---Purpose: Set field Request

fields
    theMethod: ActionMethod from StepBasic;
    theRequest: VersionedActionRequest from StepBasic;

end ActionRequestSolution;
