-- Created on: 1999-03-09
-- Created by: data exchange team
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class ShapeUpgrade from SWDRAW 

	---Purpose: Contains commands to activate package ShapeUpgrade
	--          List of DRAW commands and corresponding functionalities:
	--          DT_ShapeDivide         - ShapeUpgrade_ShapeDivide
	--          DT_PlaneDividedFace    - ShapeUpgrade_PlaneDividedFace
	--          DT_PlaneGridShell      - ShapeUpgrade_PlaneGridShell
	--          DT_PlaneFaceCommon     - ShapeUpgrade_PlaneFaceCommon
	--          DT_Split2dCurve        - ShapeUpgrade_Split2dCurve
	--          DT_SplitCurve          - ShapeUpgrade_SplitCurve
	--          DT_SplitSurface        - ShapeUpgrade_SplitSurface
	--          DT_SupportModification - ShapeUpgrade_DataMapOfShapeSurface
	--          DT_Debug               - ShapeUpgrade::SetDebug
	--          shellsolid             - ShapeAnalysis_Shell/ShapeUpgrade_ShellSewing
	
uses
    Interpretor from Draw

is

    InitCommands (myclass; theCommands: in out Interpretor from Draw);
    	---Purpose: Loads commands defined in ShapeUpgrade

end ShapeUpgrade;
