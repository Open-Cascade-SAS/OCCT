-- Created on: 1998-05-06
-- Created by: Andre LIEUTIER
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PlaneConstraint from Plate
---Purpose: constraint a point to belong to a Plane
--          

uses 
 XY from gp, 
 Pln  from  gp,
 LinearScalarConstraint from Plate

is
    Create(point2d : XY ; pln  :  Pln  from  gp; 
           iu : Integer = 0; iv : Integer = 0) returns PlaneConstraint;
-- constraint the iu th derivative in u  and iv th  derivative in v at
-- the point2d parametre to belong to the pln plane.

    -- Accessors :
    LSC(me) returns  LinearScalarConstraint ;
    ---C++: inline 
    ---C++: return const &

fields
    myLSC : LinearScalarConstraint;    
end;

