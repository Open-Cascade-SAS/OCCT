-- Created on: 1995-12-07
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PointClassifier from TopOpeBRep

uses 

    State from TopAbs,
    Face from TopoDS,
    Pnt2d from gp,
    TopolTool from BRepTopAdaptor,
    HSurface from BRepAdaptor,
    DataMapOfTopolTool from TopOpeBRep    
    
is

    Create returns PointClassifier from TopOpeBRep;
    
    Init(me:in out) is static;
    
    Load(me:in out;F:Face from TopoDS) is static;

    Classify(me:in out;F:Face from TopoDS;P:Pnt2d from gp;Tol:Real)
    ---Purpose: compute position of point <P> regarding with the face <F>. 
    returns State from TopAbs is static;

    State(me) returns State from TopAbs is static;    

fields

    myTopolTool : TopolTool from BRepTopAdaptor;
    myHSurface : HSurface from BRepAdaptor;
    myTopolToolMap : DataMapOfTopolTool from TopOpeBRep;
    myState : State from TopAbs;
    
end PointClassifier from TopOpeBRep;
