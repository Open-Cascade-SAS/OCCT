-- Created on: 1993-04-06
-- Created by: Philippe DAUTRY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class OffsetCurve from PGeom2d inherits Curve from PGeom2d

        ---Purpose :
        --  This class implements the basis services for an offset curve
        --  in 3D space.
        --  
	---See Also : OffsetCurve from Geom2d.

uses Curve from PGeom2d


is
    

  Create returns mutable OffsetCurve from PGeom2d;
    ---Purpose: Creates an OffsetCurve with default values.
	---Level: Internal 


  Create (
    	    aBasisCurve : Curve from PGeom2d;
    	    aOffsetValue : Real from Standard)
     returns mutable OffsetCurve from PGeom2d;
        ---Purpose : <aBasisCurve> is  the basis curve, <aOffsetValue>
        --         is the distance between <me> and the basis curve at
        --         any point.    <aOffsetDirection>  defines the fixed
        --         reference direction (offset direction).
	---Level: Internal 


  BasisCurve (me : mutable; aBasisCurve : Curve from PGeom2d);
	---Purpose: Set the field basisCurve with <aBasisCurve>.
	---Level: Internal 
      

  BasisCurve (me) returns Curve from PGeom2d;
        ---Purpose : The basis curve can be an offset curve.
	---Level: Internal 


  OffsetValue (me : mutable; aOffsetValue : Real from Standard);
        ---Purpose : Set the field offsetValue with <aOffsetValue>.
	---Level: Internal 


  OffsetValue (me) returns Real from Standard;
        ---Purpose : Returns the value of the field offsetValue.
	---Level: Internal 


fields

  basisCurve      : Curve from PGeom2d;
  offsetValue     : Real from Standard;

end;
