-- Created on: 1994-02-23
-- Created by: model
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

generic class GenHCurve from Adaptor3d 
    (TheCurve as Curve from Adaptor3d)

inherits HCurve from Adaptor3d 

	---Purpose: Generic class used to create a curve manipulated
      	--          with Handle from a curve described by the class Curve.

uses 
     Curve        from Adaptor3d

     
raises
    
    OutOfRange          from Standard,
    NoSuchObject        from Standard,
    DomainError         from Standard
 
is

    Create
	---Purpose: Creates an empty GenHCurve.
    	returns mutable GenHCurve from Adaptor3d; 
    

    Create(C: TheCurve)
    
	---Purpose: Creates a GenHCurve from a Curve
    	returns mutable GenHCurve from Adaptor3d; 


    Set(me: mutable; C: TheCurve)
    
	---Purpose: Sets the field of the GenHCurve.
    	is static;

    Curve(me)
    
	---Purpose: Returns the curve used to create the GenHCurve.
	--          This is redefined from HCurve, cannot be inline.
	--          
	---C++: return const &

    	returns Curve from Adaptor3d;

    GetCurve(me:mutable)
    
	---Purpose: Returns the curve used to create the GenHCurve.
	--          This is redefined from HCurve, cannot be inline.
	--          
	---C++: return  &

    	returns Curve from Adaptor3d;


    ChangeCurve(me : mutable)
    
	---Purpose: Returns the curve used to create the GenHCurve.
	--          
	---C++: return &
	---C++: inline

    	returns TheCurve;

fields

    myCurve : TheCurve is protected;

end GenHCurve;
