-- Created on: 2010-12-03
-- Created by: Artem SHAL
-- Copyright (c) 2010-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Sphere from Bnd

    ---Purpose: This class represents a bounding sphere of a geometric entity
    --          (triangle, segment of line or whatever else).

uses XYZ from gp

is

    Create returns Sphere;
	    ---Purpose: Empty constructor

    Create (theCntr : XYZ from gp; theRad : Real; theU : Integer; theV : Integer)
	    returns Sphere;
	    ---Purpose: Constructor of a definite sphere

    U (me) returns Integer;
        ---C++: inline
        ---Purpose: Returns the U parameter on shape

    V (me) returns Integer;
        ---C++: inline
        ---Purpose: Returns the V parameter on shape

    IsValid (me) returns Boolean;
        ---C++: inline
	    ---Purpose: Returns validity status, indicating that this
	    --		sphere corresponds to a real entity

    SetValid (me : in out; isValid : Boolean);
        ---C++: inline

    Center (me) returns XYZ from gp;
        ---C++: inline
	    ---C++: return const &
	    ---Purpose: Returns center of sphere object

    Radius (me) returns Real;
        ---C++: inline
	    ---Purpose: Returns the radius value

    Distances (me; theXYZ : XYZ from gp; theMin : in out Real; theMax : in out Real) is static;
	    ---Purpose: Calculate and return minimal and maximal distance to sphere.
	    --		NOTE: This function is tightly optimized; any modifications
	    --		may affect performance!
	    
    SquareDistances (me; theXYZ : XYZ from gp; theMin : in out Real; theMax : in out Real) is static;
	    ---Purpose: Calculate and return minimal and maximal distance to sphere.
	    --		NOTE: This function is tightly optimized; any modifications
	    --		may affect performance!

    Project (me; theNode : XYZ from gp; theProjNode : in out XYZ from gp; theDist : in out Real; theInside : in out Boolean)
	    ---Purpose: Projects a point on entity.
	    --		   Returns true if success
	    returns Boolean;

    Distance (me; theNode : XYZ from gp)
	    returns Real;
	    
    SquareDistance (me; theNode : XYZ from gp)
	    returns Real;

    Add (me : in out; theOther : Sphere from Bnd);

    IsOut (me; theOther : Sphere from Bnd)
	    returns Boolean;

    IsOut (me; thePnt : XYZ from gp; theMaxDist : in out Real)
	    returns Boolean;

    SquareExtent (me) returns Real;

fields

    myCenter	: XYZ from gp;
    myRadius	: Real;
    myIsValid	: Boolean;
    myU		: Integer;
    myV		: Integer;

end Sphere;
