-- Created on: 2002-12-10
-- Created by: data exchange team
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V2.0

class CurveElementFreedomMember from StepElement
inherits SelectNamed from StepData

    ---Purpose: Representation of member for  STEP SELECT type CurveElementFreedom

is
    Create returns CurveElementFreedomMember from StepElement;
	---Purpose: Empty constructor

    HasName (me) returns Boolean  is redefined;
	---Purpose: Returns True if has name

    Name (me) returns CString  is redefined;
	---Purpose: Returns set name 

    SetName (me : mutable; name : CString)  returns Boolean  is redefined;
	---Purpose: Set name 

    Matches (me; name : CString) returns Boolean  is redefined;
	---Purpose : Tells if the name of a SelectMember matches a given one;

fields

    mycase : Integer;

end CurveElementFreedomMember;
