-- Created on: 1993-06-03
-- Created by: Jean-Louis FRENKEL
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class AngleAspect from Prs3d inherits CompositeAspect from Prs3d 

    	---Purpose: A framework for defining how an angle will be
    	-- displayed in a presentation. Aspects of angle display include:
    	-- -   display of the arrow pointing to the angle
    	-- -   display of the line making up the shaft of the arrow
    	-- -   display of the text referring to the angle.
    	--   The definition set by this class is then passed to the
    	-- attribute manager Prs3d_Drawer.
    	-- Any object which requires a value for angle aspect as
    	-- an argument may then be given the attribute manager
    	-- as a substitute argument in the form of a field such as
    	-- myDrawer for example.
        
uses 

    LineAspect from Prs3d,
    TextAspect from Prs3d,
    ArrowAspect from Prs3d

is

-- 
--  Attributes for the lines.
-- 
    Create returns mutable AngleAspect from Prs3d;

    LineAspect(me) returns mutable LineAspect from Prs3d;
    	--- Purpose: Returns the setting determining how the line making
    	-- up the shaft of the arrow will be displayed.   
    
    SetLineAspect(me: mutable; anAspect: LineAspect from Prs3d);
    	---Purpose: Sets how the line making up the shaft of an arrow will be displayed.
    TextAspect(me) returns mutable TextAspect from Prs3d is static;
    	--- Purpose: Returns the setting determining how text in the
    	-- presentation of an angle will be displayed.   
    
    SetTextAspect(me:mutable; anAspect: TextAspect from Prs3d) is static;
    	---Purpose: Sets how text in the presentation of an angle will be displayed.
    ArrowAspect(me) returns mutable ArrowAspect from Prs3d is static;
    	---Purpose: Returns the setting determining how an arrow head
    	-- which points to an angle will be displayed.    
    
    SetArrowAspect(me: mutable; anAspect: ArrowAspect from Prs3d) is static;
    	---Purpose: Sets how an arrow head which points to an angle will be displayed.

fields

    myLineAspect: LineAspect from Prs3d;
    myArrowAspect: ArrowAspect from Prs3d;
    myTextAspect: TextAspect from Prs3d;
    
end AngleAspect from Prs3d;
