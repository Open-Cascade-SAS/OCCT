-- Created on: 2000-08-22
-- Created by: Andrey BETENEV
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class UOperator from ShapeProcess inherits Operator from ShapeProcess

    ---Purpose: Defines operator as container for static function
    --          OperFunc. This allows user to create new operators 
    --          without creation of new classes

uses

    OperFunc from ShapeProcess,
    Context from ShapeProcess

is

    Create (func: OperFunc from ShapeProcess);
    	---Purpose: Creates operator with implementation defined as
	--          OperFunc (static function)

    Perform (me: mutable; context: Context from ShapeProcess) 
    returns Boolean is redefined;
    	---Purpose: Performs operation and records changes in the context

fields

    myFunc: OperFunc from ShapeProcess;

end UOperator;
