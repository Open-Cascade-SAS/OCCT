-- File:        EdgeLoop.cdl
-- Created:     Mon Dec  4 12:02:26 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWEdgeLoop from RWStepShape

	---Purpose : Read & Write Module for EdgeLoop
	--           Check added by CKY , 7-OCT-1996

uses Check from Interface, ShareTool from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     EdgeLoop from StepShape,
     EntityIterator from Interface

is

	Create returns RWEdgeLoop;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable EdgeLoop from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : EdgeLoop from StepShape);

    	Share(me; ent : EdgeLoop from StepShape; iter : in out EntityIterator);

    	Check(me; ent : EdgeLoop from StepShape; shares : ShareTool; ach : in out Check);

end RWEdgeLoop;
