-- File:	StepData_SelectArrReal.cdl
-- Created:	Wed Dec 18 09:07:30 2002
-- Author:	data exchange team
--		<det@petrox.nnov.matra-dtv.fr>
---Copyright:	 Matra Datavision 2002

class SelectArrReal from StepData inherits SelectNamed from StepData

    ---Purpose :


uses

    AsciiString from TCollection,
    HArray1OfReal from TColStd

is

    Create returns mutable SelectArrReal;

--    HasName (me) returns Boolean  is redefined;

--    Name (me) returns CString  is redefined;

--    SetName (me : mutable; name : CString)  returns Boolean  is redefined;
    -- redefined to accept any name

    Kind(me) returns Integer  is redefined;
    --  fixed kind : ArrReal

    ArrReal(me) returns HArray1OfReal from TColStd;

    SetArrReal(me:mutable; arr : HArray1OfReal from TColStd);

fields

    theArr  : HArray1OfReal from TColStd;

end SelectArrReal;
