-- File:	QADBMReflex_OCC749Prs.cdl
-- Created:	Mon Oct  7 15:01:08 2002
-- Author:	QA Admin
--		<qa@russox>
---Copyright:	 Matra Datavision 2002

class OCC749Prs from QADBMReflex inherits InteractiveObject from AIS

uses
    PresentationManager3d from PrsMgr,
    Presentation          from Prs3d,
    Selection             from SelectMgr,
    Color                 from Quantity,
    MaterialAspect        from Graphic3d

is
    Create( Reflection     : Boolean from Standard;
    	    InteriorColor  : Color from Quantity;
    	    EdgeColor      : Color from Quantity;
    	    EdgeColor2     : Color from Quantity;
    	    XCount         : Integer from Standard;
    	    YCount         : Integer from Standard;
    	    BoxSize        : Integer from Standard;
    	    MaterialAspect : MaterialAspect from Graphic3d;
    	    Material       : Boolean from Standard;
    	    Timer          : Boolean from Standard )
     returns mutable OCC749Prs from QADBMReflex;

    ComputeSelection(me          : mutable;
    	    	     aSelection  : mutable Selection from SelectMgr;
    	    	     aMode       : Integer from Standard)
    is redefined virtual protected;

    SetReflection( me : mutable; Reflection : Boolean from Standard );

    GetReflection( me )
    returns Boolean from Standard;

    SetColor( me : mutable; InteriorColor : Color from Quantity;
    	    	    	    EdgeColor     : Color from Quantity );

    GetInteriorColor( me )
    returns Color from Quantity;

    GetEdgeColor( me )
    returns Color from Quantity;

    SetEdgeColor2( me : mutable; EdgeColor2 : Color from Quantity );

    GetEdgeColor2( me )
    returns Color from Quantity;

    SetXYCount( me : mutable; XCount : Integer from Standard;
    	    	    	      YCount : Integer from Standard );

    GetXCount( me )
    returns Integer from Standard;

    GetYCount( me )
    returns Integer from Standard;

    SetBoxSize( me : mutable; BoxSize : Integer from Standard );

    GetBoxSize( me )
    returns Integer from Standard;

    SetMaterialAspect( me : mutable; MaterialAspect : MaterialAspect from Graphic3d );

    GetMaterialAspect( me )
    returns MaterialAspect from Graphic3d;

    SetMaterial( me : mutable; Material : Boolean from Standard );

    GetMaterial( me )
    returns Boolean from Standard;

    SetTimer( me : mutable; Timer : Boolean from Standard );

    GetTimer( me )
    returns Boolean from Standard;

fields
    myReflection     : Boolean from Standard;
    myInteriorColor  : Color from Quantity;
    myEdgeColor      : Color from Quantity;
    myEdgeColor2     : Color from Quantity;
    myXCount         : Integer from Standard;
    myYCount         : Integer from Standard;
    myBoxSize        : Integer from Standard;
    myMaterialAspect : MaterialAspect from Graphic3d;
    myMaterial       : Boolean from Standard;
    myTimer          : Boolean from Standard;
end OCC749Prs;
