-- File:        ProductContext.cdl
-- Created:     Mon Dec  4 12:02:29 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWProductContext from RWStepBasic

	---Purpose : Read & Write Module for ProductContext

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     ProductContext from StepBasic,
     EntityIterator from Interface

is

	Create returns RWProductContext;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable ProductContext from StepBasic);

	WriteStep (me; SW : in out StepWriter; ent : ProductContext from StepBasic);

	Share(me; ent : ProductContext from StepBasic; iter : in out EntityIterator);

end RWProductContext;
