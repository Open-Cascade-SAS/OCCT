-- File:	IGESBasic_ToolHierarchy.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolHierarchy  from IGESBasic

    ---Purpose : Tool to work on a Hierarchy. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses Hierarchy from IGESBasic,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolHierarchy;
    ---Purpose : Returns a ToolHierarchy, ready to work


    ReadOwnParams (me; ent : mutable Hierarchy;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : Hierarchy;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : Hierarchy;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a Hierarchy <ent>, from
    --           its specific (own) parameters

    OwnCorrect (me; ent : mutable Hierarchy) returns Boolean  is static;
    ---Purpose : Sets automatic unambiguous Correction on a Hierarchy
    --           (NbPropertyValues forced to 6)

    DirChecker (me; ent : Hierarchy) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : Hierarchy;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : Hierarchy; entto : mutable Hierarchy;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : Hierarchy;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolHierarchy;
