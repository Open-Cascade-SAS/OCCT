-- Created on: 1995-01-31
-- Created by: Mister rmi
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class SensitiveBox from Select2D 
inherits SensitiveEntity from Select2D

	---Purpose: defines a Sensitive Box (inside or boundary)

uses
    Pnt2d from gp,
    Box2d from Bnd,
    ListOfBox2d from SelectBasics,    
    EntityOwner from SelectBasics,
    TypeOfSelection

is
    Create (OwnerId      : EntityOwner from SelectBasics;
    	    Center       : Pnt2d from gp;
    	    Height,Width : Real from Standard;
    	    Type         : TypeOfSelection = Select2D_TOS_INTERIOR)
    returns mutable SensitiveBox;
    	---Purpose: Constructs a sensitive box object defined by the
    	-- owner OwnerId, the center point Center, the height
    	-- Height, the width Width, and the selection type Type.
    	-- Type can be:
    	-- -   interior
    	-- -   boundary.

    Create (OwnerId             : EntityOwner from SelectBasics;
    	    Xmin,YMin,XMax,YMax : Real;
    	    Type         : TypeOfSelection = Select2D_TOS_INTERIOR) 
    returns mutable SensitiveBox;
    
    	---Purpose: Constructs a sensitive box object defined by the
    	-- owner OwnerId, the coordinates Xmin, YMin, XMax,
    	-- YMax, and the selection type Type.
    	-- Xmin, YMin define the minimum point in the lower left
    	-- hand corner of the box, and   XMax, YMax define the
    	-- maximum point in the upper right hand corner of the box.
    	-- Type can be:
    	-- -   interior
    	-- -   boundary.    

    Areas   (me:mutable ; aresul : in out ListOfBox2d from SelectBasics) is static;
    
    
    Matches (me   : mutable; 
    	     X,Y  : Real from Standard;
    	     aTol : Real from Standard;
    	     DMin : out Real from Standard)
    returns Boolean is static;
    
    
    Matches (me  :mutable; 
             XMin,YMin,XMax,YMax : Real from Standard;
             aTol: Real from Standard) 
    returns Boolean
    is static;


fields

    mybox    : Box2d from Bnd;
    mytype   : TypeOfSelection;
    

end SensitiveBox;
