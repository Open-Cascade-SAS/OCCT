-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SurfacePatch from StepGeom 

inherits TShared from MMgt

uses

	BoundedSurface from StepGeom, 
	TransitionCode from StepGeom, 
	Boolean from Standard
is

	Create returns mutable SurfacePatch;
	---Purpose: Returns a SurfacePatch

	Init (me : mutable;
	      aParentSurface : mutable BoundedSurface from StepGeom;
	      aUTransition : TransitionCode from StepGeom;
	      aVTransition : TransitionCode from StepGeom;
	      aUSense : Boolean from Standard;
	      aVSense : Boolean from Standard) is virtual;

	-- Specific Methods for Field Data Access --

	SetParentSurface(me : mutable; aParentSurface : mutable BoundedSurface);
	ParentSurface (me) returns mutable BoundedSurface;
	SetUTransition(me : mutable; aUTransition : TransitionCode);
	UTransition (me) returns TransitionCode;
	SetVTransition(me : mutable; aVTransition : TransitionCode);
	VTransition (me) returns TransitionCode;
	SetUSense(me : mutable; aUSense : Boolean);
	USense (me) returns Boolean;
	SetVSense(me : mutable; aVSense : Boolean);
	VSense (me) returns Boolean;

fields

	parentSurface : BoundedSurface from StepGeom;
	uTransition : TransitionCode from StepGeom; -- an Enumeration
	vTransition : TransitionCode from StepGeom; -- an Enumeration
	uSense : Boolean from Standard;
	vSense : Boolean from Standard;

end SurfacePatch;
