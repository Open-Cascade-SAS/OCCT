-- Created on: 2005-05-17
-- Created by: Eugeny NAPALKOV <eugeny.napalkov@opencascade.com>
-- Copyright (c) 2005-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class LocationDriver from BinMXCAFDoc inherits ADriver from BinMDF

uses
    MessageDriver    from CDM,
    SRelocationTable from BinObjMgt,
    RRelocationTable from BinObjMgt,
    Persistent       from BinObjMgt,
    Location         from TopLoc,
    Attribute        from TDF,
    LocationSetPtr   from BinTools
is
    Create (theMsgDriver:MessageDriver from CDM)
    returns mutable LocationDriver from BinMXCAFDoc;

    NewEmpty (me)  returns mutable Attribute from TDF
    is redefined;

    Paste(me; theSource     : Persistent from BinObjMgt;
              theTarget     : mutable Attribute from TDF;
              theRelocTable : out RRelocationTable from BinObjMgt)
    returns Boolean from Standard is redefined;

    Paste(me; theSource     : Attribute from TDF;
              theTarget     : in out Persistent from BinObjMgt;
              theRelocTable : out SRelocationTable from BinObjMgt)
    is redefined;
    
    Translate(me; theSource     : Persistent from BinObjMgt;
	               theLoc        : in out Location from TopLoc;
         	       theMap        : out RRelocationTable from BinObjMgt)
    returns Boolean from Standard;
    
    Translate(me; theLoc        : Location from TopLoc;
    	    	       theTarget     : in out Persistent from BinObjMgt;
		       theMap        : out SRelocationTable from BinObjMgt);
    ---Purpose: Translate transient location to storable
    
    SetSharedLocations(me: mutable;
                       theLocations:  in LocationSetPtr  from BinTools);
    ---C++: inline
    
fields
    myLocations : LocationSetPtr   from BinTools;
end;
