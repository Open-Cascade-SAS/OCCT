-- Created on: 1992-08-21
-- Created by: Christophe MARION
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class BiPoint from HLRBRep

    	---Purpose: Contains the colors of a shape.

uses
    Boolean from Standard,
    Real    from Standard,
    Pnt     from gp,
    Shape   from TopoDS
    
is
    Create
    returns BiPoint from HLRBRep; 
    
    Create(x1,y1,z1,x2,y2,z2   : Real    from Standard;
           S                   : Shape   from TopoDS;
           reg1,regn,outl,intl : Boolean from Standard)
    returns BiPoint from HLRBRep; 
    
    P1(me) returns Pnt from gp
    	---C++: inline
    	---C++: return const &
    is static;

    P2(me) returns Pnt from gp
    	---C++: inline
    	---C++: return const &
    is static;

    Shape(me) returns Shape from TopoDS
    	---C++: inline
    	---C++: return const &
    is static;

    Shape(me : in out; S : Shape from TopoDS)
    	---C++: inline
    is static;

    Rg1Line(me) returns Boolean from Standard
    	---C++: inline
    is static;

    Rg1Line(me : in out; B : Boolean from Standard)
    	---C++: inline
    is static;

    RgNLine(me) returns Boolean from Standard
    	---C++: inline
    is static;

    RgNLine(me : in out; B : Boolean from Standard)
    	---C++: inline
    is static;

    OutLine(me) returns Boolean from Standard
    	---C++: inline
    is static;

    OutLine(me : in out; B : Boolean from Standard)
    	---C++: inline
    is static;

    IntLine(me) returns Boolean from Standard
    	---C++: inline
    is static;

    IntLine(me : in out; B : Boolean from Standard)
    	---C++: inline
    is static;

fields
    myP1    : Pnt     from gp;
    myP2    : Pnt     from gp;
    myShape : Shape   from TopoDS;
    myFlags : Boolean from Standard;

end BiPoint;
