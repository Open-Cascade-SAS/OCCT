-- Created on: 2002-12-12
-- Created by: data exchange team
-- Copyright (c) 2002-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class FeaModel from StepFEA
inherits Representation from StepRepr

    ---Purpose: Representation of STEP entity FeaModel

uses
    HAsciiString from TCollection,
    HArray1OfRepresentationItem from StepRepr,
    RepresentationContext from StepRepr,
    HArray1OfAsciiString from TColStd

is
    Create returns FeaModel from StepFEA;
	---Purpose: Empty constructor

    Init (me: mutable; aRepresentation_Name: HAsciiString from TCollection;
                       aRepresentation_Items: HArray1OfRepresentationItem from StepRepr;
                       aRepresentation_ContextOfItems: RepresentationContext from StepRepr;
                       aCreatingSoftware: HAsciiString from TCollection;
                       aIntendedAnalysisCode: HArray1OfAsciiString from TColStd;
                       aDescription: HAsciiString from TCollection;
                       aAnalysisType: HAsciiString from TCollection);
	---Purpose: Initialize all fields (own and inherited)

    CreatingSoftware (me) returns HAsciiString from TCollection;
	---Purpose: Returns field CreatingSoftware
    SetCreatingSoftware (me: mutable; CreatingSoftware: HAsciiString from TCollection);
	---Purpose: Set field CreatingSoftware

    IntendedAnalysisCode (me) returns HArray1OfAsciiString from TColStd;
	---Purpose: Returns field IntendedAnalysisCode
    SetIntendedAnalysisCode (me: mutable; IntendedAnalysisCode: HArray1OfAsciiString from TColStd);
	---Purpose: Set field IntendedAnalysisCode

    Description (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Description
    SetDescription (me: mutable; Description: HAsciiString from TCollection);
	---Purpose: Set field Description

    AnalysisType (me) returns HAsciiString from TCollection;
	---Purpose: Returns field AnalysisType
    SetAnalysisType (me: mutable; AnalysisType: HAsciiString from TCollection);
	---Purpose: Set field AnalysisType

fields
    theCreatingSoftware: HAsciiString from TCollection;
    theIntendedAnalysisCode: HArray1OfAsciiString from TColStd;
    theDescription: HAsciiString from TCollection;
    theAnalysisType: HAsciiString from TCollection;

end FeaModel;
