-- Created on: 1997-04-14
-- Created by: Olga PILLOT
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class LinearForm from LocOpe 

	---Purpose: Defines a linear form (using Prism from BRepSweep)
	--          with modifications provided for the LinearForm feature.
uses DataMapOfShapeListOfShape from TopTools,
     Edge               from TopoDS,
     Prism            from BRepSweep,     
     Shape           from TopoDS,
     Face            from TopoDS,
     SequenceOfCurve from TColGeom, 
     ListOfShape     from TopTools,
     Curve           from Geom, 
     Vec             from gp,
     Dir             from gp,
     Plane           from Geom,     
     Pnt             from gp
    
raises NoSuchObject from Standard,
       NotDone      from StdFail

is

    Create 
     
    	returns  LinearForm  from  LocOpe;
	---C++: inline

 
    Create (Base  : Shape       from  TopoDS;
    	    V     : Vec         from  gp;
	    Pnt1  : Pnt         from  gp;
	    Pnt2  : Pnt         from  gp)
	    
	---C++: inline
	returns LinearForm from LocOpe;     

    Create (Base  : Shape       from  TopoDS;
    	    V     : Vec         from  gp;
	    Vectra: Vec         from gp;
	    Pnt1  : Pnt         from  gp;
	    Pnt2  : Pnt         from  gp)
	    
	---C++: inline
	returns LinearForm from LocOpe;     

    Perform(me:  in  out;  Base : Shape       from  TopoDS;
		    	   V    : Vec         from  gp;
		           Pnt1 : Pnt         from  gp;
		           Pnt2 : Pnt         from  gp)

	is  static;

    Perform(me:  in  out;  Base  : Shape       from  TopoDS;
		    	   V     : Vec         from  gp;
		    	   Vectra: Vec         from  gp;
		           Pnt1  : Pnt         from  gp;
		           Pnt2  : Pnt         from  gp)

	is  static;

    FirstShape(me)
    
    	returns Shape from TopoDS
	---C++: return const &
	is static;


    LastShape(me)
    
    	returns Shape from TopoDS
	---C++: return const &
	is static;


    Shape(me)
    
    	returns Shape from TopoDS 
	raises  NotDone  from  StdFail
	---C++: return const &
	is static;


    Shapes(me; S: Shape from TopoDS)
    
    	returns ListOfShape from TopTools
	---C++: return const &
    	raises NoSuchObject from Standard
	       -- The exception is raised if S is not a subshape of the profile
	is static;

    IntPerf(me:  in  out) 
     
    	is  static  private;
 

fields

    myBase       : Shape             from TopoDS;
    myVec        : Vec               from gp; 
    myTra        : Vec               from gp; 
    myDone       : Boolean           from Standard; 
    myIsTrans    : Boolean           from Standard;     
    myRes        : Shape             from TopoDS;
    myFirstShape : Shape             from TopoDS;
    myLastShape  : Shape             from TopoDS;
    myMap        : DataMapOfShapeListOfShape    from TopTools;
    myPnt1       : Pnt               from gp;
    myPnt2       : Pnt               from gp;    
    
end LinearForm;     
