-- Created on: 1993-01-09
-- Created by: CKY / Contract Toubro-Larsen (Kiran)
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class CompositeCurve from IGESGeom  inherits IGESEntity

        ---Purpose: defines IGESCompositeCurve, Type <102> Form <0>
        --          in package IGESGeom
        --          A composite curve is defined as an ordered list of entities
        --          consisting of a point, connect point and parametrised curve
        --          entities (excluding the CompositeCurve entity).

uses

        HArray1OfIGESEntity from IGESData

raises OutOfRange

is

        Create returns mutable CompositeCurve;

        -- Specific Methods pertaining to the class

        Init (me          : mutable;
              allEntities : HArray1OfIGESEntity);
         ---Purpose : This method is used to set the fields of the class
         --           CompositeCurve
         --       - allEntities : Constituent Entities of the composite curve

        NbCurves (me) returns Integer;
        ---Purpose : returns the number of curves contained in the CompositeCurve

        Curve (me; Index : Integer) returns IGESEntity
        raises OutOfRange;
        ---Purpose : returns Component of the CompositeCurve (a curve or a point)
        -- raises exception if Index <= 0 or Index > NbCurves()

fields

--
-- Class    : IGESGeom_CompositeCurve
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class CompositeCurve.
--
-- Reminder : A CompositeCurve instance is defined by :
--            The collection of constituent curves which could
--            be of type point, connect point or parametric curve
--            entities

        theEntities : HArray1OfIGESEntity;

end CompositeCurve;
