-- Created on: 2003-08-21
-- Created by: Sergey KUUL
-- Copyright (c) 2003-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class RWReprItemAndLengthMeasureWithUnit from RWStepRepr

	---Purpose : Read & Write Module for ReprItemAndLengthMeasureWithUni

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     ReprItemAndLengthMeasureWithUnit from StepRepr

is

	Create returns RWReprItemAndLengthMeasureWithUnit;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable ReprItemAndLengthMeasureWithUnit from StepRepr);

	WriteStep (me; SW : in out StepWriter; ent : ReprItemAndLengthMeasureWithUnit from StepRepr);

end RWReprItemAndLengthMeasureWithUnit;
