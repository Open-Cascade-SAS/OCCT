-- Created on: 1993-09-22
-- Created by: Didier PIFFAULT
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Vertex from BRepMesh 

  ---Purpose: 


uses    Boolean from Standard,
        Integer from Standard,
        Real from Standard,
        XY from gp,
        DegreeOfFreedom from BRepMesh


is        Create     returns Vertex from BRepMesh;

          Create         (UV      : in XY from gp;
                          Locat3d : in Integer from Standard;
                          Move    : in DegreeOfFreedom from BRepMesh)
            returns Vertex from BRepMesh;


          Create         (U, V    : Real from Standard;
                          Move    : in DegreeOfFreedom from BRepMesh)
            returns Vertex from BRepMesh;


          Initialize     (me      : in out;
                          UV      : in XY from gp; 
                          Locat3d : in Integer from Standard;
                          Move    : in DegreeOfFreedom from BRepMesh)
            is static;


          Coord          (me) 
            returns XY from gp
            ---C++: return const &
            ---C++: inline
            is static;


          Location3d    (me) 
            returns Integer from Standard
            ---C++: inline
            is static;


          Movability     (me)
            returns DegreeOfFreedom from BRepMesh
            ---C++: inline
            is static;

          SetMovability  (me   : in out;
                          Move : DegreeOfFreedom from BRepMesh)
            is static;


          HashCode       (me;
                          Upper : Integer from Standard)
            returns Integer from Standard
            ---C++: function call
            is static;


          IsEqual        (me; Other : Vertex from BRepMesh)
            returns Boolean from Standard
            ---C++: alias operator ==
            is static;


        fields  myUV         : XY from gp;
                myLocation   : Integer from Standard;
                myMovability : DegreeOfFreedom from BRepMesh;

end Vertex;
