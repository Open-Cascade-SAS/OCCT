-- Created on: 1996-12-16
-- Created by: Remi Lequette
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Builder from TNaming  

	---Purpose: A tool to create and maintain topological
    	-- attributes. 
    	-- Constructor creates an empty
    	-- TNaming_NamedShape attribute at the given
    	-- label. It allows adding "old shape" and "new
    	-- shape" pairs with the specified evolution to this
    	-- named shape. One evolution type per one
    	-- builder must be used.
        
uses
    Shape                        from TopoDS,
    Label                        from TDF,
    Data                         from TDF, 
    NamedShape                   from TNaming,	
    PtrNode                      from TNaming,	
    PtrAttribute                 from TNaming,	
    PtrDataMapOfShapePtrRefShape from TNaming
    
raises
    ConstructionError            from Standard
is

	Create (aLabel : Label from TDF) returns Builder from TNaming;
	    ---Purpose:  Create an   Builder.   
	    --  Warning:  Before Addition copies the current Value, and clear 
    	

	---Category: To Load Shape Evolution
	--           =======================
      
    	Generated(me : in out; newShape : Shape from TopoDS);
	    ---Purpose:  Records the shape newShape which was
    	    -- generated during a topological construction.
    	    --  As an example, consider the case of a face
    	    --  generated in construction of a box.
	    
	Generated(me : in out; oldShape, newShape : Shape from TopoDS);
	    ---Purpose: Records the shape newShape which was
    	    --  generated from the shape oldShape during a topological construction.
    	    -- As an example, consider the case of a face
    	    -- generated from an edge in construction of a prism.
    

	---Category: Load Modifications.

	Delete(me : in out; oldShape : Shape from TopoDS);
	    ---Purpose:  Records the shape oldShape which was deleted from the current label.
    	    -- As an example, consider the case of a face removed by a Boolean operation.
	    
	Modify(me : in out; oldShape, newShape : Shape from TopoDS);
	    ---Purpose:  Records the shape newShape which is a
    	    -- modification of the shape oldShape.
    	    -- As an example, consider the case of a face split
    	    --  or merged in a Boolean operation.
	    --          
	
    	---Category: Load Selection.
    	Select (me : in out; aShape, inShape : Shape from TopoDS);
	    ---Purpose:   Add a  Shape to the current label ,  This Shape is
	    --          unmodified.  Used for example  to define a set
	    --          of shapes under a label.
			      

        ---Category: Querying

    	NamedShape(me) returns NamedShape from TNaming;
	    ---Purpose: Returns the NamedShape which has been build or is under construction.

fields
    
    myMap         : PtrDataMapOfShapePtrRefShape from TNaming; 
    myAtt         : PtrAttribute                 from TNaming;
end Builder;
