-- Created on: 1995-03-15
-- Created by: Laurent PAINNOT
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class PolygonOnTriangulation from BRep inherits CurveRepresentation from  BRep


    	---Purpose: A representation by an array of nodes on a 
    	--          triangulation.


uses Location               from TopLoc,
     PolygonOnTriangulation from Poly,
     Triangulation          from Poly


is

    Create(P: PolygonOnTriangulation from Poly;
    	   T: Triangulation          from Poly;
	   L: Location               from TopLoc)
    returns mutable PolygonOnTriangulation from BRep;


    IsPolygonOnTriangulation(me) returns Boolean
    	---Purpose: returns True.
    is redefined;

    IsPolygonOnTriangulation(me; T : Triangulation from Poly;
                            	 L : Location from TopLoc)    returns Boolean
	---Purpose: Is it a polygon in the definition of <T> with
	--          location <L>.
    is redefined;

    PolygonOnTriangulation(me: mutable; P: PolygonOnTriangulation from Poly)
    	---Purpose: returns True.
    is redefined;

    Triangulation(me) returns any Triangulation from Poly
    	---C++: return const&
    is redefined;
    
    PolygonOnTriangulation(me) returns any PolygonOnTriangulation from Poly
    	---C++: return const&
    is redefined;

    
    Copy(me) returns mutable CurveRepresentation from BRep is virtual;
	---Purpose: Return a copy of this representation.


fields

myPolygon       : PolygonOnTriangulation    from Poly;
myTriangulation : Triangulation             from Poly;

end PolygonOnTriangulation;
