-- Created on: 1996-02-16
-- Created by: Philippe MANGIN
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Batten from DrawFairCurve inherits  BSplineCurve2d from DrawTrSurf

	---Purpose: Interactive Draw object of type "Batten"

uses Batten from FairCurve, 
     BSplineCurve2d from DrawTrSurf,
     Pnt2d from gp

is
   Create(TheBatten : Address)
   returns mutable Batten from DrawFairCurve;
   Compute(me:mutable);
   SetPoint(me: mutable; Side : Integer; Point : Pnt2d);
   SetAngle(me: mutable; Side : Integer; Angle : Real);
   SetSliding(me: mutable; Length : Real);
   SetHeight(me: mutable; Heigth : Real);
   SetSlope(me: mutable; Slope : Real);
   GetAngle(me; Side : Integer) returns Real;
   GetSliding(me) returns Real;
   FreeSliding(me:mutable);
   FreeAngle(me:mutable; Side : Integer);
   Dump(me; S : in out OStream)
	---Purpose: For variable dump.
  is redefined;
   
fields
 MyBatten : Address is protected;
end Batten;
