-- File:	RWStepShape_RWSubface.cdl
-- Created:	Fri Jan  4 17:42:45 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class RWSubface from RWStepShape

    ---Purpose: Read & Write tool for Subface

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    Subface from StepShape

is
    Create returns RWSubface from RWStepShape;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : Subface from StepShape);
	---Purpose: Reads Subface

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: Subface from StepShape);
	---Purpose: Writes Subface

    Share (me; ent : Subface from StepShape;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWSubface;
