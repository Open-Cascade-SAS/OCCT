-- Created on: 1993-05-12
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred generic class TopolTool from Contap
           ( TheVertex as any;
             TheArc    as any
           )

inherits TShared from MMgt 

    ---Purpose: Template class for an iterator the restriction of
    --          a surface.

uses Orientation from TopAbs,
     State       from TopAbs,
     Pnt2d       from gp


is

-- Arc iterator

    Init(me: mutable)

    	;


    More(me: mutable)

    	returns Boolean from Standard
    	;


    Value(me: mutable)

    	returns any TheArc
    	;


    Next(me: mutable)

    	;


-- Iterator on the vertex of an arc of restriction


    Initialize(me: mutable; A:TheArc);


    InitVertexIterator(me: mutable)

    	;


    MoreVertex(me: mutable)

    	returns Boolean from Standard
    	;



    Vertex(me: mutable)
    	returns any TheVertex
    	;


    NextVertex(me: mutable)

    	;


    Orientation(me: mutable; A: TheArc)
    
    	returns Orientation from TopAbs;


    Orientation(me: mutable; V: TheVertex)
    
    	returns Orientation from TopAbs;


    Identical(me: mutable; V1,V2: TheVertex)
    
	---Purpose: Returns True if the vertices V1 and V2 are identical.
	--          This method does not take the orientation of the
	--          vertices in account.

    	returns Boolean from Standard;


    Classify(me: mutable; P: Pnt2d from gp; Tol: Real from Standard)
    
    	returns State from TopAbs;


end TopolTool;

