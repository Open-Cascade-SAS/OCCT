-- Created on: 1991-03-07
-- Created by: Denis Pascal
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package GraphTools 

    ---Purpose: This package <GraphTools> provides  algorithms working
    --          on a directed graph.  Those algorithms are generic for
    --          user (Graph and Vertex)  data, and tool classes.


uses Standard,
     MMgt,
     TCollection,
     TColStd
     
is


    class ListOfSequenceOfInteger instantiates List from TCollection
                         (SequenceOfInteger from TColStd);

-- Requirements
-- ============

-- Data
--  Vertex
--  Graph
-- Tools
    generic class GraphIterator;
    generic class VertexIterator;

-- Services (Algorithms) 
-- =====================
    
    
    ---Purpose: Depth First Search (DFS)
    
    generic class DFSIterator,
                  DFSMap;


    ---Purpose: Breath First Search (BFS)

    generic class BFSIterator,
                  BFSMap;

		  
    ---Purpose: Sorted Strong Components (SC)

    generic class SortedStrgCmptsFromIterator,
                  SCMap;
		  
    generic class SortedStrgCmptsIterator;


    ---Purpose: Topological Sort (TS)

    class TSNode;

    generic class TopologicalSortFromIterator,
                  TSMap;  
		  
    generic class TopologicalSortIterator;
    
    
    ---Purpose: Connected Vertices (CV)

    generic class ConnectedVerticesFromIterator,
                  CVMap,
    	    	  ConnectMap;
		 
    generic class ConnectedVerticesIterator;


    ---Purpose: Reduced Graph (RG)
    
    class RGNode;
    
    class SC;
    
    class SCList instantiates List from TCollection
                (SC from GraphTools);

    generic class ReducedGraph,
		  RGMap,
		  SortedSCIterator,
		  AdjSCIterator;

end GraphTools;





