-- Created on: 1994-04-05
-- Created by: Yves FRICAUD
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

private class FunctionInter from Bisector  
inherits FunctionWithDerivative from math 

        ---Purpose:                           2                      2 
	--          F(u) =  (PC(u) - PBis1(u))   + (PC(u) - PBis2(u))

uses 
    Curve   from Geom2d,
    Curve   from Bisector
	--          

is

    Create  returns FunctionInter from Bisector;
    
    Create (C     : Curve   from Geom2d ;
            Bis1  : Curve   from Bisector;
	    Bis2  : Curve   from Bisector)  
    returns FunctionInter from Bisector;
    
    Perform (me    : in out;
    	     C     : Curve   from Geom2d ;
             Bis1  : Curve   from Bisector;
	     Bis2  : Curve   from Bisector)
    is static;	     	
	     
    Value(me : in out; X : Real; F : out Real) 
    	---Purpose: Computes the values of the Functions for the variable <X>.
    returns Boolean
    is static;
    
    Derivative(me : in out; X : Real; D : out Real) 
    returns Boolean;

    Values(me : in out ; X  : Real; F  : out Real; D  : out Real)    
    	---Purpose: Returns the values of the functions and the derivatives
    	--          for the variable <X>.
    returns Boolean
    is static;
    
fields
    
    curve     : Curve from Geom2d;
    bisector1 : Curve from Bisector;
    bisector2 : Curve from Bisector;
    
end FunctionInter;
