-- Created on: 2003-06-04
-- Created by: Galina KULIKOVA
-- Copyright (c) 2003-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class DatumReference from StepDimTol
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity DatumReference

uses
    Datum from StepDimTol

is
    Create returns DatumReference from StepDimTol;
	---Purpose: Empty constructor

    Init (me: mutable; aPrecedence: Integer;
                       aReferencedDatum: Datum from StepDimTol);
	---Purpose: Initialize all fields (own and inherited)

    Precedence (me) returns Integer;
	---Purpose: Returns field Precedence
    SetPrecedence (me: mutable; Precedence: Integer);
	---Purpose: Set field Precedence

    ReferencedDatum (me) returns Datum from StepDimTol;
	---Purpose: Returns field ReferencedDatum
    SetReferencedDatum (me: mutable; ReferencedDatum: Datum from StepDimTol);
	---Purpose: Set field ReferencedDatum

fields
    thePrecedence: Integer;
    theReferencedDatum: Datum from StepDimTol;

end DatumReference;
