-- Created on: 1992-11-17
-- Created by: Christian CAILLET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



deferred class SelectCombine  from IFSelect  inherits Selection

    ---Purpose : A SelectCombine type Selection defines algebraic operations
    --           between results of several Selections
    --           It is a deferred class : sub-classes will have to define
    --           precise what operator is to be applied

uses AsciiString from TCollection, EntityIterator,
     Graph, SelectionIterator, TSeqOfSelection

is

    Initialize;
    ---Purpose : Defines an empty SelectCombine

    NbInputs (me) returns Integer;
    ---Purpose : Returns the count of Input Selections

    Input (me; num : Integer) returns mutable Selection;
    ---Purpose : Returns an Input Selection, given its rank in the list

    InputRank (me; sel : Selection) returns Integer;
    ---Purpose : Returns the rank of an input Selection, 0 if not in the list.
    --           Most generally, its value is meaningless, except for testing
    --           the presence of an input Selection :
    --           - == 0  if <sel> is not an input for <me>
    --           - >  0  if <sel> is an input for <me>

    Add (me : mutable; sel : mutable Selection; atnum : Integer = 0);
    ---Purpose : Adds a Selection to the filling list
    --           By default, adds it to the end of the list
    --           A Positive rank less then NbInputs gives an insertion rank
    --           (InsertBefore : the new <atnum>th item of the list is <sel>)

    Remove (me : mutable; sel : Selection) returns Boolean;
    ---Purpose : Removes an input Selection.
    --           Returns True if Done, False, if <sel> is not an input for <me>

    Remove (me : mutable; num : Integer) returns Boolean;
    ---Purpose : Removes an input Selection, given its rank in the list
    --           Returns True if Done, False if <num> is out of range


    HasUniqueResult (me) returns Boolean  is redefined protected;
    ---Purpose : Returns always True, because RootResult gives a Unique list


    FillIterator (me; iter : in out SelectionIterator);
    ---Purpose : Puts in an Iterator the Selections from which "me" depends
    --           That is to say, the list of Input Selections

fields

    thelist : TSeqOfSelection;

end SelectCombine;
