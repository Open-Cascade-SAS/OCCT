-- Created on: 1991-07-24
-- Created by: Michel CHAUVAT
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



private generic class FuncExtPC from Extrema 
(Curve    as any;
 Tool     as any;
 POnC     as any;
 Pnt      as any;
 Vec      as any)
						     
    inherits FunctionWithDerivative from math
    --- Purpose: Function to find extrema of the distance between a
    --- point and a curve.

uses    SequenceOfReal    from TColStd,
	SequenceOfInteger from TColStd
	
raises  OutOfRange   from Standard,
        TypeMismatch from Standard

private class SeqPC instantiates Sequence from TCollection(POnC);	


is

    Create returns FuncExtPC;

    Create (P: Pnt; C: Curve) returns FuncExtPC;
    	---Purpose: 

    Initialize(me: in out; C: Curve)
    	---Purpose: sets the field mycurve of the function.
    is static;
    
    SetPoint(me: in out; P: Pnt)
    	---Purpose: sets the field P of the function.
    is static;


    -- In all next methods, an exception is raised if the fields 
    -- were not initialized.

    Value (me: in out; U: Real; F: out Real) returns Boolean;
    	---Purpose: Calculation of F(U).

    Derivative (me: in out; U: Real; DF: out Real) returns Boolean;
    	---Purpose: Calculation of F'(U).

    Values (me: in out; U: Real; F,DF: out Real) returns Boolean;
    	---Purpose: Calculation of F(U) and F'(U).

    GetStateNumber (me: in out) returns Integer
    	---Purpose: Save the found extremum.
    	is redefined;

    NbExt (me) returns Integer
    	---Purpose: Return the nunber of found extrema.
    raises TypeMismatch from Standard;

    SquareDistance (me; N: Integer) returns Real
    	---Purpose: Returns the Nth distance.
    	raises  OutOfRange from Standard,
                TypeMismatch from Standard;
	    	-- if N < 1 or N > NbExt(me).

    IsMin (me; N: Integer) returns Boolean
    	---Purpose: Shows if the Nth distance is a minimum.
    	raises  OutOfRange from Standard,
                TypeMismatch from Standard;
	    	-- if N < 1 or N > NbExt(me).

    Point (me; N: Integer) returns POnC
    	---Purpose: Returns the Nth extremum.
    	raises  OutOfRange from Standard,
                TypeMismatch from Standard;
	    	-- if N < 1 or N > NbExt(me).

    SubIntervalInitialize(me: in out; theUfirst, theUlast: Real from Standard);
    	---Purpose: Determines boundaries of subinterval for find of root.
    
    SearchOfTolerance(me: in out) returns Real from Standard;
    	---Purpose: Computes a Tol value. If 1st derivative of curve
    	--          |D1|<Tol, it is considered D1=0.      
    

fields
    myP    : Pnt;
    myC    : Address from Standard;

    myU    : Real;          -- current
    myPc   : Pnt;           -- current point 
    myD1f  : Real;          -- value of derivative of the function

    mySqDist: SequenceOfReal    from TColStd;
    myIsMin: SequenceOfInteger from TColStd;
    myPoint: SeqPC;
    myPinit: Boolean;
    myCinit: Boolean;
    myD1Init: Boolean;
    
    myTol: Real from Standard;  -- toolerance for derivate

--Supremum of search 1st non-zero derivative    
    myMaxDerivOrder: Integer from Standard;
    
--boundaries of subinterval for find of root
    myUinfium, myUsupremum: Real from Standard;
    

end FuncExtPC;
