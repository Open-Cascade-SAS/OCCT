-- Created on: 1992-09-18
-- Created by: Jean Louis FRENKEL
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Drawer from Prs3d inherits TShared from MMgt

	---Purpose: A graphic attribute manager which governs how
    	-- objects such as color, width, line thickness and
    	-- deflection are displayed.
    	-- Prs3d_Drawer is the mother class of AIS_Drawer.
    	-- As such, it is its set functions which are called to
    	-- modify display parameters. In the example below we
    	-- can see that the AIS_Drawer is modified to set the
    	-- value of the deviation coefficient using a method
    	-- inherited from Prs3d_Drawer.
	
uses
    DatumAspect from Prs3d,
    LineAspect from Prs3d,
    TextAspect from Prs3d,
    PointAspect from Prs3d,
    ShadingAspect from Prs3d,
    IsoAspect from Prs3d,
    DimensionAspect from Prs3d,
    PlaneAspect from Prs3d,
    ArrowAspect from Prs3d,
    TypeOfDeflection from Aspect,
    NameOfColor from Quantity,
    PlaneAngle from Quantity,
    Length from Quantity,
    TypeOfHLR from Prs3d

is
    Create returns mutable Drawer from Prs3d;

---Category: deviation definition.
-- 
-- All drawings of curves or patches are made with respect to a maximal 
-- chordial deviation. This deviation is absolute and given through
-- the method: SetMaximalChordialDeviation.
-- 
-- In the case of drawing shapes, it is allowed to ask for a relative
-- deviation.
-- This deviation will be: SizeOfObject * DeviationCoefficient where
-- DeviationCoefficient can be set through the method: SetDeviationCoefficient.
-- 
--
-- For drawing algorithms using discretisation, a default number of
-- points has been set to 17. It is possible to use the method SetDiscret
-- to change this number.
--


    SetTypeOfDeflection (me:mutable; 
    	                aTypeOfDeflection: TypeOfDeflection from  Aspect)  
    	---Purpose: Sets the type of chordal deflection.
    	-- This indicates whether the deflection value is absolute
    	-- or relative to the size of the object.         
    is virtual;
    
    TypeOfDeflection(me) returns TypeOfDeflection from Aspect
    is virtual;
    	--- Purpose: Returns the type of chordal deflection.
    	-- This indicates whether the deflection value is absolute
    	-- or relative to the size of the object.   
    
    SetMaximalChordialDeviation (me: mutable; 
    	    	    	       aChordialDeviation: Length from Quantity)
    	---Purpose: Defines the maximal chordial deviation when drawing any curve;
    	--          Even if the type of deviation is set to TOD_Relative,
    	--          this value is used by:
    	--          
    	--                   Prs3d_DeflectionCurve
    	--                   Prs3d_WFDeflectionSurface
    	--                   Prs3d_WFDeflectionRestrictedFace
    is virtual;
    
    MaximalChordialDeviation (me) returns Length from Quantity
    	---Purpose: returns the maximal chordial deviation. Default value is 0.1
    is virtual;
	    
    SetDeviationCoefficient(me: mutable; aCoefficient: Real from Standard)
    	---Purpose: Sets the deviation coefficient aCoefficient.
    is virtual;

    DeviationCoefficient(me) returns Real from Standard 
    is virtual;
    	---Purpose: Returns the deviation coefficient.
    SetHLRDeviationCoefficient(me: mutable; aCoefficient: Real from Standard)
    	---Purpose: Sets the deviation coefficient aCoefficient for removal
    	-- of hidden lines created by different viewpoints in
    	-- different presentations. The Default value is 0.02.
    is virtual;

    HLRDeviationCoefficient(me) returns Real from Standard 
    is virtual;
    	---Purpose: Returns the real number value of the hidden line
    	-- removal deviation coefficient.   
    SetHLRAngle(me: mutable; anAngle: Real from Standard)
	---Purpose: Sets anAngle, the angle of maximum chordal
    	-- deviation for removal of hidden lines created by
    	-- different viewpoints in different presentations. The
    	-- default value is 20*PI/180.
    is virtual;

    HLRAngle(me) returns Real from Standard 
    is virtual;
    	---Purpose: Returns the real number value of the deviation angle
    	-- in hidden line removal views. The default value is 20*PI/180.
    
    SetDeviationAngle(me: mutable; anAngle: Real from Standard)
	---Purpose: Sets deviation angle
    is virtual;

    DeviationAngle(me) returns Real from Standard
    	---Purpose: Returns the value for deviation angle.
    is virtual;

    SetDiscretisation(me: mutable; d: Integer from Standard)
    	---Purpose: Sets the discretisation parameter d.
    is virtual;

    Discretisation(me) returns Integer from Standard
    is virtual;
    	---Purpose: Returns the discretisation setting.
    SetMaximalParameterValue(me: mutable; Value: Real from Standard)
    	---Purpose: defines the maximum value allowed  for the first and last
	--          parameters of an infinite curve. Default value: 500. 
    is virtual;
    
    MaximalParameterValue(me) returns Real from Standard
    is virtual;
    	--- Purpose: Sets the maximum value allowed for the first and last
    	-- parameters of an infinite curve. By default, this value is 500000. 

    SetIsoOnPlane (me: mutable; OnOff: Boolean from Standard)
    	---Purpose: Sets IsoOnPlane on or off   by setting the parameter
    	-- OnOff to true or false.
    is virtual;
    
    IsoOnPlane(me) returns Boolean from Standard 
	---Purpose: Returns True if the drawing of isos on planes is enabled.
    is virtual;
    
    SetTypeOfHLR(me: mutable; theTypeOfHLR: TypeOfHLR from Prs3d)
    is virtual;
    ---Purpose: Sets the type of HLR algorithm
    --          used by drawer's interactive objects
    
    TypeOfHLR(me) returns TypeOfHLR from Prs3d
    is virtual;
     ---Purpose: Gets the myTypeOfHLR value


-- 
-- Attributes for the U Isoparametric lines of patches.
--    
    UIsoAspect (me:mutable) returns mutable IsoAspect from Prs3d
    	---Purpose: Defines the attributes which are used when drawing an 
    	--          U isoparametric curve of a face. Defines the number
    	--          of U isoparametric curves to be drawn for a single face.
    	--          The LineAspect for U isoparametric lines can be edited
    	--          (methods SetColor, SetTypeOfLine, SetWidth, SetNumber)
    	--          The default values are:
    	--          COLOR       : Quantity_NOC_GRAY75
    	--          TYPE OF LINE: Aspect_TOL_SOLID
    	--          WIDTH       : 0.5
    	--          
    	--         
    	--          These attributes are used by the following algorithms:
    	--          Prs3d_WFDeflectionSurface 
    	--          Prs3d_WFDeflectionRestrictedFace


    is virtual;    
    
    SetUIsoAspect (me:mutable; anAspect: IsoAspect from Prs3d) 
    is virtual;

-- Attributes for the V Isoparametric line of patches.


    VIsoAspect (me:mutable) returns mutable IsoAspect from Prs3d
    	---Purpose: Defines the attributes which are used when drawing an 
    	--          V isoparametric curve of a face. Defines the number
    	--          of V isoparametric curves to be drawn for a single face.
    	--          The LineAspect for V isoparametric lines can be edited
    	--          (methods SetColor, SetTypeOfLine, SetWidth, SetNumber)
    	--          The default values are:
    	--          COLOR       : Quantity_NOC_GRAY82
    	--          TYPE OF LINE: Aspect_TOL_SOLID
    	--          WIDTH       : 0.5
    	--          
    	--         
    	--          These attributes are used by the following algorithms:
    	--          Prs3d_WFDeflectionSurface 
    	--          Prs3d_WFDeflectionRestrictedFace
    is virtual;    
    
    SetVIsoAspect (me:mutable;anAspect: IsoAspect from Prs3d)
    is virtual;
    	---Purpose: Sets the appearance of V isoparameters - anAspect.

    FreeBoundaryAspect (me:mutable) returns mutable LineAspect from Prs3d
    	---Purpose:  Stores the values for presentation of free boundaries,
    	-- in other words, boundaries which are not shared.
	--          The LineAspect for the  free boundaries can be edited.
	--          The default values are:
	--          Color: Quantity_NOC_GREEN
	--          Type of line: Aspect_TOL_SOLID
	--          Width: 1.
	--          These attributes are used by the algorithm Prs3d_WFShape
    is virtual;
    
    SetFreeBoundaryAspect(me:mutable;anAspect: LineAspect from Prs3d)
    is virtual;
    	--- Purpose: Sets the parameter anAspect for the display of free boundaries.
    
    SetFreeBoundaryDraw (me: mutable; OnOff: Boolean from Standard)
    	---Purpose: Sets free boundary drawing on or off by setting the
    	-- parameter OnOff to true or false.
    
    is virtual;
    
    FreeBoundaryDraw(me) returns Boolean from Standard 
    	---Purpose: Returns True if the drawing of the shared boundaries
    	-- is disabled. True is the default setting.
    is virtual;
    

-- Attributes for the wires

    WireAspect (me:mutable) returns mutable LineAspect from Prs3d
    	---Purpose: Returns wire aspect settings.
    	--          The LineAspect for the wire can be edited.
    	--          The default values are:
    	--          Color: Quantity_NOC_RED
    	--          Type of line: Aspect_TOL_SOLID
    	--          Width: 1.           
    	--          These attributes are used by the algorithm Prs3d_WFShape
    is virtual;    

    SetWireAspect(me:mutable;anAspect: LineAspect from Prs3d)
    is virtual;

    	--- Purpose: Sets the parameter anAspect for display of wires.
        
    SetWireDraw (me: mutable; OnOff: Boolean from Standard)
    	---Purpose: Sets WireDraw on or off   by setting the parameter
    	-- OnOff to true or false.
    
    is virtual;
    
    WireDraw(me) returns Boolean from Standard 
    	---Purpose: returns True if the drawing of the wire is enabled.
    is virtual;
    

-- Attributes for the unfree boundaries

    UnFreeBoundaryAspect (me:mutable) returns mutable LineAspect from Prs3d
    	---Purpose: Returns settings for shared boundary line aspects.
    	--          The LineAspect for the unfree boundaries can be edited.
    	--          The default values are:
    	--          Color: Quantity_NOC_YELLOW
    	--          Type of line: Aspect_TOL_SOLID
    	--          Width: 1.
    	--          These attributes are used by the algorithm Prs3d_WFShape
    is virtual;

    SetUnFreeBoundaryAspect(me:mutable; anAspect: LineAspect from Prs3d)
    is virtual;
    	--- Purpose: Sets the parameter anAspect for the display of shared boundaries.   
    SetUnFreeBoundaryDraw (me: mutable; OnOff: Boolean from Standard)
    	---Purpose: Sets FreeBoundaryDraw on or off by setting the
    	-- parameter OnOff to true or false.
        --          By default the unfree boundaries  are drawn.
    
    is virtual;
    
    UnFreeBoundaryDraw(me) returns Boolean from Standard 
    	---Purpose: Returns True if the drawing of the shared boundaries is enabled.
    	-- True is the default setting.
    is virtual;
    

-- 
--  Attributes for the lines.
-- 

    LineAspect(me:mutable) returns mutable LineAspect from Prs3d
    	---Purpose:   Returns settings for line aspects.
    	-- These settings can be edited. The default values are:       
    	--          Color: Quantity_NOC_YELLOW
    	--          Type of line: Aspect_TOL_SOLID
    	--          Width: 1.
    	--          These attributes are used by the following algorithms:
    	--          Prs3d_Curve
    	--          Prs3d_Line
    	--          Prs3d_HLRShape

    is virtual;
    
    SetLineAspect(me:mutable; anAspect: LineAspect from Prs3d)
    is virtual;
    	--- Purpose: Sets the parameter anAspect for display attributes of lines.

    TextAspect(me:mutable) returns mutable TextAspect from Prs3d
    	--- Purpose: Returns settings for text aspect.
    	-- These settings can be edited. The default value is:
    	-- -   Color: Quantity_NOC_YELLOW
  
    is virtual;
    
    SetTextAspect(me:mutable; anAspect: TextAspect from Prs3d)
    is virtual;
    	--- Purpose: Sets the parameter anAspect for display attributes of text.   
    
    SetLineArrowDraw (me: mutable; OnOff: Boolean from Standard)
    	---Purpose: enables the drawing of an arrow at the end of each line.
    	--          By default the arrows are not drawn.
    
    is virtual;
    
    LineArrowDraw(me) returns Boolean from Standard 
    	---Purpose: Sets LineArrowDraw on or off by setting the
    	-- parameter OnOff to true or false.
    is virtual;
    
    ArrowAspect(me:mutable) returns mutable ArrowAspect from Prs3d 
    is virtual;
    	---Purpose: Returns the attributes for display of arrows.    
    
    SetArrowAspect(me:mutable; anAspect: ArrowAspect from Prs3d)
    is virtual ;
    	---Purpose: Sets the parameter anAspect for display attributes of arrows.
        
    PointAspect(me:mutable) returns mutable PointAspect from Prs3d
    	---Purpose: Returns the point aspect setting. The default values are
    	--        Color: Quantity_NOC_YELLOW
    	--          Type of marker: Aspect_TOM_PLUS
    	--          Scale: 1.          
	--          These attributes are used by the algorithms Prs3d_Point.
    is virtual;
    
    SetPointAspect(me:mutable; anAspect: PointAspect from Prs3d) 
    is virtual;
    	--- Purpose: Sets the parameter anAspect for display attributes of points
        
    ShadingAspect (me:mutable) returns mutable ShadingAspect from Prs3d
   is virtual;
    	---Purpose: Returns settings for shading aspects.
    	-- These settings can be edited. The default values are:
    	-- -   Color: Quantity_NOC_YELLOW
    	-- -   Material: Graphic3d_NOM_BRASS
    	--   Shading aspect is obtained through decomposition of
    	-- 3d faces into triangles, each side of each triangle
    	-- being a chord of the corresponding curved edge in
    	-- the face. Reflection of light in each projector
    	-- perspective is then calculated for each of the
    	-- resultant triangular planes.
    

    SetShadingAspect(me:mutable; anAspect: ShadingAspect from Prs3d) 
    is virtual;
    	---Purpose: Sets the parameter anAspect for display attributes of shading.
        
    SetShadingAspectGlobal(me: mutable; aValue: Boolean from Standard) 
    	---Purpose: indicates that the ShadingAspect will be apply
    	--          to the whole presentation. This allows to modify
    	--          the aspect without recomputing the content of the presentation.
    is virtual;
    
    ShadingAspectGlobal(me) returns Boolean from Standard
    is virtual;  
--
--  Attributes for hidden lines removal. These attributes are used when
--  using an algorithm such Prs3d_HLRShape for example.
--  

    DrawHiddenLine(me) returns Boolean from Standard 
    	---Purpose: returns Standard_True if the hidden lines are to be drawn.
    	--          By default the hidden lines are not drawn.
    is virtual;
    
    EnableDrawHiddenLine(me: mutable)
    	---Purpose: Enables the DrawHiddenLine function.
    is virtual;

    DisableDrawHiddenLine(me: mutable)
    	---Purpose:  Disables the DrawHiddenLine function.
    is virtual;

    HiddenLineAspect(me:mutable) returns mutable LineAspect from Prs3d
    	---Purpose: Returns settings for hidden line aspects.
    	-- These settings can be edited. The default values are:
    	--          Color: Quantity_NOC_YELLOW
    	--          Type of line: Aspect_TOL_DASH
	--          Width: 1.
    is virtual;

    SetHiddenLineAspect(me:mutable; anAspect: LineAspect from Prs3d) 
    is virtual;
    	---Purpose: Sets the parameter anAspect for the display of
    	-- hidden lines in hidden line removal mode.   
    
    SeenLineAspect(me:mutable) returns mutable LineAspect from Prs3d
	---Purpose: Returns settings for seen line aspects.
    	-- These settings can be edited. The default values are:
	--          Color: Quantity_NOC_YELLOW
    	--          Type of line: Aspect_TOL_SOLID
    	--          Width: 1.
    is virtual;

    SetSeenLineAspect(me:mutable; anAspect: LineAspect from Prs3d) 
    is virtual;
    	--- Purpose: Sets the parameter anAspect for the display of seen
    	-- lines in hidden line removal mode.

    PlaneAspect(me:mutable) returns mutable PlaneAspect from Prs3d
    is virtual;
    	---Purpose: Returns settings for the appearance of planes.
    
    SetPlaneAspect(me:mutable; anAspect: PlaneAspect from Prs3d)
    is virtual;
    	---Purpose: Sets the parameter anAspect for the display of planes.

    VectorAspect(me:mutable) returns mutable LineAspect from Prs3d
    	---Purpose: Returns settings for the appearance of vectors.
    	-- These settings can be edited. The default values are:
    	--          Color: Quantity_NOC_SKYBLUE
    	--          Type of line: Aspect_TOL_SOLID
    	--          Width: 1.
    is virtual;

    SetVectorAspect(me:mutable; anAspect: LineAspect from Prs3d) 
    is virtual;
    	---Purpose: Sets the modality anAspect for the display of vectors.    

--
--  Attributes for the presentation of a Datum.
--  

    DatumAspect(me:mutable) returns mutable DatumAspect from Prs3d
    	---Purpose: Returns settings for the appearance of datums.
    	-- These settings can be edited. The default values for
    	-- the three axes are:
    	--          Color: Quantity_NOC_PEACHPUFF
    	--          Type of line: Aspect_TOL_SOLID
    	--          Width: 1.
    is virtual;

    SetDatumAspect(me:mutable; anAspect: DatumAspect from Prs3d)
    is virtual;
    	---Purpose: Sets the modality anAspect for the display of datums.

    DimensionAspect(me:mutable) returns mutable DimensionAspect from Prs3d
    	---Purpose: Returns settings for the appearance of dimensions.
    is virtual;

    SetDimensionAspect(me:mutable; theAspect: DimensionAspect from Prs3d) 
    is virtual;
    	---Purpose: Sets the modality anAspect for display of dimensions.

    SectionAspect (me:mutable) returns mutable LineAspect from Prs3d
    	---Purpose: The LineAspect for the wire can be edited.
    	--          The default values are:
    	--          Color: Quantity_NOC_ORANGE
    	--          Type of line: Aspect_TOL_SOLID
    	--          Width: 1.
       	--          These attributes are used by the algorithm Prs3d_WFShape
    is virtual;    

    SetSectionAspect(me:mutable;anAspect: LineAspect from Prs3d)
    is virtual;
    	---Purpose: Sets the parameter anAspect for display attributes of sections.
    
    SetFaceBoundaryDraw (me           : mutable;
                         theIsEnabled : Boolean from Standard)
    is virtual;
        ---Purpose: Enables or disables face boundary drawing for shading presentations.
        -- theIsEnabled is a boolean flag indicating whether the face boundaries should be
        -- drawn or not.

    IsFaceBoundaryDraw (me) returns Boolean from Standard
    is virtual;
        ---Purpose: Checks whether the face boundary drawing is enabled or not.

    SetFaceBoundaryAspect (me        : mutable;
                           theAspect : LineAspect from Prs3d)
    is virtual;
        ---Purpose: Sets line aspect for face boundaries.
        -- theAspect is the line aspect that determines the look of the face boundaries.

    FaceBoundaryAspect (me : mutable) returns mutable LineAspect from Prs3d
    is virtual;
        ---Purpose: Returns line aspect of face boundaries.

fields
            myUIsoAspect: IsoAspect from Prs3d is protected;
            myVIsoAspect: IsoAspect from Prs3d is protected;
	    myNbPoints  : Integer   from Standard is protected;
	    myIsoOnPlane: Boolean from Standard is protected;
	    myFreeBoundaryAspect: LineAspect from Prs3d is protected;
            myFreeBoundaryDraw: Boolean from Standard is protected;
	    myUnFreeBoundaryAspect: LineAspect from Prs3d is protected;
            myUnFreeBoundaryDraw: Boolean from Standard is protected;
	    myWireAspect: LineAspect from Prs3d is protected;
            myWireDraw: Boolean from Standard is protected;
	    myLineAspect: LineAspect from Prs3d is protected;
	    myTextAspect: TextAspect from Prs3d is protected;
            myShadingAspect: ShadingAspect from Prs3d is protected;
            myShadingAspectGlobal: Boolean from Standard is protected;
            myChordialDeviation: Length from Quantity is protected;
	    myTypeOfDeflection: TypeOfDeflection from Aspect is protected;
            myMaximalParameterValue: Real from Standard is protected;
	    
            myDeviationCoefficient: Real from Standard is protected;
            myHLRDeviationCoefficient: Real from Standard is protected;

	    myDeviationAngle: Real from Standard is protected;
	    myHLRAngle:       Real from Standard is protected;
	    
            myPointAspect: PointAspect from Prs3d is protected;
            myPlaneAspect: PlaneAspect from Prs3d is protected;
            myArrowAspect: ArrowAspect from Prs3d is protected;
            myLineDrawArrow: Boolean from Standard is protected;
	    myDrawHiddenLine: Boolean from Standard is protected;
	    myHiddenLineAspect: LineAspect from Prs3d is protected;
	    mySeenLineAspect: LineAspect from Prs3d is protected;
            myVectorAspect: LineAspect from Prs3d is protected;
            myDatumAspect: DatumAspect from Prs3d is protected;
	    myDatumScale: Real from Standard is protected;
	    myDimensionAspect: DimensionAspect from Prs3d is protected;
      mySectionAspect: LineAspect from Prs3d is protected;
      myFaceBoundaryDraw    : Boolean from Standard is protected;
      myFaceBoundaryAspect  : LineAspect from Prs3d is protected;
      myTypeOfHLR           : TypeOfHLR from Prs3d is protected;
end Drawer;
