-- Created on: 1998-01-17
-- Created by: Julia GERASIMOVA
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class EqualRadiusRelation from AIS inherits Relation from AIS 

	---Purpose: 

uses
    Edge from TopoDS,
    Plane from Geom,
    PresentationManager3d from PrsMgr,
    Presentation from Prs3d,
    Projector from Prs3d,
    Transformation        from Geom,
    Selection from SelectMgr,
    Pnt from gp
    
is
    Create( aFirstEdge  : Edge from TopoDS;
    	    aSecondEdge : Edge from TopoDS; 
	    aPlane      : Plane from Geom ) 
	    ---Purpose: Creates equal relation of two arc's radiuses.
	    --          If one of edges is not in the given plane,
    	    --	        the presentation method projects it onto the plane.
    returns mutable EqualRadiusRelation from AIS;
   
-- Methods from PresentableObject

    Compute( me            : mutable;
  	     aPresentationManager: PresentationManager3d from PrsMgr;
    	     aPresentation : mutable Presentation from Prs3d;
    	     aMode         : Integer from Standard= 0 ) 
    is redefined static private;
    
    Compute( me            : mutable;
    	     aProjector    : Projector from Prs3d;
             aPresentation : mutable Presentation from Prs3d )
    is redefined static private;
    
    Compute(me            : mutable;
    	    aProjector    : Projector from Prs3d;
    	    aTrsf         : Transformation from Geom;
	    aPresentation : mutable Presentation from Prs3d)
    is redefined;
    	---Purpose: computes the presentation according to a point of view
    	--          given by <aProjector>. 
   	--          To be Used when the associated degenerated Presentations 
   	--          have been transformed by <aTrsf> which is not a Pure
    	--          Translation. The HLR Prs can't be deducted automatically
    	--          WARNING :<aTrsf> must be applied
    	--          to the object to display before computation  !!!

-- Methods from SelectableObject

    ComputeSelection( me         : mutable;
    	    	      aSelection : mutable Selection from SelectMgr;
    	    	      aMode      : Integer from Standard)
    is private;
    
    ComputeRadiusPosition(me: mutable) is private;

fields
    
    myFirstCenter  : Pnt from gp;
    mySecondCenter : Pnt from gp;
    myFirstPoint   : Pnt from gp;
    mySecondPoint  : Pnt from gp;

end EqualRadiusRelation;
