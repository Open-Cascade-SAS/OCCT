-- Created on: 1996-02-13
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class GTool from TopOpeBRepBuild

uses

    GTopo from TopOpeBRepBuild,
    ShapeEnum from TopAbs,
    OStream from Standard
    
is

    GFusUnsh(myclass; s1,s2 : ShapeEnum from TopAbs) returns GTopo;
    GFusSame(myclass; s1,s2 : ShapeEnum from TopAbs) returns GTopo;
    GFusDiff(myclass; s1,s2 : ShapeEnum from TopAbs) returns GTopo;

    GCutUnsh(myclass; s1,s2 : ShapeEnum from TopAbs) returns GTopo;
    GCutSame(myclass; s1,s2 : ShapeEnum from TopAbs) returns GTopo;
    GCutDiff(myclass; s1,s2 : ShapeEnum from TopAbs) returns GTopo;

    GComUnsh(myclass; s1,s2 : ShapeEnum from TopAbs) returns GTopo;
    GComSame(myclass; s1,s2 : ShapeEnum from TopAbs) returns GTopo;
    GComDiff(myclass; s1,s2 : ShapeEnum from TopAbs) returns GTopo;

    Dump(myclass; OS : in out OStream from Standard);
    
end GTool;
