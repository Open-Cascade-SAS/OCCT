-- Created on: 1998-04-07
-- Created by: Jean-Pierre COMBE
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class PositionStorageDriver from MPrsStd inherits ASDriver from MDF

	---Purpose: 

uses SRelocationTable from MDF,
     Attribute        from TDF,
     Attribute        from PDF, 
     MessageDriver    from CDM


is

    Create(theMessageDriver : MessageDriver from CDM)  
    returns mutable PositionStorageDriver from MPrsStd;


    VersionNumber(me) returns Integer from Standard;
	---Purpose: Returns the version number from which the driver
	--          is available: 0.

    SourceType(me) returns Type from Standard;
	---Purpose: Returns the type: ColorAttribute from TGraphicAttribute.

    NewEmpty (me) returns mutable Attribute from PDF;


    Paste(me;
    	  Source     :         Attribute from TDF;
    	  Target     : mutable Attribute from PDF;
    	  RelocTable : SRelocationTable from MDF);


end PositionStorageDriver;

