-- Created on: 1995-12-04
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.





package RWStepBasic 

uses

	StepData, Interface, TCollection, TColStd, StepBasic

is


--class ReadWriteModule;

--class GeneralModule;

class RWAddress;
class RWApplicationContext;
class RWApplicationContextElement;
class RWApplicationProtocolDefinition;
class RWApproval;
class RWApprovalPersonOrganization;
class RWApprovalRelationship;
class RWApprovalRole;
class RWApprovalStatus;
class RWCalendarDate;
class RWConversionBasedUnit;
class RWCoordinatedUniversalTimeOffset;
class RWDate;
class RWDateAndTime;
class RWDateRole;
class RWDateTimeRole;
class RWDimensionalExponents;
class RWLengthMeasureWithUnit;
class RWLengthUnit;
class RWLocalTime;
class RWMeasureWithUnit;
class RWNamedUnit;
class RWOrdinalDate;
class RWOrganization;
class RWOrganizationRole;
class RWOrganizationalAddress;
class RWPerson;
class RWPersonAndOrganization;
class RWPersonAndOrganizationRole;
class RWPersonalAddress;
class RWPlaneAngleMeasureWithUnit;
class RWPlaneAngleUnit;
class RWProduct;
class RWProductCategory;
class RWProductContext;
class RWMechanicalContext; -- FMA le 24-07-96
-- Removed from Rev2 to Rev4 : class RWProductDataRepresentationView;
class RWProductDefinition;
class RWProductDefinitionContext;
class RWProductDefinitionFormation;
class RWProductDefinitionFormationWithSpecifiedSource;
class RWProductRelatedProductCategory;
class RWProductType;
class RWRatioMeasureWithUnit;
class RWSecurityClassification;
class RWSecurityClassificationLevel;
class RWSiUnit;
class RWSolidAngleMeasureWithUnit;
class RWSolidAngleUnit; -- Added by FMA
class RWUncertaintyMeasureWithUnit;
class RWWeekOfYearAndDayDate;

class RWSiUnitAndLengthUnit;
class RWSiUnitAndPlaneAngleUnit;
class RWSiUnitAndRatioUnit;      -- Added from Rev2 to Rev4
class RWSiUnitAndSolidAngleUnit; -- Added by FMA for Rev4
class RWSiUnitAndTimeUnit;       -- Added from Rev2 to Rev4
class RWSiUnitAndAreaUnit;
class RWSiUnitAndVolumeUnit;
class RWSiUnitAndMassUnit;  -- Added for AP209 (skl 15.12.2002)
class RWSiUnitAndThermodynamicTemperatureUnit;  -- Added for AP209 (skl 15.12.2002)
class RWConversionBasedUnitAndLengthUnit;
class RWConversionBasedUnitAndPlaneAngleUnit;
class RWConversionBasedUnitAndRatioUnit;      -- Added from Rev2 to Rev4
class RWConversionBasedUnitAndSolidAngleUnit; -- Added by FMA for Rev4
class RWConversionBasedUnitAndTimeUnit;       -- Added from Rev2 to Rev4
class RWConversionBasedUnitAndAreaUnit;
class RWConversionBasedUnitAndVolumeUnit;
class RWConversionBasedUnitAndMassUnit; -- added by skl 10.02.2004 for TRJ13
class RWMassMeasureWithUnit; -- added by skl 10.02.2004 for TRJ13

    -- Added from Rev2 to Rev4

class RWApprovalDateTime;
class RWDerivedUnit;
class RWDerivedUnitElement;

    -- Added from AP214 CC1 to CC2

class RWDocument;
--class RWDigitalDocument; same as for Document

class RWDocumentRelationship;
class RWDocumentType;
class RWDocumentUsageConstraint;
class RWEffectivity;
    class RWProductDefinitionEffectivity;
class RWProductDefinitionRelationship;

class RWProductDefinitionWithAssociatedDocuments;
--class RWPhysicallyModeledProductDefinition;  same as for ProductDefinition
   
 -- Added from AP214 CC2 to DIS
    
class RWCharacterizedObject;
class RWDocumentFile;

    -- Added for AP203
class RWAction;
class RWActionAssignment;
class RWActionMethod;
class RWActionRequestAssignment;
class RWVersionedActionRequest;
class RWCertification;
class RWCertificationAssignment;
class RWCertificationType;
class RWContract;
class RWContractAssignment;
class RWContractType;
class RWProductConceptContext;
class RWProductCategoryRelationship;
class RWActionRequestSolution;

-- added for external references (CAX-IF TRJ4)
class RWDocumentRepresentationType;
class RWExternalSource;
class RWExternallyDefinedItem;
class RWGeneralProperty;
class RWObjectRole;
class RWRoleAssociation;
class RWEffectivityAssignment;
class RWExternalIdentificationAssignment;
class RWIdentificationAssignment;
class RWIdentificationRole;
class RWNameAssignment;
class RWGroup;
class RWGroupAssignment;
class RWGroupRelationship;


---Added AP209
class RWEulerAngles;
class RWMassUnit;
class RWThermodynamicTemperatureUnit;
class RWProductDefinitionFormationRelationship;

-- added for external references (CAX-IF TRJ11 2003)
class RWDocumentProductAssociation;
class RWDocumentProductEquivalence;
	---Package Method ---

--	Init;
	---Purpose: enforced the initialisation of the  libraries

end RWStepBasic;
