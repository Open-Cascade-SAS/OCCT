-- Created on: 1995-08-09
-- Created by: Arnaud BOUZY/Odile Olivier
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

--   GG  :  GER61351 17/11/1999 Change SetColor() with a compatible Quantity_Color instead
--				       the restricted NameOfColor.

class Axis from AIS inherits InteractiveObject from AIS

	---Purpose: Locates the x, y and z axes in an Interactive Object.
    	-- These are used to orient it correctly in presentations
    	-- from different viewpoints, or to construct a revolved
    	-- shape, for example, from one of the axes. Conversely,
    	-- an axis can be created to build a revolved shape and
    	-- then situated relative to one of the axes of the view.

uses 
    Line                  from Geom,
    Presentation          from Prs3d,
    PresentationManager3d from PrsMgr,
    NameOfColor           from Quantity,
    Color			  from Quantity,
    Selection             from SelectMgr,
    Projector             from Prs3d,
    Transformation        from Geom,
    Pnt                   from gp,
    Dir                   from gp,    
    LineAspect            from Prs3d,
    TypeOfAxis            from AIS, 
    Axis2Placement        from Geom,
    Axis1Placement        from Geom,
    KindOfInteractive from AIS

is
    Create(aComponent : Line from Geom) 
    returns mutable Axis from AIS;
    	--- Purpose: Initializes the line aComponent   
    
    Create( aComponent : Axis2Placement from Geom;
    	    anAxisType: TypeOfAxis from AIS)
        ---Purpose: initializes the axis2 position
    	--   aComponent. The coordinate system used is right-handed.
    returns mutable Axis from AIS;

    Create(anAxis : Axis1Placement from Geom)
    returns mutable Axis from AIS;
    	---Purpose: Initializes the axis1 position anAxis.
    
    Component(me)
   	---Purpose:
	-- Returns the axis entity aComponent and identifies it
	-- as a component of a shape.
	---C++: inline
	---C++: return const &
    returns any Line from Geom 
    is static;

    SetComponent(me: mutable;aComponent : Line from Geom)
    is static;
    	---Purpose: Sets the coordinates of the lin aComponent.
    
    Axis2Placement(me)
    	---C++: inline
    	---C++: return const &  
    	---Purpose:
    	-- Returns the position of axis2 and   positions it by
    	-- identifying it as the x, y, or z axis and giving its
    	-- direction in 3D space. The coordinate system used is right-handed.    
    returns any Axis2Placement from Geom 
    is static;

    SetAxis2Placement(me: mutable;
    	    	      aComponent : Axis2Placement from Geom;
    	    	      anAxisType : TypeOfAxis from AIS)
    is static;
    	---Purpose:
    	-- Allows you to provide settings for aComponent:the
    	-- position and direction of an axis in 3D space. The
    	-- coordinate system used is right-handed. 
    
    SetAxis1Placement(me: mutable; anAxis     : Axis1Placement from Geom)
    is static;
    	---Purpose: Constructs a new line to serve as the axis anAxis in 3D space.
        
    TypeOfAxis (me)
     	---C++: inline
    	---Purpose: Returns the type of axis.
    returns TypeOfAxis from AIS;

    SetTypeOfAxis (me : mutable;aTypeAxis: TypeOfAxis from AIS)
       ---C++: inline
       ---Purpose:
       -- Constructs the entity aTypeAxis to stock information
       -- concerning type of axis.
    is static;

    IsXYZAxis  (me) 
       ---C++: inline
       ---Purpose:
       -- Returns a signature of 2 for axis datums. When you
       -- activate mode 2 by a signature, you pick AIS objects
       -- of type AIS_Axis.
    returns Boolean from Standard;

    AcceptDisplayMode(me;aMode:Integer from Standard) returns Boolean from  Standard is redefined static;
       ---Purpose: Returns true if the interactive object accepts the display mode aMode.
        
-- -- Methods from PresentableObject

    Compute(me            : mutable;
    	    aPresentationManager: PresentationManager3d from PrsMgr;
    	    aPresentation : mutable Presentation from Prs3d;
    	    aMode         : Integer from Standard = 0) 
    is redefined static  private;
    
    Compute(me:mutable;
    	        aProjector: Projector from Prs3d;
                aPresentation: mutable Presentation from Prs3d)
    is redefined static private;

    Compute(me            : mutable;
            aProjector    : Projector from Prs3d;
            aTrsf         : Transformation from Geom;
            aPresentation : mutable Presentation from Prs3d)
    is redefined;
	 ---Purpose: computes the presentation according to a point of view
	 --          given by <aProjector>.
	 --          To be Used when the associated degenerated Presentations
	 --          have been transformed by <aTrsf> which is not a Pure
	 --          Translation. The HLR Prs can't be deducted automatically
	 --          WARNING :<aTrsf> must be applied
	 --           to the object to display before computation  !!!

-- Methods from SelectableObject

    ComputeSelection(me         : mutable;
    	    	     aSelection : mutable Selection from SelectMgr;
    	    	     aMode      : Integer from Standard)is private;


-- -- Methods from InteractiveObject

    Signature(me) returns Integer from Standard is redefined;
    ---C++: inline

    Type(me) returns KindOfInteractive from AIS is redefined;
    ---C++: inline

    SetColor(me :mutable; aColor : NameOfColor from Quantity)
    is redefined static;
 
    SetColor(me :mutable; aColor : Color from Quantity) 
    is redefined static;
    
    SetWidth(me:mutable; aValue:Real from Standard) is redefined static;

    UnsetColor(me:mutable) is redefined static;
    
    UnsetWidth(me:mutable) is redefined static;


    ComputeFields(me: mutable)
    is private;

fields

    myComponent   : Line   from Geom;    
    myAx2         : Axis2Placement from Geom;
    myPfirst      : Pnt from gp;
    myPlast       : Pnt from gp;
    myTypeOfAxis  : TypeOfAxis from AIS;
    myIsXYZAxis   : Boolean from Standard;
    myDir         : Dir from gp;
    myVal         : Real from Standard;
    myText        : CString from Standard; 
    myLineAspect  : LineAspect from Prs3d;

end Axis;
