-- File:	STEPSelections_AssemblyComponent.cdl
-- Created:	Wed Mar 24 14:14:23 1999
-- Author:	data exchange team
--		<det@friendox.nnov.matra-dtv.fr>
---Copyright:	 Matra Datavision 1999


class AssemblyComponent from STEPSelections inherits TShared from MMgt

	---Purpose: 

uses
    
    ShapeDefinitionRepresentation from StepShape,
    HSequenceOfAssemblyLink from STEPSelections

is
    
    Create returns mutable AssemblyComponent from STEPSelections;
    
    Create (sdr : ShapeDefinitionRepresentation from StepShape;
    	    list: HSequenceOfAssemblyLink from STEPSelections)
    returns mutable AssemblyComponent from STEPSelections;
    
    --Methods for getting and obtaining fields
    
    GetSDR(me) returns ShapeDefinitionRepresentation from StepShape;
    	---Purpose:
	---C++: inline
    
    GetList(me) returns HSequenceOfAssemblyLink from STEPSelections;
    	---Purpose:
	---C++: inline
    
    SetSDR(me : mutable; sdr: ShapeDefinitionRepresentation from StepShape);
    	---Purpose:
	---C++: inline
    
    SetList(me : mutable; list: HSequenceOfAssemblyLink from STEPSelections);
    	---Purpose:
	---C++: inline

fields

    mySDR : ShapeDefinitionRepresentation from StepShape;
    myList: HSequenceOfAssemblyLink from STEPSelections;

end AssemblyComponent;
