-- Created on: 1993-12-06
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- jlr le 28-07-97 F(t) in Edge/Face



package BRepBlend

uses Blend, BlendFunc, AppBlend, Approx,  Adaptor3d,Adaptor2d,
     Law,  gp, TopAbs, IntSurf, Convert,
     TCollection,TColStd,TColgp,GeomAbs,Geom,Geom2d, 
     AdvApprox, StdFail, math

is

    class PointOnRst;
    class Extremity;
    class Line;

    class HCurveTool;
    class HCurve2dTool;

    class BlendTool;
    
    alias ConstRad is ConstRad from BlendFunc;

    alias ConstRadInv is ConstRadInv from BlendFunc;

    alias Ruled is Ruled from BlendFunc;

    alias RuledInv is RuledInv from BlendFunc;
    
    alias EvolRad is EvolRad from BlendFunc;

    alias EvolRadInv is EvolRadInv from BlendFunc;

    alias CSConstRad is CSConstRad from BlendFunc;

    alias CSCircular is CSCircular from BlendFunc;

    alias Chamfer is Chamfer from BlendFunc;

    alias ChamfInv is ChamfInv from BlendFunc;

    alias ChAsym is ChAsym from BlendFunc;

    alias ChAsymInv is ChAsymInv from BlendFunc;

    imported SequenceOfPointOnRst;

    class Walking instantiates Walking from Blend
    	(HVertex              from Adaptor3d,
	 HCurve2d             from Adaptor2d,
	 HSurface             from Adaptor3d,
	 HCurve               from Adaptor3d,
	 Integer              from Standard,
	 HCurve2dTool         from BRepBlend,
	 HSurfaceTool         from Adaptor3d,
	 HCurveTool           from BRepBlend,
	 TopolTool            from Adaptor3d,
	 BlendTool            from BRepBlend,
	 PointOnRst           from BRepBlend,
	 SequenceOfPointOnRst from BRepBlend,
	 Extremity            from BRepBlend,
	 Line                 from BRepBlend);
	 
    class CSWalking instantiates CSWalking from Blend
    	(HVertex              from Adaptor3d,
	 HCurve2d             from Adaptor2d,
	 HSurface             from Adaptor3d,
	 HCurve               from Adaptor3d,
	 Integer              from Standard,
	 HCurve2dTool         from BRepBlend,
	 HSurfaceTool         from Adaptor3d,
	 HCurveTool           from BRepBlend,
	 TopolTool            from Adaptor3d,
	 BlendTool            from BRepBlend,
	 PointOnRst           from BRepBlend,
	 SequenceOfPointOnRst from BRepBlend,
	 Extremity            from BRepBlend,
	 Line                 from BRepBlend);
	 
    class AppSurf instantiates AppSurf from AppBlend
    	(AppFunction from Blend,
         Line        from BRepBlend);


    imported SequenceOfLine;


    class AppSurface; 

    deferred class AppFuncRoot;

    class AppFunc;

    class AppFuncRst;

    class AppFuncRstRst;

    class SurfRstEvolRad;

    class SurfRstConstRad;

    class RstRstEvolRad;

    class RstRstConstRad;

    class SurfPointConstRadInv;

    class SurfCurvConstRadInv;

    class SurfPointEvolRadInv;

    class CurvPointRadInv;

    class SurfCurvEvolRadInv;

    class SurfRstLineBuilder;

    class RstRstLineBuilder;

end BRepBlend;
