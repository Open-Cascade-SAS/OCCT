-- Created on: 2000-10-24
-- Created by: Peter KURNEV
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class CompareRange from IntTools 

	---Purpose: Auxiliary class to provide a sorting Ranges, 
        --          taking  into  account a value of Left .   

uses
    Range from IntTools
--raises

is
    Create   
    	returns CompareRange from IntTools; 
	---Purpose:
	--- Empty constructor
	---
	 
    Create  (aTol:Real from Standard) 
    	returns CompareRange from IntTools;
	---Purpose:
	--- Initializes me by tolerance
	---
	 
    IsLower (me; Left, Right: Range from IntTools)
	---Purpose: 
    	--- Returns True if <Left> is lower than <Right>.
	---
    	returns Boolean from Standard;
    
    IsGreater (me; Left, Right: Range from IntTools)
	---Level: Public
	---Purpose: 
    	--- Returns True if <Left> is greater than <Right>.
	---
    	returns Boolean from Standard;

    IsEqual(me; Left, Right: Range from IntTools)
	---Level: Public
	---Purpose: 
    	--- Returns True when <Right> and <Left> are equal.
	---
    	returns Boolean from Standard ;

fields
    myTol: Real from Standard; 

end CompareRange;
