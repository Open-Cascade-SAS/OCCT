-- Created on: 1992-08-18
-- Created by: Remi Lequette
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package Hatch 

	---Purpose: The  Hatch package provides   algorithm to compute
	--          cross-hatchings on a 2D face.
	--          
	--          The  Hatcher algorithms stores a   set of lines in
	--          the 2D plane.
	--          
	--          The user stores lines in the Hatcher and afterward
	--          trim them with other lines.
	--          
	--          At any moment when  trimming the user can  ask for
	--          any  line  if   it is  intersected  and how   many
	--          intervals are defined on the line by the trim.

uses
    Standard,
    TCollection,
    gp

is
    enumeration LineForm is 
	---Purpose: Form of a trimmed line
	XLINE, YLINE, ANYLINE
    end LineForm;


    private class Parameter;

    imported SequenceOfParameter;

    private class Line;

    imported SequenceOfLine;
	    
    class Hatcher;

end Hatch;
