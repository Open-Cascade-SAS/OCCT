-- Created on: 1995-12-04
-- Created by: Laurent BOURESCHE
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class TgtOnCoons from GeomFill inherits TgtField from GeomFill

	---Purpose: Defines   an   algorithmic  tangents  field   on a
	--          boundary of a CoonsAlgPatch.

uses
    Vec           from gp,
    BSpline       from Law,
    CoonsAlgPatch from GeomFill

is
    Create(K : CoonsAlgPatch from GeomFill;
           I : Integer from Standard)
    returns mutable TgtOnCoons from GeomFill;

    Value(me; W : Real from Standard)
    returns Vec from gp;
    ---Purpose: Computes  the value  of the    field of tangency    at
    --          parameter W.

    D1(me; W : Real from Standard)
    returns Vec from gp;
    ---Purpose: Computes the  derivative of  the field of  tangency at
    --          parameter W.

    D1(me; W : Real from Standard; T, DT : out Vec from gp);
    ---Purpose: Computes the value and the  derivative of the field of
    --          tangency at parameter W.

fields

    myK    : CoonsAlgPatch from GeomFill;
    ibound : Integer from Standard;

end TgtOnCoons;
