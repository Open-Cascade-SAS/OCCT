-- Created on: 1992-06-04
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class CurveToolGeo from Geom2dGcc

uses Pnt2d        from gp,
     Vec2d        from gp,
     Lin2d        from gp,
     Circ2d       from gp,
     Elips2d      from gp,
     Parab2d      from gp,
     Hypr2d       from gp,
     CurveType    from GeomAbs,
     Shape        from GeomAbs,
     Curve        from Geom2dAdaptor,
     CurveTool    from Geom2dGcc,
     OffsetCurve  from Adaptor3d

is

    TheType(myclass; C: OffsetCurve from Adaptor3d ) 
    	returns CurveType from GeomAbs;

    Line(myclass; C: OffsetCurve from Adaptor3d)
    	---Purpose: Returns the Lin2d from gp corresponding to the curve C.
	--          This method is called only when TheType returns
	--          IntCurve_Lin.
    	returns Lin2d from gp;

    Circle(myclass; C: OffsetCurve from Adaptor3d)
    	---Purpose: Returns the Circ2d from gp corresponding to the curve C.
	--          This method is called only when TheType returns
	--          IntCurve_Cir.
    	returns Circ2d from gp;

    Ellipse(myclass; C: OffsetCurve from Adaptor3d)
	---Purpose: Returns the Elips2d from gp corresponding to the curve C.
	--          This method is called only when TheType returns
	--          IntCurve_Eli.
    	returns Elips2d from gp;

    Parabola(myclass; C: OffsetCurve from Adaptor3d)
	---Purpose: Returns the Parab2d from gp corresponding to the curve C.
	--          This method is called only when TheType returns
	--          IntCurve_Prb.
    	returns Parab2d from gp;

    Hyperbola(myclass; C: OffsetCurve from Adaptor3d)
	---Purpose: Returns the Hypr2d from gp corresponding to the curve C.
	--          This method is called only when TheType returns
	--          IntCurve_Hpr.
    	returns Hypr2d from gp;

-- The following method are used only when TheType returns  IntCurve_Other.

    FirstParameter(myclass;C: OffsetCurve from Adaptor3d)
    	returns Real;

    LastParameter(myclass;C: OffsetCurve from Adaptor3d)
    	returns Real;

    EpsX (myclass                     ; 
    	  C       : OffsetCurve from Adaptor3d    ;
    	  Tol     : Real from Standard)
    	returns Real;

    NbSamples(myclass                 ;
    	      C       : OffsetCurve from Adaptor3d)
    	returns Integer;

    Value (myclass                 ;
    	   C       : OffsetCurve from Adaptor3d;
    	   X       : Real          )
    	returns Pnt2d from gp;

    D1 (myclass; C :     OffsetCurve from Adaptor3d ;
    	    	 U :     Real           ;  
                 P : out Pnt2d          ;
    	    	 T : out Vec2d          );

    D2 (myclass; C   :     OffsetCurve from Adaptor3d ;
    	    	 U   :     Real           ; 
                 P   : out Pnt2d          ;
    	    	 T,N : out Vec2d          );

    IsComposite(myclass; C:OffsetCurve from Adaptor3d)
   
    	returns Boolean from Standard;

-- The following methods are used only when IsComposite returns True.

	
    GetIntervals(myclass ; C:OffsetCurve from Adaptor3d) returns Integer from Standard;
        ---Purpose : Outputs the number of interval of continuity C1 of 
        --           the curve
        --           used if Type == Composite.

    GetInterval (myclass; C      :     OffsetCurve from Adaptor3d
                       ; Index  :     Integer  from Standard
    	    	       ; U1, U2 : out Real     from Standard);
        ---Purpose : Outputs the bounds of interval of index <Index>
        --           used if Type == Composite.

    SetCurrentInterval (myclass; C: in out OffsetCurve from Adaptor3d
                              ; Index : Integer from Standard);
        ---Purpose : Set the current valid interval of index <Index>
        --           inside which the computations will be done
        --           (used if Type == Composite).

end CurveToolGeo;




