-- Created on: 1999-10-27
-- Created by: VKH
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Updated:     SZV IMP100701 Add the "depth" field and method
--              to the pixmap object.

class PixMap from WNT

    ---Version:

    ---Purpose: This class defines a windows bitmap

    ---Keywords: Bitmap, Pixmap

inherits
    PixMap                from Aspect

uses
    Handle                from Aspect,
    Color                 from Quantity,
    Window                from Aspect

raises
    PixmapDefinitionError from Aspect,
    PixmapError           from Aspect

is

    Create ( aWindow          : Window from Aspect;
             aWidth, anHeight : Integer from Standard;
             aCDepth          : Integer from Standard = 0 )
    returns mutable PixMap from WNT
    raises PixmapDefinitionError from Aspect;
    ---Level: Public
    ---Purpose:  Warning! When <aDepth> is NULL , the pixmap is created
    -- with the SAME depth than the window <aWindow>

    ---------------------------------------------------
    -- Category: Methods to modify the class definition
    ---------------------------------------------------

    Destroy ( me : mutable )
    ---Level: Advanced
    ---Purpose: Destroies the Bitmap
    ---C++: alias ~
    --  Trigger: Raises if Bitmap is not defined properly
    raises PixmapError from Aspect is virtual;

    Dump ( me; aFilename : CString from Standard ;
           aGammaValue: Real from Standard = 1.0 )
    returns Boolean
    ---Level: Advanced
    ---Purpose:
    -- Dumps the Bitmap to an image file with
    -- an optional gamma correction value
    -- and returns TRUE if the dump occurs normaly.
    ---Category: Methods to modify the class definition
    raises PixmapError from Aspect is virtual;

    PixelColor ( me         : in;
                 theX, theY : in Integer from Standard )
    returns Color from Quantity
    is virtual;
    ---Purpose:
    -- Returns the pixel color.

    ----------------------------
    -- Category: Inquire methods
    ----------------------------

    PixmapID ( me ) returns Handle from Aspect is virtual;
    ---Level: Advanced
    ---Purpose: Returns the ID of the just created bitmap
    ---Category: Inquire methods

    ----------------------------
    -- Category: Private methods
    ----------------------------

    PreferedDepth( me ; aWindow: Window from Aspect;
                   aDepth: Integer from Standard)
    returns Integer from Standard is private;

fields
    myDC       : Handle from Aspect is protected;
    myBitmap   : Handle from Aspect is protected;
    myWND      : Window from Aspect;
end PixMap;
