-- Created on: 1993-04-06
-- Created by: Philippe DAUTRY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class Conic from PGeom2d inherits Curve from PGeom2d

        ---Purpose : Defines the general   characteristics of a  conic
        --         curve : Ellipse, Circle, Hyperbola, Parabola.
        --  
	---See Also : Conic from Geom2d

uses  Ax22d from gp

is


    Initialize;
	---Purpose: Initializes the field(s) with default value(s).
	---Level: Internal 


    Initialize(aPosition: Ax22d from gp);
	---Purpose: Initializes the field position with <aPosition>.
	---Level: Internal 


  Position (me : mutable; aPosition : Ax22d from gp);
        ---Purpose : Set the value of the field position with <aPosition>.
	---Level: Internal 


  Position (me)   returns Ax22d from gp;
        ---Purpose : Returns the value of the field <position>.
	---Level: Internal 


fields

  position : Ax22d from gp is protected;

end;
