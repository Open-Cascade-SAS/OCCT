-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class EdgeCurve from StepShape 

inherits Edge from StepShape 
-- WARNING : Multiple EXPRESS inheritance
-- Not yet automaticly managed
-- inherits GeometricRepresentationItem from StepShape 

uses

	Curve from StepGeom, 
	Boolean from Standard, 
	HAsciiString from TCollection, 
	Vertex from StepShape
is

	Create returns mutable EdgeCurve;
	---Purpose: Returns a EdgeCurve


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aEdgeStart : mutable Vertex from StepShape;
	      aEdgeEnd : mutable Vertex from StepShape) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aEdgeStart : mutable Vertex from StepShape;
	      aEdgeEnd : mutable Vertex from StepShape;
	      aEdgeGeometry : mutable Curve from StepGeom;
	      aSameSense : Boolean from Standard) is virtual;

	-- Specific Methods for Field Data Access --

	SetEdgeGeometry(me : mutable; aEdgeGeometry : mutable Curve);
	EdgeGeometry (me) returns mutable Curve;
	SetSameSense(me : mutable; aSameSense : Boolean);
	SameSense (me) returns Boolean;

fields

	edgeGeometry : Curve from StepGeom;
	sameSense : Boolean from Standard;

end EdgeCurve;
