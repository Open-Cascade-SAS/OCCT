-- Created on: 1991-10-02
-- Created by: NW,JPB,CAL
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Background from Aspect


	---Purpose: This class allows the definition of
	--	    a window background.

uses

	Color	from Quantity

is

	Create
		returns Background from Aspect;
	---Level: Public
	---Purpose: Creates a window background.
	--	    Default color : NOC_MATRAGRAY.

	Create ( AColor : Color from Quantity )
		returns Background from Aspect;
	---Level: Public
	---Purpose: Creates a window background with the colour <AColor>.

	---------------------------------------------------
	-- Category: Methods to modify the class definition
	---------------------------------------------------

	SetColor ( me		: in out;
		   AColor	: Color from Quantity );
	---Level: Public
	---Purpose: Modifies the colour of the window background <me>.
	---Category: Methods to modify the class definition

	----------------------------
	-- Category: Inquire methods
	----------------------------

	Color ( me )
		returns Color from Quantity;
	---Level: Public
	---Purpose: Returns the colour of the window background <me>.
	---Category: Inquire methods

--

fields

--
-- Class	:	Aspect_Background
--
-- Purpose	:	Declaration of variables specific to the window
--			background.
--
-- Reminder	:	A background is defined by one colour
--

	-- the colour associated with the window background
	MyColor	:	Color from Quantity;

end Background;
