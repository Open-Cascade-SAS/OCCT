-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DateAndTime from StepBasic 

inherits TShared from MMgt

uses

	Date from StepBasic, 
	LocalTime from StepBasic
is

	Create returns mutable DateAndTime;
	---Purpose: Returns a DateAndTime

	Init (me : mutable;
	      aDateComponent : mutable Date from StepBasic;
	      aTimeComponent : mutable LocalTime from StepBasic) is virtual;

	-- Specific Methods for Field Data Access --

	SetDateComponent(me : mutable; aDateComponent : mutable Date);
	DateComponent (me) returns mutable Date;
	SetTimeComponent(me : mutable; aTimeComponent : mutable LocalTime);
	TimeComponent (me) returns mutable LocalTime;

fields

	dateComponent : Date from StepBasic;
	timeComponent : LocalTime from StepBasic;

end DateAndTime;
