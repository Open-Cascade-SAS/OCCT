-- File:        PcurveOrSurface.cdl
-- Created:     Fri Dec  1 11:11:11 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993



class PcurveOrSurface from StepGeom inherits SelectType from StepData

	-- <PcurveOrSurface> is an EXPRESS Select Type construct translation.
	-- it gathers : Pcurve, Surface

uses

	Pcurve,
	Surface
is

	Create returns PcurveOrSurface;
	---Purpose : Returns a PcurveOrSurface SelectType

	CaseNum (me; ent : Transient) returns Integer;
	---Purpose: Recognizes a PcurveOrSurface Kind Entity that is :
	--        1 -> Pcurve
	--        2 -> Surface
	--        0 else

	Pcurve (me) returns any Pcurve;
	---Purpose : returns Value as a Pcurve (Null if another type)

	Surface (me) returns any Surface;
	---Purpose : returns Value as a Surface (Null if another type)


end PcurveOrSurface;

