-- Created on: 1993-04-06
-- Created by: Philippe DAUTRY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class VectorWithMagnitude from PGeom2d inherits Vector from PGeom2d

        ---Purpose : Defines a vector  with  magnitude.  A vector with
        --         magnitude can have a zero length.
        --         
	---See Also : VectorWithMagnitude from Geom2d.

uses Vec2d from gp

is


  Create returns mutable VectorWithMagnitude;
        ---Purpose : Creates a VectorWithMagnitude with default values.
	---Level: Advanced 


  Create (aVec : Vec2d from gp) returns mutable VectorWithMagnitude;
        ---Purpose : Creates a VectorWithMagnitude with <aVec>.
	---Level: Advanced 


end;
