-- Created on: 1994-03-30
-- Created by: Laurent BUCHARD
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

generic class Classifier3d from TopClass 
    	(TheIntersector as any)  -- as Intersection3d from TopClass

	---Purpose: 

uses
    Lin             from gp,
    CurveTransition from TopTrans,
    Orientation     from TopAbs,
    State           from TopAbs,
    Face            from TopoDS

raises
    DomainError from Standard
    
is
    Create returns Classifier3d from TopClass;
	---Purpose: Creates an undefined classifier.
	
    Reset(me : in out; L   : Lin  from gp;
                       P   : Real from Standard; 
                       Tol : Real from Standard)
	---Purpose: Starts  a  classification process.   The  point to
	--          classify is the origin of  the  line <L>.  <P>  is
	--          the original length of the segment on <L>  used to
	--          compute  intersections.   <Tol> is the   tolerance
	--          attached to the intersections.
    is static;
    
    Compare(me : in out; F   : Face        from TopoDS;
                         Or  : Orientation from TopAbs)
	---Purpose: Updates  the classification process with  the face
	--          <F> from the boundary. 
    raises
    	DomainError  -- The classifier has not been set
    is static;

    Parameter(me) returns Real
	---Purpose: Returns the current value of the parameter.
	---C++: inline
    is static;

    HasIntersection(me) returns Boolean from Standard
    	---Purpose: Returns True if an intersection is computed.
    is static;

    Intersector(me : in out) returns TheIntersector
	---Purpose: Returns the intersecting algorithm.
	--          
	---C++: inline
	---C++: return &
    is static;
    
    State(me) returns State from TopAbs
	---Purpose: Returns the current state of the point.
	--          
	---C++: inline
    is static;
    

fields
    isSet          : Boolean          from Standard;
    myFace         : Face             from TopoDS;
    myLin          : Lin              from gp;
    myParam        : Real             from Standard;
    myTolerance    : Real             from Standard;
    myState        : State            from TopAbs;
    hasIntersect   : Boolean          from Standard;
    myIntersector  : TheIntersector;
    
end Classifier3d;

