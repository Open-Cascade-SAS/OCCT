-- Created on: 1997-02-10
-- Created by: Alexander BRIVIN
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Info from Vrml 

	---Purpose:  defines a Info node of VRML specifying properties of geometry
	---          and its appearance. 
    	--  It  is  used  to  store  information  in  the  scene  graph, 
	--  Typically  for  application-specific  purposes,  copyright  messages, 
	--  or  other  strings.
uses

     AsciiString from TCollection
is
 
    Create  (  aString  :  AsciiString from TCollection  =  "<Undefined info>")    
        returns Info from Vrml; 

    SetString ( me : in out;  aString  :  AsciiString from TCollection ); 
    String ( me  )  returns  AsciiString from TCollection; 
   
    Print  ( me;  anOStream: in out OStream from Standard ) returns OStream from Standard;
    ---C++:  return  & 

fields
 
    myString  :  AsciiString from TCollection;  -- Info string

end Info;

