-- Created on: 1993-06-17
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class WireEdgeClassifier from TopOpeBRepBuild
    inherits CompositeClassifier from TopOpeBRepBuild
    
---Purpose: 
-- Classify edges and wires.
-- shapes are Wires, Element are Edge.

uses
    
    ShapeEnum from TopAbs,
    State from TopAbs,
    Shape from TopoDS,
    Pnt2d from gp,
    Edge from BRepClass,
    FacePassiveClassifier from BRepClass,
    BlockBuilder from TopOpeBRepBuild,
    Loop from TopOpeBRepBuild
    
is

    Create(F : Shape from TopoDS;
    	   BB : BlockBuilder) returns WireEdgeClassifier;
    ---Purpose: Creates a classifier on edge <F>.  
    -- Used to compare edges and wires on the edge <F>.

    Compare(me : in out; L1,L2 : Loop) returns State from TopAbs
    is redefined;

    LoopToShape(me : in out; L : Loop)
    returns Shape from TopoDS;

    CompareShapes(me : in out; B1,B2 : Shape from TopoDS)
    ---Purpose: classify wire <B1> with wire <B2>
    returns State from TopAbs;
    
    CompareElementToShape(me : in out; E,B : Shape from TopoDS)
    ---Purpose: classify edge <E> with wire <B>
    returns State from TopAbs;
    
    ResetShape(me : in out; B : Shape from TopoDS);
    ---Purpose: prepare classification involving wire <B>
    -- calls ResetElement on first edge of <B>
    
    ResetElement(me : in out; E : Shape from TopoDS);
    ---Purpose: prepare classification involving edge <E>
    -- define 2D point (later used in Compare()) on first vertex of edge <E>.
    
    CompareElement(me : in out; E : Shape from TopoDS);
    ---Purpose: Add the edge <E> in the set of edges used in 2D point
    -- classification.
    
    State(me : in out) returns State from TopAbs;
    ---Purpose: Returns state of classification of 2D point, defined by 
    -- ResetElement, with the current set of edges, defined by Compare.

fields
    
    myFirstCompare : Boolean;
    myPoint2d : Pnt2d from gp;
    myBCEdge : Edge from BRepClass;
    myFPC : FacePassiveClassifier from BRepClass; 
    myShape : Shape from TopoDS;
    
end WireEdgeClassifier from TopOpeBRepBuild;
