-- Created on: 1995-10-26
-- Created by: Yves FRICAUD
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class AsDes from BRepAlgo inherits TShared from MMgt

	---Purpose: SD to store descendants and ascendants of Shapes.

uses
    DataMapOfShapeListOfShape from TopTools,
    ListOfShape               from TopTools,
    Shape                     from TopoDS

raises
    ConstructionError from Standard 

is
    Create returns AsDes from BRepAlgo;
	---Purpose: Creates an empty AsDes.
    
    Clear(me : mutable);
    
    Add  (me : mutable ; S  : Shape from TopoDS;
    	    	         SS : Shape from TopoDS)
       ---Purpose: Stores <SS> as a futur subshape of <S>. 
    is static;		       

    Add (me : mutable ; S  : Shape from TopoDS;
    	    	        SS : ListOfShape from TopTools)
       ---Purpose: Stores <SS> as futurs SubShapes of <S>. 		       
    is static;		       

    HasAscendant(me; S : Shape from TopoDS)
    returns Boolean from Standard;

    HasDescendant(me; S : Shape from TopoDS)
    returns Boolean from Standard;
		       
    Ascendant (me; S : Shape from TopoDS)
    	---Purpose: Returns the Shape containing <S>. 
    	---C++: return const &
    returns ListOfShape from TopTools;

    Descendant (me; S : Shape from TopoDS)
	---Purpose: Returns futur subhapes of <S>.
    	---C++: return const &
    returns ListOfShape from TopTools;
    
    ChangeDescendant (me : mutable; S : Shape from TopoDS)
	---Purpose: Returns futur subhapes of <S>.
    	---C++: return &
    returns ListOfShape from TopTools;
    
    Replace ( me : mutable; OldS, NewS : Shape from TopoDS)
    	---Purpose: Replace <OldS> by <NewS>.
    	--          <OldS> disapear from <me>.
    is static;
        
    Remove  (me  :  mutable; 
    	     S   :  Shape  from  TopoDS) 
    	---Purpose: Remove <S> from me.
    raises 
	ConstructionError -- if <S> HasDescendant.    
    is static; 
     
    HasCommonDescendant  (me ;   
    	    	    	  S1 :           Shape        from  TopoDS;   
			  S2 :           Shape        from  TopoDS;  
    	    	    	  LC :  in  out  ListOfShape  from  TopTools)  
	 ---Purpose: Returns  True if (S1> and <S2>  has  common 
	 --           Descendants.  Stores in <LC> the Commons Descendants.
    returns  Boolean  from  Standard; 
     
    BackReplace ( me : mutable; 
    	    	  OldS : Shape       from TopoDS;
    	    	  NewS : Shape       from TopoDS;
    	    	  L    : ListOfShape from TopTools;
		  InUp : Boolean     from Standard)  
    	---Purpose: Replace <OldS> by <NewS>.
    	--          <OldS> disapear from <me>.
    is static private; 
     
	     
fields

    up   : DataMapOfShapeListOfShape from TopTools;
    down : DataMapOfShapeListOfShape from TopTools;

end AsDes;
