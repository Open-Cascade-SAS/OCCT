-- File:	IGESGraph_ToolNominalSize.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolNominalSize  from IGESGraph

    ---Purpose : Tool to work on a NominalSize. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses NominalSize from IGESGraph,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolNominalSize;
    ---Purpose : Returns a ToolNominalSize, ready to work


    ReadOwnParams (me; ent : mutable NominalSize;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : NominalSize;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : NominalSize;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a NominalSize <ent>, from
    --           its specific (own) parameters

    OwnCorrect (me; ent : mutable NominalSize) returns Boolean  is static;
    ---Purpose : Sets automatic unambiguous Correction on a NominalSize
    --           (NbPropertyValues forced to 2 or 3 according HasStandardName)

    DirChecker (me; ent : NominalSize) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : NominalSize;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : NominalSize; entto : mutable NominalSize;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : NominalSize;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolNominalSize;
