-- Created by: DAUTRY Philippe
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

--      	---------------------

---Version:	0.0
--Version	Date		Purpose
--		0.0	Jul  6 1998	Creation
--		1.0	Jul  6 1998	Separation Forget/Resume

class DeltaOnResume from TDF inherits AttributeDelta from TDF

	---Purpose: This class provides default services for an
	--          AttributeDelta on an Resume action.
	--          
	--          Applying this AttributeDelta means FORGETTING its
	--          attribute.

uses

    Attribute from TDF

is

    Create(anAtt : Attribute from TDF)
    	returns mutable DeltaOnResume from TDF;
	---Purpose: Creates a TDF_DeltaOnResume.

    Apply (me : mutable)
    	is redefined static;
    	---Purpose: Applies the delta to the attribute.

end DeltaOnResume;
