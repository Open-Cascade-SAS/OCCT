-- Created on: 1995-01-25
-- Created by: Jean-Louis Frenkel
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package PrsMgr
    	---Purpose: The PrsMgr package provides low level services
    	-- and is only to be used when you do not want to use
    	-- the services provided by AIS.
    	-- PrsMgr manages display through the following services:
    	-- -   supplying a graphic structure for the object to be presented
    	-- -   recalculating presentations when required, e.g. by
    	--   moving the object or changing its color
    	-- -   defining the display mode of the object to be
    	--   presented; in the case of AIS_Shape, for example,
    	--   this determines whether the object is to be displayed in:
    	--   -   wireframe 0
    	--   -   shading 1.
    	-- Note that each new Interactive Object must have all its display modes defined.
        
uses

    MMgt,TCollection,
    TopLoc,
    Aspect,
    Prs3d,
    Graphic3d,
    Quantity,Geom,
    Visual3d,
    V3d,
    TColStd, 
    gp
 
is

    enumeration TypeOfPresentation3d is TOP_AllView, TOP_ProjectorDependant
    end TypeOfPresentation3d;
    	---Purpose: To declare the type of presentation as follows
    	-- -   AllView for display involving no recalculation for
    	--   new projectors (points of view)in hidden line removal mode
    	-- -   ProjectorDependant for display in hidden line
    	--   removal mode, where every new point of view
    	--   entails recalculation of the display.

    class PresentationManager;
    alias PresentationManager3d is PresentationManager;
    class Presentation;
    alias Presentation3d is Presentation;
    deferred class PresentableObject;

    imported ListOfPresentations;
    imported ListOfPresentableObjects;

    class Prs;

    class ModedPresentation;
    class Presentations  instantiates Sequence from TCollection
    	(ModedPresentation from PrsMgr);
    pointer PresentationPointer to Presentation from PrsMgr;
    pointer PresentableObjectPointer to PresentableObject from PrsMgr;
end PrsMgr;
