-- Created on: 2003-10-13
-- Created by: Alexander SOLOVYOV
-- Copyright (c) 2003-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class TextPrsBuilder from MeshVS inherits PrsBuilder from MeshVS

	---Purpose: This class provides methods to create text data presentation.
        -- It store map of texts assigned with nodes or elements.

uses
  Real from Standard,

  Presentation from Prs3d,

  Boolean from Standard,
  Integer from Standard,

  Mesh                        from MeshVS,
  MeshPtr                     from MeshVS,
  DisplayModeFlags            from MeshVS,
  DataSource                  from MeshVS,
  DataMapOfIntegerAsciiString from MeshVS,
  BuilderPriority             from MeshVS,
  Color                       from Quantity,
  AsciiString                 from TCollection,
  PackedMapOfInteger          from TColStd

is

  Create  ( Parent   : Mesh from MeshVS;
            Height   : Real;
            Color    : Color from Quantity;
            Flags    : DisplayModeFlags from MeshVS = MeshVS_DMF_TextDataPrs;
            DS       : DataSource from MeshVS = 0;
            Id       : Integer = -1;
            Priority : BuilderPriority from MeshVS = MeshVS_BP_Text ) returns mutable TextPrsBuilder from MeshVS;

  Build   ( me; Prs        : Presentation from Prs3d;
            IDs            : PackedMapOfInteger;
            IDsToExclude   : in out PackedMapOfInteger;
            IsElement      : Boolean;
            theDisplayMode : Integer ) is virtual;
	---Purpose: Builds presentation of text data

  GetTexts ( me; IsElement : Boolean ) returns DataMapOfIntegerAsciiString from MeshVS;
	---C++: return const &
	---Purpose: Returns map of text assigned with nodes ( IsElement = False ) or elements ( IsElement = True )

  SetTexts ( me : mutable;
             IsElement     : Boolean;
             Map           : DataMapOfIntegerAsciiString from MeshVS );
	---Purpose: Sets map of text assigned with nodes or elements

  HasTexts ( me; IsElement : Boolean )    returns Boolean;
	---Purpose: Returns True if map isn't empty

  GetText  ( me; IsElement : Boolean;
             ID            : Integer;
             Text          : out AsciiString from TCollection )   returns Boolean;
	---Purpose: Returns text assigned with single node or element

  SetText  ( me : mutable;
             IsElement     : Boolean;
             ID            : Integer;
             Text          : AsciiString from TCollection );
	---Purpose: Sets text assigned with single node or element

fields
  myNodeTextMap         : DataMapOfIntegerAsciiString from MeshVS;
  myElemTextMap         : DataMapOfIntegerAsciiString from MeshVS;

end TextPrsBuilder;
