-- File:	STEPSelections_AssemblyLink.cdl
-- Created:	Wed Mar 24 12:40:23 1999
-- Author:	data exchange team
--		<det@friendox.nnov.matra-dtv.fr>
---Copyright:	 Matra Datavision 1999


class AssemblyLink from STEPSelections inherits TShared from MMgt

	---Purpose: 

uses
    
    NextAssemblyUsageOccurrence from StepRepr,
    ContextDependentShapeRepresentation from StepShape,
    AssemblyComponent from STEPSelections

is

    Create returns mutable AssemblyLink from STEPSelections;
    
    Create(nauo: NextAssemblyUsageOccurrence from StepRepr;
    	   item: Transient from Standard;
	   part: AssemblyComponent from STEPSelections)
    returns mutable AssemblyLink from STEPSelections;
    
    --Methods for setting and obtaining fields
    
    GetNAUO(me) returns NextAssemblyUsageOccurrence from StepRepr;
    	---Purpose:
	---C++: inline
	
    GetItem(me) returns Transient from Standard;
    	---Purpose:
	---C++: inline
	
    GetComponent(me) returns AssemblyComponent from STEPSelections;
    	---Purpose:
	---C++: inline
    
    SetNAUO(me: mutable; nauo: NextAssemblyUsageOccurrence from StepRepr);
    	---Purpose:
	---C++: inline
	
    SetItem(me: mutable; item: Transient from Standard);
    	---Purpose:
	---C++: inline
    
    SetComponent(me: mutable; part: AssemblyComponent from STEPSelections);
	---Purpose:
	---C++: inline

fields

    myNAUO     : NextAssemblyUsageOccurrence from StepRepr;
    myItem     : Transient from Standard;
    myComponent: AssemblyComponent from STEPSelections;

end AssemblyLink;
