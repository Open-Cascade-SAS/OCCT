-- Created on: 1994-06-24
-- Created by: Yves FRICAUD
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Inter from Bisector 

	---Purpose: Intersection between two <Bisec> from Bisector.

inherits 
    Intersection from IntRes2d
    
uses   
    Domain  from IntRes2d,
    Bisec   from Bisector,
    Curve   from Bisector,
    BisecCC from Bisector,
    Curve   from Geom2d,
    Line    from Geom2d
    
raises ConstructionError from Standard

is
    Create returns Inter from Bisector;
    
    Create (C1: Bisec from Bisector; D1: Domain from IntRes2d;
            C2: Bisec from Bisector; D2: Domain from IntRes2d;
    	    TolConf,Tol  : Real    from Standard;
    	    ComunElement : Boolean from Standard) 
	---Purpose: Intersection between 2 curves.  
	--          C1 separates the element A and B. 
	--          C2 separates the elements C et D.
	--          If B an C have the same geometry. <ComunElement>
	--          Has to be True. 
	--          It Permits an optimiztion of the computation.

    returns  Inter from Bisector
    raises   ConstructionError from Standard;

    
    Perform (me: in out;
             C1: Bisec from Bisector; D1: Domain from IntRes2d;
             C2: Bisec from Bisector; D2: Domain from IntRes2d;
    	     TolConf,Tol  : Real    from Standard;
    	     ComunElement : Boolean from Standard) 
	---Purpose: Intersection between 2 curves.          
    	--          C1 separates the element A and B. 
	--          C2 separates the elements C et D.
	--          If B an C have the same geometry. <ComunElement>
	--          Has to be True. 
	--          It Permits an optimiztion of the computation.

    raises   ConstructionError from Standard
    is static;
    
    SinglePerform (me: in out;
             	   C1: Curve from Geom2d ; D1: Domain from IntRes2d;
             	   C2: Curve from Geom2d ; D2: Domain from IntRes2d;
    	           TolConf,Tol  : Real    from Standard;
    	           ComunElement : Boolean from Standard) 
	---Purpose: Intersection between 2 curves.          
    
    raises   ConstructionError from Standard
    is static private;
	
    NeighbourPerform (me : in out;
    	    	      C1 : BisecCC from Bisector; D1: Domain from IntRes2d;
                      C2 : BisecCC from Bisector; D2: Domain from IntRes2d;
    	              Tol: Real    from Standard)
    is static private;
    
    TestBound (me : in out;
    	       C1 : Line  from Geom2d  ; D1      : Domain  from IntRes2d;
    	       C2 : Curve from Geom2d  ; D2      : Domain  from IntRes2d;
	       Tol: Real  from Standard; Reverse : Boolean from Standard)
    is static private;
    
end Inter;
