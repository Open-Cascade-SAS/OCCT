-- File:	IGESGraph_ToolDrawingUnits.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolDrawingUnits  from IGESGraph

    ---Purpose : Tool to work on a DrawingUnits. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses DrawingUnits from IGESGraph,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolDrawingUnits;
    ---Purpose : Returns a ToolDrawingUnits, ready to work


    ReadOwnParams (me; ent : mutable DrawingUnits;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : DrawingUnits;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : DrawingUnits;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a DrawingUnits <ent>, from
    --           its specific (own) parameters

    OwnCorrect (me; ent : mutable DrawingUnits) returns Boolean  is static;
    ---Purpose : Sets automatic unambiguous Correction on a DrawingUnits
    --           (NbPropertyValues forced to 2)

    DirChecker (me; ent : DrawingUnits) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : DrawingUnits;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : DrawingUnits; entto : mutable DrawingUnits;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : DrawingUnits;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolDrawingUnits;
