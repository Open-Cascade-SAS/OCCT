-- Created by: PLOTNIKOV Eugeny
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Image from WNT inherits TShared from MMgt

	---Purpose: Internal class for image management

 uses

    Handle from Aspect

 is

    Create ( aBitmap : Handle from Aspect; aHashCode : Integer from Standard )
     returns mutable Image from WNT;
    	---Purpose: Creates a class.

    Destroy ( me : mutable ) is virtual;
	---Level:   Public
	---Purpose: Destroys all ressources attached to the Image
    ---C++:     alias ~

    HBITMAP ( me ) returns Handle from Aspect;
    ---Level:   Public
    ---Purpose: Returns bitmap handle
    ---C++:     inline

    Image ( me ) returns Address from Standard;
    ---Level:   Public
    ---Purpose: Returns pointer to internal structure
    ---C++:     inline

 fields

    myImage    : Address from Standard is protected;
    myHashCode : Integer from Standard is protected;

end Image;
