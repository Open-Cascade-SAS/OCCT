-- Created on: 1992-11-17
-- Created by: Christian CAILLET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DispPerOne  from IFSelect  inherits Dispatch

    ---Purpose : A DispPerOne gathers all the input Entities into as many
    --           Packets as there Root Entities from the Final Selection,
    --           that is, one Packet per Entity

uses AsciiString from TCollection, Graph, SubPartsIterator

is

    Create returns mutable DispPerOne;
    ---Purpose : Creates a DispPerOne

    Label (me) returns AsciiString from TCollection;
    ---Purpose : Returns as Label, "One File per Input Entity"

    	--  --    Evaluation    --  --

    LimitedMax (me; nbent : Integer; max : out Integer) returns Boolean
    	is redefined;
    ---Purpose : Returns True, maximum limit is given as <nbent>

    PacketsCount (me; G : Graph; count : out Integer) returns Boolean
    	is redefined;
    ---Purpose : Returns True (count is easy to know) and count is the length
    --           of the input list (RootResult from FinalSelection)

    Packets (me; G : Graph; packs : in out SubPartsIterator);
    ---Purpose : Returns the list of produced Packets. It defines one Packet
    --           per Entity given by RootResult from the Final Selection.

end DispPerOne;
