-- File:        BSplineSurfaceWithKnotsAndRationalBSplineSurface.cdl
-- Created:     Mon Dec  4 12:02:34 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWBSplineSurfaceWithKnotsAndRationalBSplineSurface from RWStepGeom

	---Purpose : Read & Write Module for BSplineSurfaceWithKnotsAndRationalBSplineSurface
	--           Check added by CKY , 7-OCT-1996

uses Check from Interface, ShareTool from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     BSplineSurfaceWithKnotsAndRationalBSplineSurface from StepGeom,
     EntityIterator from Interface

is

	Create returns RWBSplineSurfaceWithKnotsAndRationalBSplineSurface;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable BSplineSurfaceWithKnotsAndRationalBSplineSurface from StepGeom);

	WriteStep (me; SW : in out StepWriter; ent : BSplineSurfaceWithKnotsAndRationalBSplineSurface from StepGeom);

	Share(me; ent : BSplineSurfaceWithKnotsAndRationalBSplineSurface from StepGeom; iter : in out EntityIterator);

    	Check(me; ent : BSplineSurfaceWithKnotsAndRationalBSplineSurface from StepGeom; shares : ShareTool; ach : in out Check);

end RWBSplineSurfaceWithKnotsAndRationalBSplineSurface;
