-- Created on: 1996-04-10
-- Created by: Joelle CHAUVET
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Modified:	Wed Jan 15 09:45:42 1997
--    by:	Joelle CHAUVET
--		G1135 : Methods CutSense with criterion, Coefficients,
--		                CritValue, SetCritValue,
--		        Field 'myCritValue'

class Patch from AdvApp2Var

uses

    Boolean,Integer,Real from Standard,
    HArray1OfReal,HArray2OfReal from TColStd,
    HArray2OfPnt from TColgp,
    EvaluatorFunc2Var,Context,Framework,Criterion from AdvApp2Var

is

    Create returns Patch;
    Create(U0,U1,V0,V1 : Real; iu,iv : Integer) returns Patch;
    Create(P : Patch) returns Patch is private;
    IsDiscretised(me) returns Boolean;
    Discretise(me: in out; Conditions : Context;
    	    	    	   Constraints: Framework;
    	    	    	   func : EvaluatorFunc2Var);
    IsApproximated(me) returns Boolean;
    HasResult(me) returns Boolean;
    MakeApprox(me: in out; Conditions : Context;
    	    	    	   Constraints: Framework;
    	    	    	   NumDec : Integer);
    AddConstraints(me: in out; Conditions : Context;
    	    	    	       Constraints: Framework);
    AddErrors(me: in out; Constraints: Framework);
    ChangeDomain(me: in out; a,b,c,d : Real);
    ResetApprox(me: in out);
    OverwriteApprox(me: in out);
    U0(me) returns Real;
    U1(me) returns Real;
    V0(me) returns Real;
    V1(me) returns Real;
    UOrder(me) returns Integer;
    VOrder(me) returns Integer;
    CutSense(me) returns Integer;
    CutSense(me; Crit : Criterion; NumDec : Integer) returns Integer;
    NbCoeffInU(me) returns Integer;
    NbCoeffInV(me) returns Integer;
    ChangeNbCoeff(me: in out; NbCoeffU, NbCoeffV : Integer);
    Poles(me; SSPIndex : Integer; Conditions : Context) returns HArray2OfPnt;
    Coefficients(me; SSPIndex : Integer; Conditions : Context) returns HArray1OfReal;
    MaxErrors(me) returns HArray1OfReal;
    AverageErrors(me) returns HArray1OfReal;
    IsoErrors(me) returns HArray2OfReal;
    CritValue(me) returns Real;
    SetCritValue(me: in out; dist : Real);

fields

    myU0, myU1    : Real;
    myV0, myV1    : Real;
    myOrdInU      : Integer;
    myOrdInV      : Integer;
    myNbCoeffInU  : Integer;
    myNbCoeffInV  : Integer;
    myApprIsDone  : Boolean;
    myHasResult   : Boolean;
    myEquation    : HArray1OfReal;
    myMaxErrors   : HArray1OfReal;
    myMoyErrors   : HArray1OfReal;
    myIsoErrors   : HArray2OfReal;
    myCutSense    : Integer;
    myDiscIsDone  : Boolean;
    mySosoTab     : HArray1OfReal;
    myDisoTab     : HArray1OfReal;
    mySodiTab     : HArray1OfReal;
    myDidiTab     : HArray1OfReal;
    myCritValue   : Real;

end Patch;
















