-- File:	MeshAlgo_Vertex.cdl
-- Created:	Tue May 11 16:17:57 1993
-- Author:	Didier PIFFAULT
--		<dpf@nonox>
---Copyright:	 Matra Datavision 1993

-- signature
deferred class Vertex from MeshAlgo 

	---Purpose: Describes the data  structure for  a  vertex in  a
	--          Delaunay triangulation.

uses    Boolean from Standard,
    	Integer from Standard,
        Real from Standard,
        XY from gp,
    	DegreeOfFreedom from MeshDS


is      Initialize (x, y   : Real from Standard;
    	    	    theMov : DegreeOfFreedom from MeshDS) ; 

	Coord      (me) 
	    ---C++: return const &
    	    returns XY from gp;

	Movability (me)
    	    	    returns DegreeOfFreedom from MeshDS;

	SetMovability (me : in out; mov : DegreeOfFreedom from MeshDS);


---Purpose: For maping the Vertices.
--          Same Vertex -> Same HashCode
--          Different Vertices -> Not IsEqual but can have same HashCode 

	HashCode       (me;
    	    	    	Upper : Integer from Standard)
	---C++: function call
	    returns Integer from Standard;


	IsEqual        (me; Other : Vertex from MeshAlgo)
	---C++: alias operator ==
	    returns Boolean from Standard;


end Vertex;
