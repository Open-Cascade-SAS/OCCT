-- Created on: 1997-05-13
-- Created by: Alexander BRIVIN
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class IsoAspect from VrmlConverter inherits LineAspect from VrmlConverter

 	---Purpose: qualifies the aspect properties for  
	--          the VRML conversation of iso curves . 

uses 

    Material    from   Vrml

is

    Create
    returns mutable IsoAspect from VrmlConverter;

    ---Purpose: create a default IsoAspect. 
    --  Default value: myNumber  - 10.

    Create  (aMaterial: Material from Vrml; 
    	    	 OnOff: Boolean from Standard;
               aNumber: Integer from Standard)
    returns mutable IsoAspect from VrmlConverter;
	    

    SetNumber (me: mutable; aNumber: Integer from Standard) 
    --Purpose: defines the number of U or V isoparametric curves 
    --         to be drawn for a single face.
    is static;

    Number (me) returns Integer from Standard 
    ---Purpose: returns the number of U or V isoparametric curves drawn for a
    --          single face.
    is static;

    
fields

    myNumber: Integer from Standard;

end IsoAspect;
