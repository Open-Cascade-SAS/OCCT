-- Created on: 1997-02-12
-- Created by: Alexander BRIVIN
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Translation from Vrml 

	---Purpose:  defines a Translation of VRML specifying transform
	---          properties.
    	--  This  node  defines  a  translation  by  3D  vector. 
    	--  By  default  : 
	--    myTranslation (0,0,0) 

uses
 
    Vec  from  gp

is
 
    Create returns  Translation from Vrml; 
 
    Create  ( aTranslation  :  Vec  from  gp ) 
    	returns  Translation from Vrml; 

    SetTranslation ( me : in out;  aTranslation : Vec  from  gp );
    Translation ( me )  returns Vec  from  gp;

    Print  ( me;  anOStream: in out OStream from Standard) returns OStream from Standard;
    ---C++:  return  & 

fields
 
    myTranslation  :  Vec  from  gp;  -- Translation vector

end Translation;

