-- Created by: GG
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class IconBox from Xw inherits Window from Xw

	---Version:

	---Purpose: This class defines a X11 IconBox
	--  Warning: The IconBox is not visible at the creation time .
	--	    To show the Icon Box use the method Show () .
	--	    In this case the Icon Box appears at the DSU position
	--	    specified given in [0,1] space .
	--	    The size of the Icon Box grows depending of the number
	--	    of the Icons loaded inside .

	---References:

uses

	NameOfColor 	from Quantity,
	GraphicDevice	from Xw,
	TypeOfVisual 	from Xw,
	Handle		from Aspect,
	WindowQuality   from Xw

raises

	WindowDefinitionError	from Aspect,
	WindowError		from Aspect

is

	Create ( Device	: GraphicDevice from Xw ;
		 Name	: CString from Standard ;
		 Xc	: Real from Standard = 0.5 ;
		 Yc	: Real from Standard = 0.5 ;
		 BackColor : NameOfColor from Quantity = Quantity_NOC_MATRAGRAY;
		 aQuality : WindowQuality from Xw = Xw_WQ_SAMEQUALITY)
	returns mutable IconBox from Xw
	---Level: Public
	---Purpose: Creates a IconBox n Preferred PseudoColor Visual
	--	    defined by his Center in DSU and connects it to the
	--	    X server at the first call depending of the GraphicDevice
	--	    connexion .
	--	    ALL Icons are loaded from the Icon File Directory Name :
	--	    "[$SYMBOL]xxxxxxx[.ifd]"
	--  Warning: Raises if the Position is out of the Screen Space
	--	    or the Icon File Directory Name don't exist
	raises WindowDefinitionError from Aspect ;

	---------------------------------------------------
	-- Category: Methods to modify the class definition
	---------------------------------------------------

	LoadIcons ( me : mutable ; Name : CString from Standard ) 
					returns Integer from Standard is static;
	---Level: Public
	---Purpose: Loads Icon Box from an Other Icon File Directory Name
	--  and returns the loaded icons number.
	--  Warning: The Icons previously loaded are NOT cleared .
	---Category: Methods to modify the class definition

	Show ( me )  is static;
	---Level: Public
	---Purpose: Shows Icon Box to the screen
	--  Warning: The Icon Box is displayed at the centered position
	--	    specified at the creation time and the size depend
	--	    of the Icon number really loaded inside .

	UnloadIcons ( me : mutable ; Name : CString from Standard ) 
					returns Integer from Standard is static;
	---Level: Public
	---Purpose: Unloads All previously loaded Icons in the IconBox
        --  and returns the unloaded icons number.
	---Category: methods to modify the class definition

	Destroy ( me : mutable) is redefined ;
	---Level: Public
	---Purpose: Destroies the IconBox
	---C++: alias ~
	---Category: Methods to modify the class definition

	AddIcon ( me : mutable ; W : Window from Xw ;
	      Name : CString from Standard;
	      aWidth : Integer from Standard = 0;
	      aHeight : Integer from Standard = 0) is static;
	---Level: Public
	---Purpose: Adds an Icon of Size aWidth,aHeight given in PIXEL
	--  to the Icon Box from a FULL Existing Window
	--  NOTE that if aWidth or aHeight is 0 the default icon size is taken.
	---Category: methods to modify the class definition

	SaveIcons ( me ) returns Integer from Standard is static;
	---Level: Public
	---Purpose:  Saves all new created Icons as iconname.xwd file in the user
	--  directory and returns the saved icons number.
	
	----------------------------
	-- Category: Inquire methods
	----------------------------

	IconNumber ( me )
	returns Integer from Standard is static;
	---Level: Public
	---Purpose: Returns the Number of Icons loaded in the Icon Box .

	IconName ( me ; Index : Integer from Standard )
	returns CString from Standard
	---Level: Public
	---Purpose: Returns the Name of the N ime Icon
	--  Warning: Raises if Index if out of range depending of the
	--	    Number of Loaded Icons .
	raises WindowError from Aspect is static;

	IconSize ( me ; Name : CString from Standard ;
			Width, Height : out Integer from Standard )
	returns Boolean from Standard is static;
	---Level: Public
	---Purpose: Returns the Pixmap Size attached to the Icon Name
	--  Warning: May return FALSE if Icon doesn't exist in the IconBox .
	---Category: Inquire methods

	IconPixmap ( me ; Name : CString from Standard )
	returns Handle from Aspect is static;
	---Level: Public
	---Purpose: Returns the Pixmap attached to the Icon Name
	--  Warning: May return 0 if Icon doesn't exist in the IconBox .
	---Category: Inquire methods

	IconPixmap ( me ; Name : CString from Standard ;
			  Width, Height : Integer from Standard )
	returns Handle from Aspect is static;
	---Level: Public
	---Purpose: Returns the Centered part of the Pixmap of required Size
	--	    attached to the Icon Name
	--  Warning: May return 0 if Icon doesn't exist in the IconBox .
	---Category: Inquire methods

fields

	MyNumberOfIcons	: Integer from Standard ;

end IconBox ;
