-- Created on: 1999-11-26
-- Created by: Andrey BETENEV
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0

class ProductCategoryRelationship from StepBasic
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity ProductCategoryRelationship

uses
    HAsciiString from TCollection,
    ProductCategory from StepBasic

is
    Create returns ProductCategoryRelationship from StepBasic;
	---Purpose: Empty constructor

    Init (me: mutable; aName: HAsciiString from TCollection;
                       hasDescription: Boolean;
                       aDescription: HAsciiString from TCollection;
                       aCategory: ProductCategory from StepBasic;
                       aSubCategory: ProductCategory from StepBasic);
	---Purpose: Initialize all fields (own and inherited)

    Name (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Name
    SetName (me: mutable; Name: HAsciiString from TCollection);
	---Purpose: Set field Name

    Description (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Description
    SetDescription (me: mutable; Description: HAsciiString from TCollection);
	---Purpose: Set field Description
    HasDescription (me) returns Boolean;
	---Purpose: Returns True if optional field Description is defined

    Category (me) returns ProductCategory from StepBasic;
	---Purpose: Returns field Category
    SetCategory (me: mutable; Category: ProductCategory from StepBasic);
	---Purpose: Set field Category

    SubCategory (me) returns ProductCategory from StepBasic;
	---Purpose: Returns field SubCategory
    SetSubCategory (me: mutable; SubCategory: ProductCategory from StepBasic);
	---Purpose: Set field SubCategory

fields
    theName: HAsciiString from TCollection;
    theDescription: HAsciiString from TCollection; -- optional
    theCategory: ProductCategory from StepBasic;
    theSubCategory: ProductCategory from StepBasic;
    defDescription: Boolean; -- flag "is Description defined"

end ProductCategoryRelationship;
