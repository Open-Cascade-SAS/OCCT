-- Created on: 1994-06-01
-- Created by: Modelistation
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class SetGlobalParameter  from IGESSelect  inherits ModelModifier from IGESSelect

    ---Purpose : Sets a Global (Header) Parameter to a new value, directly given
    --           Controls the form of the parameter (Integer, Real, String
    --           with such or such form), but not the consistence of the new
    --           value regarding the rest of the file.
    --           
    --           The new value is given under the form of a HAsciiString, even
    --           for Integer or Real values. For String values, Hollerith forms
    --           are accepted but not mandatory
    --  Warning : a Null (not set) value is not accepted. For an empty string,
    --           give a Text Parameter which is empty

uses AsciiString from TCollection, HAsciiString from TCollection,
     IGESModel, CopyTool, ContextModif

is

    Create (numpar : Integer) returns mutable SetGlobalParameter;
    ---Purpose : Creates an SetGlobalParameter, to be applied on Global
    --           Parameter <numpar>

    GlobalNumber (me) returns Integer;
    ---Purpose : Returns the global parameter number to which this modifiers
    --           applies

    SetValue (me : mutable; text : mutable HAsciiString);
    ---Purpose : Sets a Text Parameter for the new value

    Value (me) returns mutable HAsciiString;
    ---Purpose : Returns the value to set to the global parameter (Text Param)


    Performing (me; ctx : in out ContextModif;
    	        target  : mutable IGESModel;
                TC      : in out CopyTool);
    ---Purpose : Specific action : only <target> is used : the form of the new
    --           value is checked regarding the parameter number (given at
    --           creation time).

    Label (me) returns AsciiString from TCollection;
    ---Purpose : Returns a text which is
    --           "Sets Global Parameter <numpar> to <new value>"

fields

    thenum : Integer;
    theval : HAsciiString from TCollection;

end SetGlobalParameter;
