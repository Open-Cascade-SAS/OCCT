-- Created on: 1998-11-23
-- Created by: Philippe MANGIN
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class IsPlanarSurface from GeomLib 

	---Purpose: Find if a surface is a planar  surface.          

uses 
  Surface  from  Geom, 
  Pln     from  gp

raises 
  NotDone  from  StdFail

is 
  Create(S  :  Surface;  Tol  :  Real  =  1.0e-7) 
  returns  IsPlanarSurface  from  GeomLib; 
   
  IsPlanar(me)  
  ---Purpose: Return if the Surface is a plan
  returns  Boolean; 
   
  Plan(me)   
  ---Purpose: Return the plan definition        
  ---C++: return const &     
  returns  Pln  from  gp 
  raises  NotDone;  --  if  <me>  is  not  Planar

fields 
  myPlan  :  Pln  from  gp; 
  IsPlan  :  Boolean;

end IsPlanarSurface;
