-- File:        ProductType.cdl
-- Created:     Mon Dec  4 12:02:30 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWProductType from RWStepBasic

	---Purpose : Read & Write Module for ProductType

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     ProductType from StepBasic,
     EntityIterator from Interface

is

	Create returns RWProductType;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable ProductType from StepBasic);

	WriteStep (me; SW : in out StepWriter; ent : ProductType from StepBasic);

	Share(me; ent : ProductType from StepBasic; iter : in out EntityIterator);

end RWProductType;
