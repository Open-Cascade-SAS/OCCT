-- Created on: 1993-06-17
-- Created by: Christian CAILLET
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DispatchControl  from Transfer  inherits CopyControl from Interface

    ---Purpose : This is an auxiliary class for TransferDispatch, which allows
    --           to record simple copies, as CopyControl from Interface, but
    --           based on a TransientProcess. Hence, it allows in addition
    --           more actions (such as recording results of adaptations)

uses Transient, TransientProcess, InterfaceModel

raises InterfaceError

is

    Create (model : InterfaceModel; TP : mutable TransientProcess)
    	returns mutable DispatchControl;
    ---Purpose : Creates the DispatchControl, ready for use

    TransientProcess (me) returns mutable TransientProcess;
    ---Purpose : Returns the content of the DispatchControl : it can be used
    --           for a direct call, if the basic methods do not suffice
    ---C++ : return const &

    StartingModel (me) returns any InterfaceModel;
    ---Purpose : Returns the Model from which the transfer is to be done
    ---C++ : return const &

    	--  Now, inherited methods used for Copy (the minimum set)

    Clear (me : mutable);
    ---Purpose : Clears the List of Copied Results

    Bind (me : mutable; ent : Transient; res : mutable Transient)
    ---Purpose : Binds a (Transient) Result to a (Transient) Starting Entity
    	raises InterfaceError;
    --           Error if <ent> is already bound

    Search (me; ent : Transient; res : out mutable Transient)
    	returns Boolean;
    ---Purpose : Searches for the Result bound to a Starting Entity
    --           If Found, returns True and fills <res>
    --           Else, returns False and nullifies <res>

fields

    theTP    : TransientProcess;
    themodel : InterfaceModel;

end DispatchControl;
