-- Created on: 2001-05-03
-- Created by: Igor FEOKTISTOV
-- Copyright (c) 2001-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

class Limitation from QANewModTopOpe inherits MakeShape from BRepBuilderAPI

---Purpose: provides  cutting  shape  by  face  or  shell;

uses

    Shape from TopoDS, 
    ListOfShape from TopTools, 
    ModeOfLimitation  from  QANewModTopOpe, 
    State  from  TopAbs,  
    CutPtr  from  QANewModTopOpe, 
    CommonPtr  from  QANewModTopOpe
is 
  
    Create(theObjectToCut,  theCutTool : Shape from TopoDS;
    	    theMode : ModeOfLimitation  from  QANewModTopOpe = QANewModTopOpe_Forward)
    ---Purpose: initializes and  fills data structure for  cutting and
    --          makes  cutting according to orientation theCutTool and
    --          theMode.
    --          if theCutTool is not face or shell does nothing.
    
    returns Limitation from QANewModTopOpe;    
     
    Cut(me  :  in  out);
    ---Purpose: makes cutting  according to  orientation theCutTool
    --          and  current value   of  myMode.  Does nothing  if
    --          result already  exists.

    SetMode(me  :  in  out;  theMode  :  ModeOfLimitation  from  QANewModTopOpe); 
     
    GetMode(me)  returns  ModeOfLimitation  from  QANewModTopOpe;  
     
    Shape1(me)  returns  Shape  from  TopoDS
    ---Purpose: Returns the first shape.
    ---C++: return const &
    ---Level: Public
    is static;
     
    Shape2(me)  returns  Shape  from  TopoDS
    ---Purpose: Returns the second shape.
    ---C++: return const &
    ---Level: Public
    is static; 
    
    Modified (me: in out; S : Shape from TopoDS)
    	---Purpose: Returns the list  of shapes modified from the shape
    	--          <S>. 
        ---C++: return const & 
        ---Level: Public
    returns ListOfShape from TopTools
    is redefined;
 
    Modified2 (me: in out;  
    	    	aS : Shape from TopoDS) 
    	returns ListOfShape from TopTools;
    ---Purpose: Returns the list  of shapes modified from the shape <S>.
    ---         For use in BRepNaming.
    ---C++: return const & 
    ---Level: Public

    Generated (me: in out; S : Shape from TopoDS)
    	returns ListOfShape from TopTools
	is redefined;
    	---Purpose: Returns the list  of shapes generated from the shape <S>.
    	---         For use in BRepNaming.
    	---C++:  return const &
    
    HasModified (me)
    	returns Boolean from Standard
	is virtual;
    	---Purpose: Returns true if there is at least one modified shape.
    	---         For use in BRepNaming.

    HasGenerated (me)
    	returns Boolean from Standard
	is virtual;
    	---Purpose: Returns true if there is at least one generated shape.
    	---         For use in BRepNaming.

    HasDeleted (me)
    	returns Boolean from Standard
	is virtual;
    	---Purpose: Returns true if there is at least one deleted shape.
    	---         For use in BRepNaming.

    IsDeleted (me: in out; S : Shape from TopoDS)
    returns Boolean from Standard
    is redefined;
      
    Delete(me  :  in  out)  is  redefined; 
    ---C++:  alias  "Standard_EXPORT  ~QANewModTopOpe_Limitation()  {Delete();}"
  

fields 

    myResultFwd     :  Shape  from  TopoDS;  
    myResultRvs     :  Shape  from  TopoDS;  
    myObjectToCut   :  Shape  from  TopoDS;  
    myCutTool       :  Shape  from  TopoDS;  
    myCut           :  CutPtr  from  QANewModTopOpe;
    myCommon        :  CommonPtr  from  QANewModTopOpe;
    myFwdIsDone     :  Boolean  from  Standard;
    myRevIsDone     :  Boolean  from  Standard;  
    myMode          :  ModeOfLimitation  from  QANewModTopOpe;
    
end  Limitation;
