-- Created on: 1998-05-20
-- Created by: Christian CAILLET
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




deferred class SignText  from MoniTool    inherits TShared
 
        ---Purpose : Provides the basic service to get a text which identifies
        --           an object in a context
        --           It can be used for other classes (general signatures ...)
        --           It can also be used to build a message in which an object
        --           is to be identified
 
uses CString, Transient, AsciiString from TCollection
 
is
 
    Name (me) returns CString  is deferred;
    ---Purpose : Returns an identification of the Signature (a word), given at
    --           initialization time

    TextAlone (me; ent : any Transient)
    	returns AsciiString from TCollection  is virtual;
    ---Purpose : Gives a text as a signature for a transient object alone, i.e.
    --           without defined context.
    --           By default, calls Text with undefined context (Null Handle) and
    --           if empty, then returns DynamicType

    Text (me; ent : any Transient; context : any Transient)
    	returns AsciiString from TCollection  is deferred;
    ---Purpose : Gives a text as a signature for a transient object in a context
    --           If the context is senseless, it can be given as Null Handle
    --           empty result if nothing to give (at least the DynamicType could
    --           be sent ?)

end SignText;
