-- Created by: TCL
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class DrawSymbol from Prs2d inherits Line from Graphic2d

	---Purpose: The primitive symbol for drawing

uses

	Drawer		    from Graphic2d,
	GraphicObject	from Graphic2d, 
    TypeOfSymbol    from Prs2d,
    FStream         from Aspect

raises

	SymbolDefinitionError from Prs2d

is
	-------------------------
	-- Category: Constructor
	-------------------------

	Create( aGO       : GraphicObject from Graphic2d;
		    aSymbType : TypeOfSymbol  from Prs2d;
		    aX, aY    : Real          from Standard;
		    aWidth    : Real          from Standard = 10.0;
		    aHeight   : Real          from Standard = 10.0;
		    anAngle   : Real          from Standard = 0.0 )
	 returns mutable DrawSymbol from Prs2d 
     raises SymbolDefinitionError from Prs2d;

	---Level: Public
	---Purpose: Creates the predefined marker index <anIndex> 
	--	    at position <aX>, <aY> and size <aWidth>,<aHeight>.
    ---Category: Constructor
	---Purpose:  Trigger  -   Raises SymbolDefinitionError if the
	--	    symbol type isn't defined,
	--      or the symbol size < aWidth, aHeight > is null.

	----------------------------------------------------
	-- Category: Draw and Pick
	----------------------------------------------------

	Draw( me: mutable; aDrawer: Drawer from Graphic2d ) is static protected;
	---Level: Internal
	---Purpose: Draws the symbol <me>.

	Pick( me : mutable; 
          X, Y       : ShortReal from Standard;
		  aPrecision : ShortReal from Standard;
		  aDrawer    : Drawer from Graphic2d ) returns Boolean from Standard
	  is static protected;
	---Level: Internal
	---Purpose: Returns Standard_True if the symbol <me> is picked,
	--	    Standard_False if not.
	--  Warning: Checks only if the point <X>, <Y> is in the
	--	    boundary rectangle of <me>

   Save( me; aFStream: in out FStream from Aspect ) is virtual;

fields

	myTypeSymb : TypeOfSymbol from Prs2d;
	myX        : ShortReal from Standard;
	myY        : ShortReal from Standard;
	myWidth    : ShortReal from Standard;
	myHeight   : ShortReal from Standard;
	myAngle    : ShortReal from Standard;

end Marker from Graphic2d;
