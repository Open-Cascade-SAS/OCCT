-- Created on: 1993-04-06
-- Created by: Philippe DAUTRY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class BezierCurve from PGeom2d inherits BoundedCurve from PGeom2d

        ---Purpose : Defines a rational or non rational Bezier curve.
        --         
	---See Also : BezierCurve from Geom2d.

uses  HArray1OfReal from PColStd,
      HArray1OfPnt2d  from PColgp

is 


  Create returns mutable BezierCurve from PGeom2d;
        ---Purpose : Creates a non rational  Bezier curve with default
        --         values.
	---Level: Internal 


  Create(aPoles    : HArray1OfPnt2d;
         aWeights  : HArray1OfReal;
	 aRational : Boolean from Standard)
     returns mutable BezierCurve from PGeom2d;
        ---Purpose : Creates a non rational Bezier curve with a set of
        --         poles aCurvePoles and a set of weights aPoleWeight.
	---Level: Internal 


  Rational (me: mutable; aRational: Boolean from Standard);
        ---Purpose : Set the value of the field rational with <aRational>.
	---Level: Internal 


  Rational (me) returns Boolean;
        ---Purpose : Returns the value of the field rational.
	---Level: Internal 


  Poles (me: mutable; aPoles : HArray1OfPnt2d from PColgp);
        ---Purpose : Set the value of the field poles with <aPoles>.
	---Level: Internal 


  Poles (me) returns HArray1OfPnt2d from PColgp;
        ---Purpose : Returns the value of the field poles.
	---Level: Internal 


  Weights (me: mutable; aWeights : HArray1OfReal from PColStd);
        ---Purpose : Set the value of the field weights.
	---Level: Internal 


  Weights (me)returns HArray1OfReal from PColStd;
        ---Purpose : Returns the value of the field weights.
	---Level: Internal 


fields

   rational : Boolean from Standard;
   poles    : HArray1OfPnt2d  from PColgp;
   weights  : HArray1OfReal from PColStd;

end;
