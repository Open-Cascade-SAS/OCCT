-- File:	Dynamic_EnumerationParameter.cdl
-- Created:	Thu Feb  3 14:44:37 1994
-- Author:	Gilles DEBARBOUILLE
--		<gde@metrox>
---Copyright:	 Matra Datavision 1994


generic class EnumerationParameter from Dynamic (Enum as any)

inherits

    Parameter from Dynamic     
    
    ---Purpose: This  generic class defines  a  parameter with a given
    --          enumeration.  For correct use an instanciation of this
    --          class,  the  Convert  method  must  be  defined.  This
    --          method is automaticaly called by the constructor which
    --          takes a  CString  as value for  the  enumeration.  The
    --          prototype  of the Convert method  must be described as
    --          follows :
    --          
    --          void Convert(const Standard_CString,Enum);
    --          
    --          The  prototype  and the body of  this   method, can be
    --          written  in   the  file   <mypackage.cxx>   where  the
    --          enumeration  is described.    No declaration  of   the
    --          Convert method in any .cdl file is necessary.


uses
    CString from Standard,
    OStream from Standard 

is

    Create(aparameter : CString from Standard)
    
    ---Level: Public 
    
    ---Purpose: Creates an  EnumerationParameter  of  <aparameter>  as
    --          name.

    returns mutable EnumerationParameter from Dynamic;

    Create(aparameter : CString from Standard; avalue : Enum)
    
    ---Level: Public 
    
    ---Purpose: Creates  an  EnumerationParameter  of  <aparameter> as
    --          name and <avalue> as value.

    returns mutable EnumerationParameter from Dynamic;
    
    Create(aparameter , avalue : CString from Standard) 

    ---Level: Public 
    
    ---Purpose: Creates an  EnumerationParameter  of  <aparameter>  as
    --          name  and <avalue> as value. The user has to define  a
    --          Convert method to translate  the string <avalue> in an
    --          enumeration term.

    returns mutable EnumerationParameter from Dynamic;
    
    Value(me) returns Enum
    
    ---Level: Public 
    
    ---Purpose: Returns the enumeration value <thevalue>.
    
    is static;
    
    Value (me : mutable ; avalue : Enum)
    
    ---Level: Public 
    
    ---Purpose: Sets the field <thevalue> with the enumeration value <avalue>

    is static;
    
    Dump(me ; astream : in out OStream from Standard)
    
    ---Level: Internal 
    
    ---Purpose: useful for debugging.
    
    is redefined;
    
fields

    thevalue : Enum;

end EnumerationParameter;
