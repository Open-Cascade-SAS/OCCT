-- Created on: 1992-06-22
-- Created by: Gilles DEBARBOUILLE
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Lexicon from Units 

inherits

    TShared from MMgt 

	---Purpose: This class defines a lexicon useful to analyse and
	--          recognize the  different key words  included  in a
	--          sentence.  The lexicon is stored  in a sequence of
	--          tokens.

uses

    HAsciiString   from TCollection,
    AsciiString    from TCollection,
    TokensSequence from Units

is

    Create returns mutable Lexicon from Units;
    
    ---Level: Internal 
    
    ---Purpose: Creates an empty instance of Lexicon.
    
    Creates(me : mutable ; afilename : CString)
    
    ---Level: Internal 
    
    ---Purpose: Reads the file <afilename> to create a sequence  of tokens
    --          stored in <thesequenceoftokens>.
    
    is static;
    
    Sequence(me) returns any TokensSequence from Units
    
    ---Level: Internal 
    
    ---C++: inline
    
    ---Purpose: Returns the first item of the sequence of tokens.
    
    is static;
    
    FileName(me) returns AsciiString from TCollection
    
    ---Level: Internal 
    
    ---Purpose: Returns in a AsciiString from TCollection the name of the file.
    
    is static;
    
    UpToDate(me) returns Boolean
    
    ---Level: Internal 
    
    ---Purpose: Returns true if  the  file has not  changed  since the
    --          creation   of   the  Lexicon   object.   Returns false
    --          otherwise.

    is virtual;
    
    AddToken(me : mutable ; aword , amean : CString ; avalue : Real)
    
    ---Level: Internal 
    
    ---Purpose: Adds to the lexicon a new token with <aword>, <amean>,
    --          <avalue>  as  arguments.  If there is  already a token
    --          with   the  field  <theword>  equal    to <aword>, the
    --          existing token is updated.
    
    is static;
    
    Dump(me)
    
    ---Level: Internal 
    
    ---C++: inline
    ---Purpose: Useful for debugging.

    is virtual;
    
fields

    thefilename         : HAsciiString from TCollection;
    thetime             : Time from Standard;
    thesequenceoftokens : TokensSequence from Units;

end Lexicon;
