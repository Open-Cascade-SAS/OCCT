-- Created on: 1997-01-08
-- Created by: VAUTHIER Jean-Claude
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package QADNaming 

	---Purpose: 

	--           FOR OLD TOPOLOGY ONLY!
uses 
    Draw,
    TCollection, 
    TColStd,
    TDF,
    TNaming,
    TopoDS,
    TopTools
is
         
    class DataMapOfShapeOfName instantiates
    	DataMap from TCollection(Shape          from TopoDS,
	    	    	    	 AsciiString    from TCollection,
                                 ShapeMapHasher from TopTools);  				  			       								   
    CurrentShape (ShapeEntry      : CString  from Standard; 
    	    	  Data            : Data     from TDF)
    returns Shape from TopoDS;		  

    GetShape (ShapeEntry  :        CString     from Standard; 
    	      Data        :        Data        from TDF;
    	      Shapes      : in out ListOfShape from TopTools);
    

    GetEntry (Shape      : in     Shape   from TopoDS; 
              Data       : in     Data    from TDF; 
              Status     : in out Integer from Standard)
    	---Purpose: Status = 0  Not  found, 
    	--          Status = 1  One  shape,
    	--          Status = 2  More than one shape. 
    returns AsciiString from TCollection;
    
    Entry (theArguments : Address from Standard;
    	   theLabel : in out Label from TDF) returns Boolean from Standard;
    --- Purpose: returns label by first two arguments (df and entry string)

    AllCommands        (DI : in out Interpretor from Draw);
    
    BasicCommands      (DI : in out Interpretor from Draw);
    ---Purpose: commands relatives to NamedShape

    BuilderCommands    (DI : in out Interpretor from Draw);
    ---Purpose: loading NamedShape to the Data Framework

    IteratorsCommands  (DI : in out Interpretor from Draw);
    ---Purpose: loading NamedShape to the Data Framework

    ToolsCommands      (DI : in out Interpretor from Draw);
    
    SelectionCommands  (DI : in out Interpretor from Draw);
    ---Purpose: commands relatives to Naming 

end QADNaming;




