-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class AutoDesignDateAndPersonAssignment from StepAP214 

inherits PersonAndOrganizationAssignment from StepBasic

uses

	HArray1OfAutoDesignDateAndPersonItem from StepAP214, 
	AutoDesignDateAndPersonItem from StepAP214, 
	PersonAndOrganization from StepBasic,
	PersonAndOrganizationRole from StepBasic
is

	Create returns mutable AutoDesignDateAndPersonAssignment;
	---Purpose: Returns a AutoDesignDateAndPersonAssignment


	Init (me : mutable;
	      aAssignedPersonAndOrganization : mutable PersonAndOrganization from StepBasic;
	      aRole : mutable PersonAndOrganizationRole from StepBasic) is redefined;

	Init (me : mutable;
	      aAssignedPersonAndOrganization : mutable PersonAndOrganization from StepBasic;
	      aRole : mutable PersonAndOrganizationRole from StepBasic;
	      aItems : mutable HArray1OfAutoDesignDateAndPersonItem from StepAP214) is virtual;

	-- Specific Methods for Field Data Access --

	SetItems(me : mutable; aItems : mutable HArray1OfAutoDesignDateAndPersonItem);
	Items (me) returns mutable HArray1OfAutoDesignDateAndPersonItem;
	ItemsValue (me; num : Integer) returns AutoDesignDateAndPersonItem;
	NbItems (me) returns Integer;

fields

	items : HArray1OfAutoDesignDateAndPersonItem from StepAP214; -- a SelectType

end AutoDesignDateAndPersonAssignment;
