-- Created on: 1993-01-09
-- Created by: CKY / Contract Toubro-Larsen ( TCD )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Planar from IGESDraw  inherits IGESEntity

        ---Purpose: defines IGESPlanar, Type <402> Form <16>
        --          in package IGESDraw
        --
        --          Indicates that a collection of entities is coplanar.The
        --          entities may be geometric, annotative, and/or structural.

uses

        TransformationMatrix    from IGESGeom,
        HArray1OfIGESEntity from IGESData

raises OutOfRange

is

        Create returns mutable Planar;

        -- Specific Methods pertaining to the class

        Init (me                    : mutable;
              nbMats                : Integer;
              aTransformationMatrix : TransformationMatrix;
              allEntities           : HArray1OfIGESEntity);
        ---Purpose : This method is used to set the fields of the class Planar
        --       - nbMats                : Number of Transformation matrices
        --       - aTransformationMatrix : Pointer to the Transformation matrix
        --       - allEntities           : Pointers to the entities specified

        NbMatrices (me) returns Integer;
        ---Purpose : returns the number of Transformation matrices in <me>

        NbEntities (me) returns Integer;
        ---Purpose : returns the number of Entities in the plane pointed to by this
        -- associativity

        IsIdentityMatrix (me) returns Boolean;
        ---Purpose : returns True if TransformationMatrix is Identity Matrix,
        -- i.e:- No Matrix defined.

        TransformMatrix (me) returns TransformationMatrix;
        ---Purpose : returns the Transformation matrix moving data from the XY plane
        -- into space or zero

        Entity (me; EntityIndex : Integer) returns IGESEntity
        raises OutOfRange;
        ---Purpose : returns the Entity on the specified plane, indicated by EntityIndex
        -- raises an exception if EntityIndex <= 0 or
        -- EntityIndex > NbEntities()

fields

--
-- Class    : IGESDraw_Planar
--
-- Purpose  : Declaration of the variables specific to a Planar Entity.
--
-- Reminder : A Planar Entity is defined by :
--                    - Number of Transformation matrices
--                    - Pointer to the Transformation matrix
--                    - Pointers to the entities specified
--

        theNbMatrices           : Integer;

        theTransformationMatrix : TransformationMatrix;

        theEntities             : HArray1OfIGESEntity;

end Planar;
