-- Created on: 1993-02-05
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



package Contap

	---Purpose: 

uses Standard,StdFail,MMgt, GeomAbs, TopAbs, TCollection, gp, TColgp,
     math, IntSurf, IntStart, IntWalk,
     Geom2d, TColStd, Geom, Adaptor3d,  Adaptor2d

is

    deferred generic class ArcTool;        -- template class
    
    deferred generic class SurfaceTool;    -- template class
    
    deferred generic class TopolTool;      -- template class
    
    generic class Point;

    generic class Line;

    generic class SurfFunction;
    
    generic class ArcFunction;
    
    generic class SurfProps;

    generic class ContourGen, ThePoint,TheSequenceOfPoint,TheHSequenceOfPoint,
                              TheLine, TheSequenceOfLine,
			      TheSurfProps, TheSurfFunction, TheArcFunction,
                              TheSearch, TheIWalking, TheSearchInside;
    	    	    	      ---TheLineConstructor;

    class ContAna;		   

    enumeration TFunction is
    	ContourStd,
	ContourPrs,
	DraftStd,
	DraftPrs
    end TFunction;	

    enumeration IType is  -- a replacer dans IntSurf et fusionner avec IntPatch
    -- type of the line of contour

    	Lin,       -- pour conflit avec deferred class Line
    	Circle,
        Walking,
    	Restriction
    end IType;
	
    generic class HContToolGen;
    
    generic class HCurve2dToolGen;
    
    class HCurve2dTool instantiates 
    	HCurve2dToolGen from Contap ( 
	    HCurve2d from Adaptor2d);

    class HContTool instantiates 
        HContToolGen from Contap (
    	 HVertex       from Adaptor3d,
	 HCurve2d      from Adaptor2d,
	 HSurface      from Adaptor3d,
    	 HCurve2dTool  from Contap,
	 HSurfaceTool  from Adaptor3d);
	 
    class Contour instantiates ContourGen from Contap
    	(HVertex       from Adaptor3d,
	 HCurve2d      from Adaptor2d,
	 HSurface      from Adaptor3d,
	 HCurve2dTool  from Contap,
	 HSurfaceTool  from Adaptor3d,
	 HContTool     from Contap,
	 TopolTool     from Adaptor3d);


end Contap;
