-- Created on: 1993-03-23
-- Created by: BBL
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ColorMapEntry from Aspect inherits Storable from Standard

	---Version: 0.0

	---Purpose: This class defines a colormap entry.
	--	    A colormap entry is an association between
	--	    a RGB object and a index in the colormap.
	---Keywords:
	---Warning:
	---References:

uses
	Color from Quantity

raises
	OutOfRange 	from Standard,
	BadAccess 	from Aspect

is
	Create
	returns ColorMapEntry from Aspect;
	---Level: Public
	---Purpose: Creates an unallocated colormap entry
	
	Create ( index : in Integer from Standard;
		 rgb : in Color from Quantity)
 	returns ColorMapEntry;
	---Level: Public
	---Purpose: Creates an allocated colormap entry

	Create ( entry : in ColorMapEntry from Aspect )
 	returns ColorMapEntry
	---Level: Public
	---Purpose: Creates an allocated colormap entry.
	--  Warning: Raises error if the colormap entry <entry>
	--	    is unallocated.
	raises BadAccess from Aspect;

	SetValue ( me: in out; index : in Integer from Standard;
			rgb : in Color from Quantity );
	---Level: Public
 	---Purpose: Sets colormap entry value and allocates it.
 
	SetValue ( me: in out; entry : in ColorMapEntry from Aspect);
	---Level: Public
 	---Purpose: Sets colormap entry value and allocates it.
	---C++: alias operator =
 
	SetColor ( me: in out; rgb : in Color from Quantity );
	---Level: Public
 	---Purpose: Sets color <rgb> of colormap entry.

	Color ( me : in ) returns Color from Quantity
	---Warning: Raises error if the colormap entry is unallocated .
	raises BadAccess from Aspect;
	---C++: return const & 

	SetIndex ( me: in out; index : in Integer from Standard);
	---Level: Public
 	---Purpose: Sets index value of a colormap entry.

	Index ( me : in ) returns Integer from Standard 
	---Warning: Raises error if the colormap entry is unallocated .
	raises BadAccess from Aspect;

	Free ( me : in out );
	---Level: Public
	---Purpose: Unallocates the colormap entry.

	IsAllocated ( me : in )
	returns Boolean from Standard;
	---Level: Public
	---Purpose: Returns True if the colormap entry is allocated.
	--  Warning: A colormap entry is allocated when the color and
	--	    the index is defined.

        Dump( me : in ) ;
	---Level: Internal

fields
	allocated 	: Boolean from Standard;
	mycolor		: Color from Quantity;
	myindex 	: Integer from Standard;
	myColorIsDef	: Boolean from Standard;
	myIndexIsDef	: Boolean from Standard;

end ColorMapEntry from Aspect;
