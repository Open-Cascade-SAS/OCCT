-- File:	TCompound.cdl
-- Created:	Mon Dec 17 11:18:44 1990
-- Author:	Remi Lequette
--		<rle@topsn3>
---Copyright:	 Matra Datavision 1990, 1992



class TCompound from PTopoDS inherits TShape from PTopoDS

	---Purpose: A topological Compound object containing shapes.

uses
    ShapeEnum from TopAbs

is
    Create returns mutable TCompound from PTopoDS;
	---Purpose: the new TCompound is empty.
    ---Level: Internal 
    	
    ShapeType(me) returns ShapeEnum from TopAbs;
    ---Level: Internal 

end TCompound;

