-- Created on: 1992-09-29
-- Created by: Didier PIFFAULT
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class InterferencePolyhedron from IntPatch inherits Interference from Intf

	---Purpose: Computes the  interference between two polyhedra or the
	--          self interference of a polyhedron. Points of intersection,
  --          polylines  of intersection and zones of tangence.

uses    Pnt               from gp,
        XYZ               from gp,
    	Box               from Bnd,
    	SectionPoint      from Intf,
    	SeqOfSectionPoint from Intf,
    	SectionLine       from Intf,
    	SeqOfSectionLine  from Intf,
    	TangentZone       from Intf,
    	SeqOfTangentZone  from Intf,
        Polyhedron        from IntPatch,
        PolyhedronTool    from IntPatch

is

-- Interface :

    Create          returns InterferencePolyhedron from IntPatch;
    ---Purpose: Constructs an empty interference of Polyhedron.

    Create         (Obje1  : in Polyhedron from IntPatch;
    	    	    Obje2  : in Polyhedron from IntPatch) 
    	            returns InterferencePolyhedron from IntPatch;
    ---Purpose: Constructs  and computes  an  interference between  the two
    --          Polyhedra.

    Create         (Obje   : in Polyhedron from IntPatch) 
    	            returns InterferencePolyhedron from IntPatch;
    ---Purpose: Constructs  and  computes   the self   interference  of   a
    --          Polyhedron.

    Perform        (me     : in out;
    	    	    Obje1  : in Polyhedron from IntPatch;
    	    	    Obje2  : in Polyhedron from IntPatch);
    ---Purpose: Computes the interference between the two Polyhedra.

    Perform        (me     : in out;
    	    	    Obje   : in Polyhedron from IntPatch);
    ---Purpose: Computes the self interference of a Polyhedron.

-- Implementation :

    Interference   (me     : in out;
    	    	    Obje1  : in Polyhedron from IntPatch)
    	    	    is private;
    Interference   (me     : in out;
    	    	    Obje1  : in Polyhedron from IntPatch;
     	    	    Obje2  : in Polyhedron from IntPatch)
    	    	    is private;
    ---Purpose: Compares the bounding volumes between the facets of <Obje1>
    --          and the facets of <Obje2> and intersects the facets when the
    --          bounding volumes have a common part.

    Intersect      (me     : in out;
		    TriF   : in Integer from Standard;
    	    	    Obje1  : in Polyhedron from IntPatch;
		    TriS   : in Integer from Standard;
    	    	    Obje2  : in Polyhedron from IntPatch)
    	    	    is private;
    ---Purpose: Computes  the intersection between    the  facet <Tri1>  of
    --          <FirstPol> and the facet <Tri2> of <SecondPol>.

    TangentZoneValue
    	    	   (me;
    	    	    TheTZ  : in out TangentZone from Intf;
		    Obje1  : Polyhedron from IntPatch;
		    Tri1   : Integer from Standard;
    	    	    Obje2  : Polyhedron from IntPatch;
    	    	    Tri2   : Integer from Standard)
		    returns Boolean from Standard
    	    	    is private;
    ---Purpose: Computes the  zone of tangence between the  facet <Tri1> of
    --          <FirstPol> and the facet <Tri2> of <SecondPol>.

    CoupleCharacteristics (me: in out;
            FirstPol: Polyhedron from IntPatch;
            SeconPol: Polyhedron from IntPatch) is private;
fields
    OI       : Integer from Standard[3]; -- index des sommets de l objet
    TI       : Integer from Standard[3]; -- index des sommets du tool
    dpOpT    : Real from Standard[3, 3]; -- distance point Objet - point Tool
    dpOeT    : Real from Standard[3, 3]; -- distance point Objet - edge  Tool
    deOpT    : Real from Standard[3, 3]; -- distance edge  Objet - point Tool
    voo      : XYZ from gp[3];           -- vecteur point point Obje
    vtt      : XYZ from gp[3];           -- vecteur point point Tool
    Incidence: Real from Standard;       -- angle entre les deux plans

end InterferencePolyhedron;
