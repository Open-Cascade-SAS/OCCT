-- Created on: 1993-06-08
-- Created by: Laurent BOURESCHE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Tool from BRepSweep -- as Tool from Sweep

    ---Purpose: Provides  the  indexation and type  analysis  services
    --          required by the TopoDS generating Shape of BRepSweep.
    --          

uses

    Shape from TopoDS,
    IndexedMapOfShape from TopTools,
    ShapeEnum from TopAbs,
    Orientation from TopAbs

raises 

    OutOfRange from Standard

is

    Create(aShape: Shape from TopoDS);
	---Purpose: Initialize the tool  with <aShape>.  The IndexTool
	--          must prepare an indexation for  all  the subshapes
	--          of this shape.

    NbShapes(me) returns Integer
	---Purpose: Returns the number of subshapes in the shape.
    is static;

    Index(me; aShape : Shape from TopoDS) returns Integer
	---Purpose: Returns the index of <aShape>.
    is static;
    
    Shape(me; anIndex : Integer from Standard) returns Shape from TopoDS
	---Purpose: Returns the Shape at Index anIdex.
    is static;
    
    Type(me; aShape : Shape from TopoDS) returns ShapeEnum from TopAbs
	---Purpose: Returns the type of <aShape>.
    is static;

    Orientation (me; aShape : Shape from TopoDS) 
    returns Orientation from TopAbs
	---Purpose: Returns the Orientation of <aShape>.
    is static;

    SetOrientation (me; 
    	    	    aShape : in out Shape from TopoDS; 
    	    	    Or     : Orientation  from  TopAbs) 
	---Purpose: Set the Orientation of <aShape> with Or.
    is static;

fields

    myMap : IndexedMapOfShape from TopTools;
    
end Tool from BRepSweep;



