-- Created on: 2002-10-29
-- Created by: Michael SAZONOV
-- Copyright (c) 2002-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class ADriverTable from BinMDF inherits TShared from MMgt

        ---Purpose: A driver table is an object building links between
        --          object types and object drivers. In the
        --          translation process, a driver table is asked to
        --          give a translation driver for each current object
        --          to be translated.

uses
    Type               from Standard,
    ADriver            from BinMDF,    
    TypeADriverMap     from BinMDF,
    IndexedMapOfTransient from TColStd,
    SequenceOfAsciiString from TColStd,
    TypeIdMap from BinMDF

is
    Create returns mutable ADriverTable from BinMDF;
        ---Purpose: Constructor

    AddDriver(me : mutable; theDriver : ADriver from BinMDF);
        ---Purpose: Adds a translation driver <theDriver>.

    AssignId(me : mutable; theType	: Type from Standard;
			   theId	: Integer from Standard)
    	is private;
	---C++: inline
        ---Purpose: Assigns the ID to the driver of the Type

    AssignIds(me : mutable; theTypes	: IndexedMapOfTransient from TColStd);
        ---Purpose: Assigns the IDs to the drivers of the given Types.
        --          It uses indices in the map as IDs.
        --          Useful in storage procedure.

    AssignIds(me : mutable; theTypeNames : SequenceOfAsciiString from TColStd);
        ---Purpose: Assigns the IDs to the drivers of the given Type Names;
        --          It uses indices in the sequence as IDs.
        --          Useful in retrieval procedure.

    GetDriver(me; theType     : Type from Standard;
                  theDriver   : in out ADriver from BinMDF)
        returns Integer from Standard;
	---C++: inline
        ---Purpose: Gets a driver <theDriver> according to <theType>.
        --          Returns Type ID if the driver was assigned an ID; 0 otherwise.

    GetDriver(me; theTypeId   : Integer from Standard)
    	returns ADriver from BinMDF;
	---C++: inline
        ---Purpose: Returns a driver according to <theTypeId>.
        --          Returns null handle if a driver is not found

fields
    myMap	: TypeADriverMap from BinMDF;
    myMapId	: TypeIdMap from BinMDF;

end ADriverTable;
