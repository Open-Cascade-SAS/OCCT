-- Created on: 1991-03-28
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package IntWalk

	---Purpose: This package defines the "walking" (marching) algorithmes
	--          for the intersection between two surfaces.
	--          One of the surfaces is a parametric one.
	--          If the other is an implicit one, the "IWalking" class will
	--          be used.
	--          If both surfaces are parametric, the "PWalking" class will
	--          be used.

        ---Level: Internal
        --
        -- All the methods of the classes of this package are Internal.
	-- 
uses   
     Standard, MMgt, TCollection, TColStd, gp, math, StdFail, IntSurf, IntImp

is

    enumeration StatusDeflection is 
                PasTropGrand, PointConfondu, ArretSurPointPrecedent,
                ArretSurPoint, OK;

-- StepTooGreat, ConfusedPoint, StopOnPreviousPoint, StopOnPoint, OK
    
--class of result objects marching on a biparametric surface

    generic class IWLine;
    
    
--algorithm marching/solution

    generic class IWalking, TheIWLine, SequenceOfIWLine;
    
    imported VectorOfWalkingData;
    ---Purpose: Defines a dynamic vector of work data.
    
    imported VectorOfInteger;
    ---Purpose: Defines a dynamic vector of integer.

    
--algorithm/solution for a marching on intersection between
-- 2 biparametric surfaces

    generic class PWalking, TheInt2S;


end IntWalk;
