-- Created by: DAUTRY Philippe
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

--      	-------

---Version:	0.0
--Version	Date		Purpose
--		0.0	Feb 10 1997	Creation



package DDF 

	---Purpose: Provides facilities to manipulate data framework
	--          in a Draw-Commands environment.

uses

    Standard,
    Draw,
    TCollection,
    TDF

is

    -- ----------------------------------------------------------------------
    -- Classes
    -- ----------------------------------------------------------------------

    class Data;
    	---Purpose : Encapsulates a data framework from TDF.

    class Browser;
    	---Purpose : Browses a data framework from TDF.

    class Transaction;
	---Purpose: Encapsulates a Transaction from TDF.

    class TransactionStack
    	instantiates Stack from TCollection (Transaction from DDF);

    -- ----------------------------------------------------------------------
    -- Package methods
    -- ----------------------------------------------------------------------


    GetDF (Name     : in out CString from Standard; 
           DF       : in out Data    from TDF;
           Complain : in     Boolean from Standard = Standard_True)
    returns Boolean;
   	---Purpose: Search in draw  directory the framewok  identified
   	--          by its name <Name>. returns True if found. In that
   	--          case <DF> is setted.


    FindLabel (DF      : in     Data    from TDF; 
    	      Entry    : in     CString from Standard;
	      Label    : in out Label   from TDF;
              Complain : in     Boolean from Standard = Standard_True)
    returns Boolean;
   	---Purpose: Search in <DF>  the label identified by its  entry
   	--          <Entry>.  returns  <True> if  found. In  that case
   	--          <Label> is setted.

    AddLabel (DF      : in     Data    from TDF;
    	      Entry   : in     CString from Standard; 
    	      Label   : in out Label   from TDF)
    returns  Boolean;
    	---Purpose : Search in <DF> the  label identified by its entry
    	--         <Entry>.   if label doesn't  exist, create  and add
    	--         the Label in <DF>. In that case return True.


    Find (DF       : in     Data      from TDF;
          Entry    : in     CString   from Standard;
    	  ID       : in     GUID      from Standard;
          A        : in out Attribute from TDF;
          Complain : Boolean from Standard = Standard_True)
    returns Boolean;
    	---Purpose: Search   in <DF> the  attribute  identified by its 
    	--          <ID> and its <entry>.  returns <True> if found. In
    	--          that case A is setted. 


    ReturnLabel(theCommands : in out Interpretor from Draw; L : Label from TDF)
    returns Interpretor from Draw;
    	---C++: return &

    -- ----------------------------------------------------------------------
    -- Commands
    -- ----------------------------------------------------------------------

    AllCommands   (theCommands : in out Interpretor from Draw);    


    BasicCommands (theCommands : in out Interpretor from Draw);    
    	---Purpose : Basic commands.

    DataCommands (theCommands : in out Interpretor from Draw);    
    	---Purpose : Data framework commands 
    	--           create, clear & copy.

    TransactionCommands (theCommands : in out Interpretor from Draw);    
    	---Purpose : open commit abort a transaction
    	--           undo facilities.

    BrowserCommands (theCommands : in out Interpretor from Draw);    
    	---Purpose : Browser commands .

end DDF;



