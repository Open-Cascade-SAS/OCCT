-- File:	RWStepShape_RWDimensionalLocation.cdl
-- Created:	Tue Apr 18 16:42:58 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0
-- Copyright:	Matra Datavision 1999

class RWDimensionalLocation from RWStepShape

    ---Purpose: Read & Write tool for DimensionalLocation

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    DimensionalLocation from StepShape

is
    Create returns RWDimensionalLocation from RWStepShape;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : DimensionalLocation from StepShape);
	---Purpose: Reads DimensionalLocation

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: DimensionalLocation from StepShape);
	---Purpose: Writes DimensionalLocation

    Share (me; ent : DimensionalLocation from StepShape;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWDimensionalLocation;
