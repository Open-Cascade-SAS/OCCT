-- Created on: 2000-05-10
-- Created by: Andrey BETENEV
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1

class ExternalIdentificationItem from StepAP214
inherits SelectType from StepData

    ---Purpose: Representation of STEP SELECT type ExternalIdentificationItem

uses
    DocumentFile from StepBasic,
    ExternallyDefinedClass from StepAP214,
    ExternallyDefinedGeneralProperty from StepAP214,
    ProductDefinition from StepBasic

is
    Create returns ExternalIdentificationItem from StepAP214;
	---Purpose: Empty constructor

    CaseNum (me; ent: Transient) returns Integer;
	---Purpose: Recognizes a kind of ExternalIdentificationItem select type
	--          1 -> DocumentFile from StepBasic
	--          2 -> ExternallyDefinedClass from StepAP214
	--          3 -> ExternallyDefinedGeneralProperty from StepAP214
	--          4 -> ProductDefinition from StepBasic
	--          0 else

    DocumentFile (me) returns DocumentFile from StepBasic;
	---Purpose: Returns Value as DocumentFile (or Null if another type)

    ExternallyDefinedClass (me) returns ExternallyDefinedClass from StepAP214;
	---Purpose: Returns Value as ExternallyDefinedClass (or Null if another type)

    ExternallyDefinedGeneralProperty (me) returns ExternallyDefinedGeneralProperty from StepAP214;
	---Purpose: Returns Value as ExternallyDefinedGeneralProperty (or Null if another type)

    ProductDefinition (me) returns ProductDefinition from StepBasic;
	---Purpose: Returns Value as ProductDefinition (or Null if another type)

end ExternalIdentificationItem;
