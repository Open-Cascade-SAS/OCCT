-- Created on: 1994-02-03
-- Created by: Jean Marc LACHAUME
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package Geom2dHatch

uses
    Geom2dAdaptor,
    Geom2dInt,
    gp,
    HatchGen,
    TCollection,
    TColStd,
    TopClass,
    TopAbs

is
    
    class Intersector ;
    
    class Hatcher;
    
    class Element;
    class Elements;
    class Hatching;
    
    class Hatchings instantiates DataMap from TCollection
    (Integer          from Standard,
     Hatching         from Geom2dHatch,
     MapIntegerHasher from TColStd) ;

    class Classifier instantiates FaceClassifier from  TopClass 
    (Elements    from Geom2dHatch,
     Curve       from Geom2dAdaptor,
     Intersector from Geom2dHatch);

    private class MapOfElements instantiates DataMap from TCollection
    (Integer          from Standard,
     Element          from Geom2dHatch,
     MapIntegerHasher from TColStd);

end Geom2dHatch ;
