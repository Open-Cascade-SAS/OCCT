-- Created on: 1992-12-02
-- Created by: Isabelle GRIGNON
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class CelGProps  from GProp inherits GProps from GProp

	--- Purpose  : 
	--  Computes the  global properties of bounded curves 
	--  in 3D space. 
	--  It can be an elementary curve from package gp such as 
	--  Lin, Circ, Elips, Parab .

uses  Circ  from gp,
      Lin   from gp,
      Parab from gp,
      Pnt   from gp
       
is

    Create returns CelGProps;
  
    Create (C : Circ from gp; CLocation : Pnt)   returns CelGProps;

    Create (C : Circ from gp; U1, U2 : Real; CLocation : Pnt)returns CelGProps;

    Create (C : Lin from gp; U1, U2 : Real; CLocation : Pnt) returns CelGProps;

    SetLocation(me : in out;CLocation : Pnt) ;

    Perform(me : in out; C :Circ; U1,U2 : Real);
    
    Perform(me : in out; C : Lin ; U1,U2 : Real);

end CelGProps;


