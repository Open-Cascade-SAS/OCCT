-- Created on: 1991-02-06
-- Created by: Arnaud BOUZY
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class RUIterator from Expr

	---Purpose: Iterates on NamedUnknowns in a GeneralRelation. 
    	---Level : Internal

uses GeneralRelation from Expr,
    NamedUnknown from Expr,
    MapOfNamedUnknown from Expr
    
raises NoMoreObject from Standard,
    NoSuchObject from Standard

is

    Create(rel : GeneralRelation)
    ---Purpose: Creates an iterator on every NamedUnknown contained in 
    --          <rel>.
    returns RUIterator;
    
    More(me)
    ---Purpose: Returns False if on other unknown remains.
    returns Boolean
    is static;
    
    Next(me : in out)
    raises NoMoreObject
    is static;
    
    Value(me)
    ---Purpose: Returns current NamedUnknown.
    --          Raises exception if no more unknowns remain.
    returns NamedUnknown
    raises NoSuchObject
    is static;

fields

    myMap : MapOfNamedUnknown;
    myCurrent : Integer;

end RUIterator;
