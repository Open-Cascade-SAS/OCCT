-- Created on: 1995-02-01
-- Created by: Marie Jose MARTZ
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Geom2dVector from Geom2dToIGES inherits Geom2dEntity from Geom2dToIGES

    ---Purpose: This class implements the transfer of the Vector from Geom2d
    --          to IGES . These can be :
    --          . Vector
    --              * Direction
    --              * VectorWithMagnitude
  
uses
 
    Vector               from Geom2d,
    VectorWithMagnitude  from Geom2d,
    Direction            from Geom2d,
    Direction            from IGESGeom,
    Geom2dEntity         from Geom2dToIGES

     
is 
    
    Create returns Geom2dVector from Geom2dToIGES;


    Create(G2dE : Geom2dEntity from Geom2dToIGES)  
    	 returns Geom2dVector from Geom2dToIGES;
    ---Purpose : Creates a tool Geom2dVector ready to run and sets its
    --         fields as G2dE's.

    Transfer2dVector   (me    : in out;
                        start : Vector from Geom2d)
    	 returns mutable Direction from IGESGeom;
    ---Purpose :  Transfert  a  GeometryEntity which  answer True  to  the
    --            member : BRepToIGES::IsGeomVector(Geometry).  If this
    --            Entity could not be converted, this member returns a NullEntity.


    Transfer2dVector   (me    : in out;
                        start : VectorWithMagnitude from Geom2d)
    	 returns mutable Direction from IGESGeom;


    Transfer2dVector   (me    : in out;
                        start : Direction from Geom2d)
    	 returns mutable Direction from IGESGeom;


end Geom2dVector;


