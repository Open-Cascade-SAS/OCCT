-- Created on: 1993-01-07
-- Created by: Christian CAILLET
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



deferred class SelectInList  from IFSelect  inherits SelectAnyList

    ---Purpose : A SelectInList kind Selection selects a List of an Entity,
    --           which is composed of single Entities
    --           To know the list on which to work, SelectInList has two
    --           deferred methods : NbItems (inherited from SelectAnyList) and
    --           ListedEntity (which gives an item as an Entity) which must be
    --           defined to get a List in an Entity of the required Type (and
    --           consider that list is empty if Entity has not required Type)
    --           
    --           As for SelectAnyList, if a type of Entity defines several
    --           lists, a given sub-class of SelectInList is attached on one

uses AsciiString from TCollection, Transient, EntityIterator, Graph, IntParam

raises OutOfRange

is

--    NbItems (me; ent : Transient) returns Integer  is deferred;
--    KeepInputEntity (me; iter : in out EntityIterator) is deferred; 
--    these method are inherited as deferred and remain to be defined

    ListedEntity (me; num : Integer; ent : Transient)
    	returns Transient  raises OutOfRange  is deferred;
    ---Purpose : Returns an Entity, given its rank in the list

    FillResult (me; n1,n2 : Integer; ent : Transient;
    	result : in out EntityIterator);
    ---Purpose : Puts into the result, the sub-entities of the list, from n1 to
    --           n2 included. Remark that adequation with Entity's type and
    --           length of list has already been made at this stage
    --           Called by RootResult; calls ListedEntity (see below)

end SelectInList;
