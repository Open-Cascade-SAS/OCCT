-- File:        ColourSpecification.cdl
-- Created:     Fri Dec  1 11:11:16 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class ColourSpecification from StepVisual 

inherits Colour from StepVisual 

uses

	HAsciiString from TCollection
is

	Create returns mutable ColourSpecification;
	---Purpose: Returns a ColourSpecification

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection) is virtual;

	-- Specific Methods for Field Data Access --

	SetName(me : mutable; aName : mutable HAsciiString);
	Name (me) returns mutable HAsciiString;

fields

	name : HAsciiString from TCollection;

end ColourSpecification;
