-- File:	StepFEA_FeaRepresentationItem.cdl
-- Created:	Thu Dec 12 17:51:06 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class FeaRepresentationItem from StepFEA
inherits RepresentationItem from StepRepr

    ---Purpose: Representation of STEP entity FeaRepresentationItem

uses
    HAsciiString from TCollection

is
    Create returns FeaRepresentationItem from StepFEA;
	---Purpose: Empty constructor

end FeaRepresentationItem;
