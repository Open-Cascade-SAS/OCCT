-- File:        CurveReplica.cdl
-- Created:     Fri Dec  1 11:11:17 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class CurveReplica from StepGeom 

inherits Curve from StepGeom 

uses

	CartesianTransformationOperator from StepGeom, 
	HAsciiString from TCollection
is

	Create returns mutable CurveReplica;
	---Purpose: Returns a CurveReplica


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aParentCurve : mutable Curve from StepGeom;
	      aTransformation : mutable CartesianTransformationOperator from StepGeom) is virtual;

	-- Specific Methods for Field Data Access --

	SetParentCurve(me : mutable; aParentCurve : mutable Curve);
	ParentCurve (me) returns mutable Curve;
	SetTransformation(me : mutable; aTransformation : mutable CartesianTransformationOperator);
	Transformation (me) returns mutable CartesianTransformationOperator;

fields

	parentCurve : Curve from StepGeom;
	transformation : CartesianTransformationOperator from StepGeom;

end CurveReplica;
