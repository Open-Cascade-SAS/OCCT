-- Created on: 1995-12-04
-- Created by: Laurent BOURESCHE
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class TgtOnCoons from GeomFill inherits TgtField from GeomFill

	---Purpose: Defines   an   algorithmic  tangents  field   on a
	--          boundary of a CoonsAlgPatch.

uses
    Vec           from gp,
    BSpline       from Law,
    CoonsAlgPatch from GeomFill

is
    Create(K : CoonsAlgPatch from GeomFill;
           I : Integer from Standard)
    returns mutable TgtOnCoons from GeomFill;

    Value(me; W : Real from Standard)
    returns Vec from gp;
    ---Purpose: Computes  the value  of the    field of tangency    at
    --          parameter W.

    D1(me; W : Real from Standard)
    returns Vec from gp;
    ---Purpose: Computes the  derivative of  the field of  tangency at
    --          parameter W.

    D1(me; W : Real from Standard; T, DT : out Vec from gp);
    ---Purpose: Computes the value and the  derivative of the field of
    --          tangency at parameter W.

fields

    myK    : CoonsAlgPatch from GeomFill;
    ibound : Integer from Standard;

end TgtOnCoons;
