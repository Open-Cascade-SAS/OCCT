-- File:        UniformCurveAndRationalBSplineCurve.cdl
-- Created:     Mon Dec  4 12:02:33 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWUniformCurveAndRationalBSplineCurve from RWStepGeom

	---Purpose : Read & Write Module for UniformCurveAndRationalBSplineCurve

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     UniformCurveAndRationalBSplineCurve from StepGeom,
     EntityIterator from Interface

is

	Create returns RWUniformCurveAndRationalBSplineCurve;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable UniformCurveAndRationalBSplineCurve from StepGeom);

	WriteStep (me; SW : in out StepWriter; ent : UniformCurveAndRationalBSplineCurve from StepGeom);

	Share(me; ent : UniformCurveAndRationalBSplineCurve from StepGeom; iter : in out EntityIterator);

end RWUniformCurveAndRationalBSplineCurve;
