-- Created on: 1997-01-10
-- Created by: Christophe MARION
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PolyInternalNode from HLRAlgo inherits TShared from MMgt

uses
    Address from Standard,
    Integer from Standard
    
is
    Create returns mutable PolyInternalNode from HLRAlgo; 
    	---C++: inline
    
    Indices(me) returns Address from Standard
    	---C++: inline
    is static;

    RValues(me) returns Address from Standard
    	---C++: inline
    is static;

fields
    myIndices : Integer from Standard[4];
    myRValues : Real    from Standard[11];
    
end PolyInternalNode;
