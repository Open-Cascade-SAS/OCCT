-- Created on: 1993-03-03
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Update:      fma


package PTopLoc 

	---Purpose: The  PTopLoc     package      describes persistent
	--          structures for 3D local coordinate systems.
	--          
	--          The  class Datum3D describes  an  elementary local
	--          coordinate system.   It is a linear transformation
	--          (Trsf  from  gp).   The  transformation  is  rigid
	--          (Rotation +  Translation).
	--          
	--          The private    class  ItemLocation represents   an
	--          elementary  local   coordinate   system  (Datum3D)
	--          raised to  an Integer power  elevation. It is used
	--          to link coordinate systems in a Location.
	--          
	--          The  class Location  describes a local  coordinate
	--          system.   It   is  a  chain   of  elementary local
	--          coordinate systems raised to power elevations. The
	--          Location keeps track  of how the coordinate system
	--          was built.

uses

    Standard,
    gp

is
    class Datum3D;
    -- inherits Persistent from Standard
	---Purpose: Persistent elementary local coordinate system.
	
    private class ItemLocation;
    -- inherits Persistent from Standard
	---Purpose: Persistent class  used to  implement Locations.
	
    class Location;
    -- inherits Storable from Standard
	---Purpose: Storable composite local coordinate system.

end PTopLoc;
