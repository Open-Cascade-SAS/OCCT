-- Created on: 1993-03-02
-- Created by: Philippe DAUTRY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Plane from PGeom inherits ElementarySurface from PGeom

        ---Purpose : This class describes the infinite plane.
        --         
	---See Also : Plane from Geom.


uses Ax3      from gp

is


  Create returns mutable Plane from PGeom;
	---Purpose: Create a plane with default values.
    	---Level: Internal 


  Create (aPosition : Ax3 from gp)
    	returns mutable Plane from PGeom;
	---Purpose: Creates a Plane with these field values.
    	---Level: Internal 


end;

