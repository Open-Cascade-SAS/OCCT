-- Created on: 1992-09-23
-- Created by: Christian CAILLET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Articulations  from IFGraph  inherits GraphContent

    	---Purpose : this class gives entities which are Articulation points
    	--           in a whole Model or in a sub-part
    	--           An Articulation Point divides the graph in two (or more)
    	--           disconnected sub-graphs
    	--           Identifying Articulation Points allows improving
    	--           efficiency of spliting a set of Entities into sub-sets

uses Transient, HSequenceOfInteger, EntityIterator, Graph

is

    Create (agraph : Graph; whole : Boolean) returns Articulations;
    ---Purpose : creates Articulations to evaluate a Graph
    --           whole True : works on the whole Model
    --           whole False : remains empty, ready to work on a sub-part

    GetFromEntity (me : in out; ent : any Transient);
    ---Purpose : adds an entity and its shared ones to the list

    GetFromIter (me : in out; iter : EntityIterator);
    ---Purpose : adds a list of entities (as an iterator)

    ResetData (me : in out);
    ---Purpose : Allows to restart on a new data set

    	-- --   Results   -- --
    	--   More-Next-Value give Articulation points

    Evaluate (me : in out) is redefined;
    ---Purpose : Evaluates the list of Articulation points

    Visit (me : in out; num : Integer) returns Integer  is private;
    ---Purpose : basic routine of computation
    --           (see book Sedgewick "Algorithms", p 392)

fields

    thegraph : Graph;
    thenow   : Integer;  -- for Visit algorithm
    thelist  : HSequenceOfInteger;  -- results from Visiting

end Articulations;
