-- Created on: 1993-04-07
-- Created by: Laurent BUCHARD
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class IntersectionSegment from IntCurveSurface
 

    ---Purpose: A IntersectionSegment describes a segment of curve 
    --          (w1,w2) where distance(C(w),Surface) is less than a  
    --          given tolerances. 
    
    ---Level: Public

uses

    IntersectionPoint    from IntCurveSurface

is

    Create
    	returns IntersectionSegment from IntCurveSurface;
	
    Create(P1: IntersectionPoint from IntCurveSurface;
    	   P2: IntersectionPoint from IntCurveSurface)
	returns IntersectionSegment from IntCurveSurface;
	
    SetValues(me: in out;
    	     P1: IntersectionPoint from IntCurveSurface;
	     P2: IntersectionPoint from IntCurveSurface)
	 is static;
	 
    Values(me;
    	  P1: out IntersectionPoint from IntCurveSurface;
	  P2: out IntersectionPoint from IntCurveSurface)
	 is static;
	 
    FirstPoint(me;
	       P1: out IntersectionPoint from IntCurveSurface)
	 is static;	 

    SecondPoint(me;
	        P2: out IntersectionPoint from IntCurveSurface)
	 is static;

	 
    FirstPoint(me)
	returns IntersectionPoint from IntCurveSurface 
	---C++: return const &
        is static;	 

    SecondPoint(me)
    	 returns IntersectionPoint from IntCurveSurface
	 ---C++: return const &
	 is static;
 
    Dump(me)
          is static;

fields

    myP1 : IntersectionPoint from IntCurveSurface;
    myP2 : IntersectionPoint from IntCurveSurface;
 
end IntersectionSegment;

