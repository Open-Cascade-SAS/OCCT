-- Created on: 1996-04-10
-- Created by: Joelle CHAUVET
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Modified:	Mon Dec  9 10:30:56 1996
--    by:	Joelle CHAUVET
--		G1135 : Empty constructor


class Network from AdvApp2Var

uses

    Boolean,Integer,Real from Standard,
    SequenceOfReal,HArray1OfReal from TColStd,
    IsoType from GeomAbs,
    Patch, SequenceOfPatch, Framework from AdvApp2Var

raises NoSuchObject from Standard 

is
    Create returns Network;
    Create(Net : SequenceOfPatch; TheU,TheV : SequenceOfReal) returns Network;
    FirstNotApprox(me; Index :  out Integer)
    ---Purpose: search the Index of the first Patch not approximated,
    --          if all Patches are approximated Standard_False is returned
    returns Boolean; 
    ChangePatch(me: in out; Index : Integer) 
    ---C++: alias operator()
    ---C++: return &
    ---C++: inline
    returns Patch;
    UpdateInU(me: in out; CuttingValue : Real);
    UpdateInV(me: in out; CuttingValue : Real);
    SameDegree(me : in out; iu, iv : Integer; ncfu, ncfv : out Integer);
    NbPatch(me) returns Integer;
    NbPatchInU(me) returns Integer;
    NbPatchInV(me) returns Integer;
    UParameter(me; Index : Integer) returns Real;
    VParameter(me; Index : Integer) returns Real;
    Patch(me; UIndex, VIndex : Integer) 
    ---C++: alias operator()
    ---C++: return const &
    ---C++: inline
    returns Patch;
    

fields

    myNet         : SequenceOfPatch;
    myUParameters : SequenceOfReal;
    myVParameters : SequenceOfReal;

end Network;

