-- Created on: 1993-03-23
-- Created by: BBL
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Modified:	02-06-98 : FMN ; Suppression appel Clear (deja fait dans ALienData)

class SGIRGBAlienImage from AlienImage inherits AlienUserImage from AlienImage

    	---Purpose: Defines an SGI .rgb Alien image, i.e. an image using
    	-- the image format for Silicon Graphics workstations.

uses
	File 			from OSD,
	AsciiString 		from TCollection,
	ColorImage 		from Image,
	PseudoColorImage 	from Image,
	Image			from Image,
	SGIRGBAlienData 	from AlienImage

is
	Create returns mutable SGIRGBAlienImage from AlienImage;
    	---Purpose: Constructs an empty SGI .rgb Alien image.
    
	Clear( me : in out mutable) ;
	---Level: Public
	---Purpose: Frees memory allocated by SGIRGBAlienImage

	SetName( me : in out mutable;
		 aName : in AsciiString from TCollection) ;
	---Level: Public
	---Purpose: Set Image name .

	Name( me : in immutable ) returns AsciiString from TCollection ;
		  ---C++: return const &
    		  ---Purpose: Reads the  Image name .

	ToImage( me : in immutable ) 
	  returns mutable Image from Image ;
	---Level: Public
	---Purpose : Converts a SGIRGBAlienImage object to a Image object.

	FromImage( me : in out mutable ; anImage : in Image from Image ) ;
	---Level: Public
	---Purpose : Converts a Image object to a SGIRGBAlienImage object.

	Read ( me : in out mutable; afile : in out File from OSD )
	  returns Boolean from Standard ;
	---Purpose: Reads content of a SGIRGBAlienImage object from a file
	--          Returns True if file is a XWD file .

	Write( me : in immutable; afile : in out File from OSD )
	  returns Boolean from Standard ;
	---Purpose: Writes content of a SGIRGBAlienImage object to a file

fields
	myData : SGIRGBAlienData  from  AlienImage;

end ;
 
