-- Created on: 1997-03-26
-- Created by: Christian CAILLET
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DerivedUnitElement  from StepBasic    inherits TShared

    ---Purpose : Added from StepBasic Rev2 to Rev4

uses
     NamedUnit from StepBasic

is

    Create returns DerivedUnitElement;

    Init (me : mutable; aUnit : NamedUnit from StepBasic; aExponent : Real);

    SetUnit (me : mutable; aUnit : NamedUnit from StepBasic);
    Unit (me) returns NamedUnit from StepBasic;

    SetExponent (me : mutable; aExponent : Real);
    Exponent (me) returns Real;

fields

    theUnit : NamedUnit from StepBasic;
    theExponent : Real;

end DerivedUnitElement;
