-- Created on: 1994-08-30
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Modification from Draft inherits Modification from BRepTools

	---Purpose: 

uses Shape       from TopoDS,
     Face        from TopoDS,
     Edge        from TopoDS,
     Vertex      from TopoDS,
     Location    from TopLoc,
     ListOfShape                      from TopTools,
     IndexedDataMapOfShapeListOfShape from TopTools,
     
     Orientation from TopAbs,
     Shape       from GeomAbs,

     Surface  from Geom,
     Curve    from Geom,
     Curve    from Geom2d,
     
     Pnt      from gp,
     Lin      from gp,
     Pln      from gp,
     Dir      from gp,
     
     ErrorStatus               from Draft,
     DataMapOfFaceFaceInfo     from Draft,
     DataMapOfEdgeEdgeInfo     from Draft,
     DataMapOfVertexVertexInfo from Draft


raises NotDone           from StdFail,
       NoSuchObject      from Standard,
       ConstructionError from Standard

is

    Create(S: Shape from TopoDS)
    
    	returns mutable Modification from Draft;


    Clear(me: mutable)
	---Purpose: Resets on the same shape.
        is static;
    

    Init(me: mutable; S: Shape from TopoDS)
	---Purpose: Changes the basis shape and resets.
    is static;


    Add(me: mutable; F           : Face    from TopoDS; 
                     Direction   : Dir     from gp;
                     Angle       : Real    from Standard; 
		     NeutralPlane: Pln     from gp; 
                     Flag        : Boolean from Standard = Standard_True)
	---Purpose: Adds  the  face  F    and propagates    the  draft
	--          modification to  its  neighbour faces if they  are
	--          tangent. If an error occurs, will return False and
	--          ProblematicShape  will  return the "bad" face.

    	returns Boolean from Standard
        raises ConstructionError from Standard
	       -- The exception is raised if ProblematicShape does not
	       -- return a null shape
    	is static;


    Remove(me: mutable; F: Face from TopoDS)
	---Purpose: Removes the face F and the neighbour faces if they
	--          are tangent.   It will be  necessary to  call this
	--          method if  the  method Add returns Standard_False,
	--          to unset ProblematicFace.


    	raises NoSuchObject from Standard
	       -- The exception is raised if F has not been added.
    	is static;



    Perform(me: mutable)
	---Purpose: Performs the draft angle modification and sets the
	--          value returned by the method  IsDone.  If an error
	--          occurs, IsDone  will return Standard_False, and an
	--          error status will  be  given by the  method Error,
	--          and the  shape on which  the problem appeared will
	--          be given by ProblematicShape

	raises ConstructionError from Standard
	--- The exception   is  raised  if  ProblematicShape  does not
	--  return a null shape.
    	is static;


    IsDone(me)
	---Purpose: Returns  True  if   Perform has  been  succesfully
	--          called. Otherwise more information can be obtained
	--          using the methods Error() and ProblematicShape().
    	returns Boolean from Standard
	is static;


    Error(me)
    
    	returns ErrorStatus from Draft
	is static;


    ProblematicShape(me)
	---Purpose: Returns the shape (Face,  Edge or Vertex) on which
	--          an error occured.
    
    	returns Shape from TopoDS
	---C++: return const&
	is static;


    ConnectedFaces(me: mutable; F: Face from TopoDS)
    
    	returns ListOfShape from TopTools
	---Purpose: Returns all  the  faces   which  have been   added
	--          together with the face <F>.
	--          
	---C++: return const&

    	raises NoSuchObject from Standard,
	       -- The exception is raised if F has not been added.
               NotDone from StdFail
	       -- The exception is raised if IsDone returns False.
	is static;


    ModifiedFaces(me: mutable)
    
    	returns ListOfShape from TopTools
	---Purpose: Returns all the faces  on which a modification has
	--          been given.
	--          
	---C++: return const&

    	raises NotDone from StdFail
	-- The exception is raised if ProblematicShape does not return
	-- a null shape.
	is static;




-- Methods inherited from BRepTools_Modification

    NewSurface(me: mutable; F       :     Face     from TopoDS;
                            S       : out Surface  from Geom;
		            L       : out Location from TopLoc;
		            Tol     : out Real     from Standard;
                            RevWires : out Boolean from Standard;
                            RevFace  : out Boolean from Standard)



      	---Purpose: Returns Standard_True if   the face <F>  has  been
      	--          modified.  In this case,  <S> is the new geometric
      	--          support of the  face,  <L> the new  location,<Tol>
      	--          the   new tolerance.<RevWires>  has  to  be set to
      	--          Standard_True when   the modification reverses the
      	--          normal   of  the  surface.(the  wires   have to be
      	--          reversed).  <RevFace>    has    to  be   set    to
      	--          Standard_True  if  the orientation of the modified
      	--          face changes in  the shells which contain it. Here
      	--          it will be set to Standard_False.
      	--          
      	--          Otherwise, returns Standard_False, and <S>,   <L>,
      	--          <Tol> , <RevWires> ,<RevFace> are not  significant.
    
    	returns Boolean from Standard
	;
	

    NewCurve(me: mutable; E  :     Edge     from TopoDS;
                          C  : out Curve from Geom;
		          L  : out Location from TopLoc;
		          Tol: out Real     from Standard)
    
    	returns Boolean from Standard
	;
	
	---Purpose: Returns Standard_True  if  the edge  <E> has  been
	--          modified.  In this case,  <C> is the new geometric
	--          support of the  edge, <L> the  new location, <Tol>
	--          the         new    tolerance.   Otherwise, returns
	--          Standard_False,    and  <C>,  <L>,   <Tol> are not
	--          significant.
    

    NewPoint(me: mutable; V  :     Vertex from TopoDS;
                          P  : out Pnt    from gp;
		          Tol: out Real   from Standard)
    
    	returns Boolean from Standard
	;
	
	---Purpose: Returns  Standard_True if the  vertex <V> has been
	--          modified.  In this  case, <P> is the new geometric
	--          support of the vertex,   <Tol> the new  tolerance.
	--          Otherwise, returns Standard_False, and <P>,  <Tol>
	--          are not significant.
    

    NewCurve2d(me: mutable;  E    :     Edge  from TopoDS;
                             F    :     Face  from TopoDS;
                             NewE :     Edge     from TopoDS;
                             NewF :     Face     from TopoDS;
                             C    : out Curve from Geom2d;
		             Tol  : out Real  from Standard)
    
    	returns Boolean from Standard
	;
	
	---Purpose: Returns Standard_True if  the edge  <E> has a  new
	--          curve on surface on the face <F>.In this case, <C>
	--          is the new geometric support of  the edge, <L> the
	--          new location, <Tol> the new tolerance.
	--          
	--          Otherwise, returns  Standard_False, and <C>,  <L>,
	--          <Tol> are not significant.
	--          
	--          <NewE> is the new  edge created from  <E>.  <NewF>
	--          is the new face created from <F>. They may be usefull.


    NewParameter(me: mutable; V  :     Vertex from TopoDS;
                              E  :     Edge   from TopoDS;
                              P  : out Real   from Standard;
  		              Tol: out Real   from Standard)
    
    	returns Boolean from Standard
	;
	
	---Purpose: Returns Standard_True if the Vertex  <V> has a new
	--          parameter on the  edge <E>. In  this case,  <P> is
	--          the parameter,    <Tol>  the     new    tolerance.
	--          Otherwise, returns Standard_False, and <P>,  <Tol>
	--          are not significant.

    

    Continuity(me: mutable; E          : Edge from TopoDS;
    	                    F1,F2      : Face from TopoDS;
			    NewE       : Edge from TopoDS;
			    NewF1,NewF2: Face from TopoDS)
    
    	returns Shape from GeomAbs;
	
	---Purpose: Returns the  continuity of  <NewE> between <NewF1>
	--          and <NewF2>.
	--          
	--          <NewE> is the new  edge created from <E>.  <NewF1>
	--          (resp. <NewF2>) is the new  face created from <F1>
	--          (resp. <F2>).


-- Private implementation methods

    InternalAdd(me: mutable; F           : Face    from TopoDS; 
                             Direction   : Dir     from gp;
                             Angle       : Real    from Standard; 
		             NeutralPlane: Pln     from gp; 
    	    	    	     Flag        : Boolean from Standard = Standard_True)

	returns Boolean from Standard	     
    	is static private;
			     
			     
    Propagate(me: mutable)
    
	returns Boolean from Standard	     
    	is static private;
    
    
    NewCurve(me: mutable; C           : Curve       from Geom;
                          S           : Surface     from Geom;
                          OriS        : Orientation from TopAbs;
                          Direction   : Dir         from gp;
                          Angle       : Real        from Standard; 
			  NeutralPlane: Pln         from gp; 
                          Flag        : Boolean     from Standard = Standard_True)

	returns mutable Curve from Geom
	is static private;


    NewSurface(me: mutable; S           : Surface     from Geom;
                            OriS        : Orientation from TopAbs;
                            Direction   : Dir         from gp;
                            Angle       : Real        from Standard; 
			    NeutralPlane: Pln         from gp)

	returns mutable Surface from Geom
	is static private;


fields

    myFMap  : DataMapOfFaceFaceInfo     from Draft;
    myEMap  : DataMapOfEdgeEdgeInfo     from Draft;
    myVMap  : DataMapOfVertexVertexInfo from Draft;
    myComp  : Boolean                   from Standard;
    myShape : Shape                     from TopoDS;
    badShape: Shape                     from TopoDS;
    errStat : ErrorStatus               from Draft;
    curFace : Face                      from TopoDS;
    conneF  : ListOfShape               from TopTools;
    myEFMap : IndexedDataMapOfShapeListOfShape from TopTools;
    
end Modification;
