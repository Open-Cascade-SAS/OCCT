-- Created on: 1994-05-31
-- Created by: Christian CAILLET
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SelectLevelNumber  from IGESSelect  inherits SelectExtract

    ---Purpose : This selection looks at Level Number of IGES Entities :
    --           it considers items attached, either to a single level with a
    --           given value, or to a level list which contains this value
    --           
    --           Level = 0  means entities not attached to any level
    --           
    --           Remark : the class CounterOfLevelNumber gives informations
    --             about present levels in a file.

uses AsciiString from TCollection, Transient, InterfaceModel, IntParam

is

    Create returns SelectLevelNumber;
    ---Purpose : Creates a SelectLevelNumber, with no Level criterium : see
    --           SetLevelNumber. Empty, this selection filters nothing.

    SetLevelNumber (me : mutable; levnum : IntParam);
    ---Purpose : Sets a Parameter as Level criterium

    LevelNumber (me) returns IntParam;
    ---Purpose : Returns the Level criterium. NullHandle if not yet set
    --           (interpreted as Level = 0 : no level number attached)

    Sort (me; rank : Integer; ent : Transient; model : InterfaceModel)
    	returns Boolean;
    ---Purpose : Returns True if <ent> is an IGES Entity with Level Number
    --           admits the criterium (= value if single level, or one of the
    --           attached level numbers = value if level list)

    ExtractLabel (me) returns AsciiString from TCollection;
    ---Purpose : Returns the Selection criterium :
    --           "IGES Entity, Level Number admits <nn>" (if nn > 0) or
    --           "IGES Entity attached to no Level" (if nn = 0)

fields

    thelevnum : IntParam;

end SelectLevelNumber;
