-- Created on: 2002-04-09
-- Created by: QA Admin
-- Copyright (c) 2002-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class PresentableObject from QARoutelous inherits InteractiveObject from AIS
uses
    Selection from SelectMgr,
    PresentationManager3d from PrsMgr,
    Presentation from Prs3d,
    TypeOfPresentation3d from PrsMgr
is
    
    Create(aTypeOfPresentation3d: TypeOfPresentation3d from PrsMgr = PrsMgr_TOP_AllView) returns mutable PresentableObject from QARoutelous;
    
    ComputeSelection(me:mutable; aSelection :mutable Selection from SelectMgr;
                                 aMode      : Integer) is redefined virtual protected;

    Compute(me:mutable;
    	    aPresentationManager: PresentationManager3d from PrsMgr;
            aPresentation: mutable Presentation from Prs3d;
            aMode: Integer from Standard = 0)
    is redefined virtual protected;
	    
end PresentableObject;
    
