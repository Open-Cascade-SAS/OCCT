-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class BSplineCurveWithKnots from StepGeom 

inherits BSplineCurve from StepGeom 

uses

	HArray1OfInteger from TColStd, 
	HArray1OfReal from TColStd, 
	KnotType from StepGeom, 
	Integer from Standard, 
	Real from Standard, 
	HAsciiString from TCollection, 
	HArray1OfCartesianPoint from StepGeom, 
	BSplineCurveForm from StepGeom, 
	Logical from StepData
is

	Create returns mutable BSplineCurveWithKnots;
	---Purpose: Returns a BSplineCurveWithKnots


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aDegree : Integer from Standard;
	      aControlPointsList : mutable HArray1OfCartesianPoint from StepGeom;
	      aCurveForm : BSplineCurveForm from StepGeom;
	      aClosedCurve : Logical from StepData;
	      aSelfIntersect : Logical from StepData) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aDegree : Integer from Standard;
	      aControlPointsList : mutable HArray1OfCartesianPoint from StepGeom;
	      aCurveForm : BSplineCurveForm from StepGeom;
	      aClosedCurve : Logical from StepData;
	      aSelfIntersect : Logical from StepData;
	      aKnotMultiplicities : mutable HArray1OfInteger from TColStd;
	      aKnots : mutable HArray1OfReal from TColStd;
	      aKnotSpec : KnotType from StepGeom) is virtual;

	-- Specific Methods for Field Data Access --

	SetKnotMultiplicities(me : mutable; aKnotMultiplicities : mutable HArray1OfInteger);
	KnotMultiplicities (me) returns mutable HArray1OfInteger;
	KnotMultiplicitiesValue (me; num : Integer) returns Integer;
	NbKnotMultiplicities (me) returns Integer;
	SetKnots(me : mutable; aKnots : mutable HArray1OfReal);
	Knots (me) returns mutable HArray1OfReal;
	KnotsValue (me; num : Integer) returns Real;
	NbKnots (me) returns Integer;
	SetKnotSpec(me : mutable; aKnotSpec : KnotType);
	KnotSpec (me) returns KnotType;

fields

	knotMultiplicities : HArray1OfInteger from TColStd;
	knots : HArray1OfReal from TColStd;
	knotSpec : KnotType from StepGeom; -- an Enumeration

end BSplineCurveWithKnots;
