-- Created on: 1996-02-13
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class GTool from TopOpeBRepBuild

uses

    GTopo from TopOpeBRepBuild,
    ShapeEnum from TopAbs,
    OStream from Standard
    
is

    GFusUnsh(myclass; s1,s2 : ShapeEnum from TopAbs) returns GTopo;
    GFusSame(myclass; s1,s2 : ShapeEnum from TopAbs) returns GTopo;
    GFusDiff(myclass; s1,s2 : ShapeEnum from TopAbs) returns GTopo;

    GCutUnsh(myclass; s1,s2 : ShapeEnum from TopAbs) returns GTopo;
    GCutSame(myclass; s1,s2 : ShapeEnum from TopAbs) returns GTopo;
    GCutDiff(myclass; s1,s2 : ShapeEnum from TopAbs) returns GTopo;

    GComUnsh(myclass; s1,s2 : ShapeEnum from TopAbs) returns GTopo;
    GComSame(myclass; s1,s2 : ShapeEnum from TopAbs) returns GTopo;
    GComDiff(myclass; s1,s2 : ShapeEnum from TopAbs) returns GTopo;

    Dump(myclass; OS : in out OStream from Standard);
    
end GTool;
