-- Created on: 2000-08-15
-- Created by: data exchange team
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Location from PXCAFDoc inherits Attribute from PDF

	---Purpose: 

uses 
--    Location from TopLoc,
    Location from PTopLoc
is
    Create returns mutable Location from PXCAFDoc;
    
    Create (Loc: Location from PTopLoc) returns mutable Location from PXCAFDoc;
    
    Set (me: mutable; Loc: Location from PTopLoc);
    
    Get (me) returns Location from PTopLoc;
    
fields
    myPLocation : Location from PTopLoc;
    
end Location;
