-- Created on: 1993-04-15
-- Created by: Gilles DEBARBOUILLE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Color from Materials

	---Purpose: This class  encapsulates   a Quantity_Color  in  a
	--          Transient object, to be used in an ObjectProperty
	--          from the package Dynamic.

inherits

    Transient
    
uses

    Color from Quantity, TypeOfColor from Quantity, NameOfColor from Quantity

--raises

is

    Create returns mutable Color from Materials;    
    ---Level: Internal     
    ---Purpose: Creates an empty instance of Color.
    
    Create(acolor : Color from Quantity)
    ---Level: Internal     
    ---Purpose: Creates an instance of Color, with <acolor> as color.
    
    returns mutable Color from Materials;
    
    Color(me : mutable ; acolor : Color from Quantity)    
    ---Level: Internal     
    ---Purpose: Sets <acolor> into <me>.    
    is static;

    Color(me) returns Color from Quantity   
    ---Level: Internal     
    ---Purpose: Returns a Quantity_Color corresponding to <me>.    
    is static;

    Color(me; aTypeOfColor : in TypeOfColor from Quantity; Reel1, Reel2, Reel3 : out Real from Standard);
    ---Purpose: Get the values ( RGB or HLS )  between 0.0 and 1.0

    Color255(me; aTypeOfColor : in TypeOfColor from Quantity; Reel1, Reel2, Reel3 : out Real from Standard);
    ---Purpose: Get the values ( RGB or HLS )  between 0.0 and 255.0

    SetColor(me : mutable; aTypeOfColor : in TypeOfColor from Quantity; Reel1, Reel2, Reel3 : in Real from Standard);
    ---Purpose: Set the values ( RGB or HLS )  between 0.0 and 1.0

    SetColor255(me : mutable; aTypeOfColor : in TypeOfColor from Quantity; Reel1, Reel2, Reel3 : in Real from Standard);
   ---Purpose: Set the values ( RGB or HLS )  between 0.0 and 255.0

fields

    thecolor : Color from Quantity;

end Color;
