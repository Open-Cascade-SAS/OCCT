-- Created on: 1993-06-17
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


package TopOpeBRep 

	---Purpose: This package provides  the topological  operations
	--          on the BRep data structure.

uses

    Standard,
    MMgt,
    TColStd,
    TopAbs,
    TopoDS,
    TopTools,
    TopExp,
    gp,
    Geom,
    Geom2d,
    GeomAbs,
    Geom2dAdaptor,
    Bnd,
    BRep,
    BRepClass,
    BRepAdaptor,
    BRepTopAdaptor,
    ProjLib,
    IntRes2d,
    Geom2dInt,    
    
    IntSurf,
    IntPatch,

    GeomAdaptor,
    IntCurveSurface,
    BRepIntCurveSurface,

    TopOpeBRepDS,
    TopOpeBRepTool,
    TCollection
    
is

    enumeration TypeLineCurve is
    	ANALYTIC,RESTRICTION,WALKING,
        LINE,CIRCLE,ELLIPSE,PARABOLA,HYPERBOLA,
	OTHERTYPE
    end TypeLineCurve;

    class VPointInter;

    class Array1OfVPointInter instantiates Array1 from TCollection
    	(VPointInter from TopOpeBRep);

    class HArray1OfVPointInter instantiates HArray1 from TCollection
    	(VPointInter from TopOpeBRep, Array1OfVPointInter from TopOpeBRep);

    pointer PThePointOfIntersection to Point from IntPatch;
    class VPointInterIterator;

    pointer PPntOn2S to PntOn2S from IntSurf;
    class WPointInter;
    
    class WPointInterIterator;
	 
    class LineInter;
    pointer PLineInter to LineInter from TopOpeBRep;
	
    class Array1OfLineInter instantiates Array1 from TCollection
    	(LineInter from TopOpeBRep);

    class HArray1OfLineInter instantiates HArray1 from TCollection
    	(LineInter from TopOpeBRep, Array1OfLineInter from TopOpeBRep);

    class DataMapOfTopolTool instantiates DataMap from TCollection 
    	(Shape          from TopoDS,
     	 TopolTool from BRepTopAdaptor,
     	 ShapeMapHasher from TopTools);

    pointer PIntRes2d_IntersectionPoint to IntersectionPoint from IntRes2d;
    class Hctxff2d;
    class Hctxee2d;

    enumeration P2Dstatus is
    	P2DUNK,P2DINT,P2DSGF,P2DSGL,P2DNEW 
    end P2Dstatus;
    
    class Point2d;
    class SequenceOfPoint2d instantiates Sequence from TCollection(Point2d from TopOpeBRep);
    
    class PointClassifier;

    class VPointInterClassifier;

    class GeomTool;
     
    class FacesIntersector;
    ---Purpose: Describes the intersection of two faces.
    pointer PFacesIntersector to FacesIntersector from TopOpeBRep;
	
    class EdgesIntersector;
    ---Purpose: Describes the intersection of two edges on the same surface
    pointer PEdgesIntersector to EdgesIntersector from TopOpeBRep;

    class FaceEdgeIntersector;
    ---Purpose: Describes the intersection of a face and an edge.
	
    class ShapeScanner;

    class ShapeIntersector;

    class ShapeIntersector2d;

    class PointGeomTool;
    
    class FFTransitionTool;

    class Bipoint;
    class ListOfBipoint instantiates List from TCollection(Bipoint);
    
    class FacesFiller;
    pointer PFacesFiller to FacesFiller from TopOpeBRep;
    class FFDumper;

    class EdgesFiller;

    class FaceEdgeFiller;

    class DSFiller;

    Print(TLC  : TypeLineCurve from TopOpeBRep; OS  : in out OStream) 
    ---C++: return &
    returns OStream;
    ---Purpose: Prints the name  of  <TLC>  as  a String  on the
    --          Stream <S> and returns <S>.

end TopOpeBRep;
