-- Created on: 2002-12-12
-- Created by: data exchange team
-- Copyright (c) 2002-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class Curve3dElementProperty from StepFEA
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity Curve3dElementProperty

uses
    HAsciiString from TCollection,
    HArray1OfCurveElementInterval from StepFEA,
    HArray1OfCurveElementEndOffset from StepFEA,
    HArray1OfCurveElementEndRelease from StepFEA

is
    Create returns Curve3dElementProperty from StepFEA;
	---Purpose: Empty constructor

    Init (me: mutable; aPropertyId: HAsciiString from TCollection;
                       aDescription: HAsciiString from TCollection;
                       aIntervalDefinitions: HArray1OfCurveElementInterval from StepFEA;
                       aEndOffsets: HArray1OfCurveElementEndOffset from StepFEA;
                       aEndReleases: HArray1OfCurveElementEndRelease from StepFEA);
	---Purpose: Initialize all fields (own and inherited)

    PropertyId (me) returns HAsciiString from TCollection;
	---Purpose: Returns field PropertyId
    SetPropertyId (me: mutable; PropertyId: HAsciiString from TCollection);
	---Purpose: Set field PropertyId

    Description (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Description
    SetDescription (me: mutable; Description: HAsciiString from TCollection);
	---Purpose: Set field Description

    IntervalDefinitions (me) returns HArray1OfCurveElementInterval from StepFEA;
	---Purpose: Returns field IntervalDefinitions
    SetIntervalDefinitions (me: mutable; IntervalDefinitions: HArray1OfCurveElementInterval from StepFEA);
	---Purpose: Set field IntervalDefinitions

    EndOffsets (me) returns HArray1OfCurveElementEndOffset from StepFEA;
	---Purpose: Returns field EndOffsets
    SetEndOffsets (me: mutable; EndOffsets: HArray1OfCurveElementEndOffset from StepFEA);
	---Purpose: Set field EndOffsets

    EndReleases (me) returns HArray1OfCurveElementEndRelease from StepFEA;
	---Purpose: Returns field EndReleases
    SetEndReleases (me: mutable; EndReleases: HArray1OfCurveElementEndRelease from StepFEA);
	---Purpose: Set field EndReleases

fields
    thePropertyId: HAsciiString from TCollection;
    theDescription: HAsciiString from TCollection;
    theIntervalDefinitions: HArray1OfCurveElementInterval from StepFEA;
    theEndOffsets: HArray1OfCurveElementEndOffset from StepFEA;
    theEndReleases: HArray1OfCurveElementEndRelease from StepFEA;

end Curve3dElementProperty;
