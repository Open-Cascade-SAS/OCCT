-- Created on: 1997-01-08
-- Created by: Robert COUBLANC
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

--Modified by rob on Jul-28-97		


class ConnectedShape from AIS inherits ConnectedInteractive from AIS

	---Purpose: Constructs a Connected Interactive Object with an
    	-- AIS_Shape presentation as its reference Interactive Object.
    	-- In topological decomposition of the shape, this class
    	-- assigns the same owners to the sensitive primitives
    	-- as those in AIS_Shape. Like AIS_Shape, it allows a
    	-- presentation of hidden parts. These are calculated
    	-- automatically from the shape of its reference entity.

    

uses

    Shape                from TopoDS,
    Projector            from Prs3d,
    Presentation         from Prs3d,
    Selection            from SelectMgr,
    Integer              from Standard,
    Shape                from AIS,
    TypeOfPresentation3d from PrsMgr,
    PresentationManager3d from PrsMgr,
    InteractiveObject    from AIS,
    KindOfInteractive    from AIS,
    Location             from TopLoc,
    Transformation       from Geom
raises
    NotImplemented from Standard

is

    Create (aTypeOfPresentation : TypeOfPresentation3d from PrsMgr 
    	    	    	    	  =PrsMgr_TOP_ProjectorDependant) 
    returns mutable  ConnectedShape  from  AIS;
    	---Purpose: Initializes the type of 3d presentation aTypeOfPresentation
        
    Create (aInteractiveShape   : Shape from AIS;
    	    aTypeOfPresentation : TypeOfPresentation3d from PrsMgr 
    	    	    	    	  =PrsMgr_TOP_ProjectorDependant)  
    returns  mutable  ConnectedShape  from  AIS;
    	---Purpose: Initializes the entity aInteractiveShape and the type of 3d presentation aTypeOfPresentation.

    Create(aConnectedShape     : ConnectedShape from AIS;
     	   aTypeOfPresentation : TypeOfPresentation3d from PrsMgr 
    	    	    	    	=PrsMgr_TOP_ProjectorDependant)  
    returns  mutable  ConnectedShape  from  AIS;
    	---Purpose: Initializes the entity aConnectedShape and the type of 3d presentation aTypeOfPresentation.
    
    ---Category:  Redefined methods...

    Type(me) returns KindOfInteractive from AIS
    is redefined virtual;

    Signature(me) returns Integer from Standard
    is redefined virtual;

    AcceptShapeDecomposition(me) 
    returns Boolean from Standard is redefined;



	   
    Connect(me          : mutable; 
    	    anotherIObj : InteractiveObject from AIS) is redefined ;
	---Purpose:  Establishes the connection between the Connected
    	-- Interactive Object, anotherIobj, and its reference
    	-- entity. If there is already a previous connection with
    	-- an Interactive Object, this connection is removed.

    Connect(me:mutable;
    	    anotherIobj: InteractiveObject from AIS;
	    aLocation : Location from TopLoc) is redefined;
	---Purpose: Establishes the connection between the Connected
    	-- Interactive Object, anotherIobj, and its reference
    	-- entity. If there is already a previous connection with
    	-- an Interactive Object, this connection is removed.
    	-- This syntax also initiates the location of the Connected Interactive Object.


    Compute(me:mutable;
    	        aProjector   :         Projector    from Prs3d;
                aPresentation: mutable Presentation from Prs3d)
    is redefined virtual private;
 
    Compute(me                   : mutable;
    	    aProjector           : Projector from Prs3d;
	    aTrsf                : Transformation from Geom;
	    aPresentation        : mutable Presentation from Prs3d)
    is redefined virtual private;

    ComputeSelection(me:mutable; aSelection :mutable Selection from SelectMgr;
                                 aMode      :        Integer   from Standard)
    is redefined virtual private;
    	---Purpose: Generates sensitive entities by copying 
        -- them from myReferense selection specified by aMode,  
        -- creates and sets an entity owner for this entities and adds 
        -- them to aSelection.
    
    Shape(me:mutable) returns Shape from TopoDS;
        ---C++: return const&
    	---Purpose: Returns the topological shape which is the reference
    	-- for the connected shape. Sets hilight mode to index
    	-- 0. This returns a wireframe presentation.
	

    UpdateShape(me:mutable;WithLocation:Boolean from Standard = Standard_True)
    is static private;
    
    Compute(me:mutable;
    	        aProjector   :         Projector    from Prs3d;
                aPresentation: mutable Presentation from Prs3d;
    	    	aShape       :         Shape from TopoDS)
    is  private;

    
fields
    
    myOwnSh : Shape   from TopoDS; -- used for HLR and selection...
    
end ConnectedShape;
