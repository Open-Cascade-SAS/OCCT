-- Created on: 1994-03-30
-- Created by: Laurent BUCHARD
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

generic class SolidClassifier from TopClass
    (TheSolidExplorer    as any;
     TheIntersection3d   as any)
     
     ---Purpose: Provides an algorithm to classify a point in a solid.



uses 
    Pnt     from gp,
    Face    from TopoDS,
    Shape   from TopoDS,
    State   from TopAbs

raises
    DomainError from Standard
    
    
    
is 
       
    Create 
    	---Purpose: Empty constructor.
    returns SolidClassifier from TopClass;
    
    
    Create(S   : in out TheSolidExplorer;
           P   :        Pnt from gp;
	   Tol :        Real from Standard)
    	---Purpose: Constructor to classify the point P with the 
    	--          tolerance Tol on the solid S.
    returns SolidClassifier from TopClass;
    
    
    Perform(me  : in out;
            S   : in out  TheSolidExplorer;
            P   :         Pnt from gp;
	    Tol :         Real from Standard);
    	---Purpose: Classify the point P with the 
    	--          tolerance Tol on the solid S.

    
    Rejected(me)
    	---Purpose: Returns True if the classification has been 
    	--          computed by rejection. 
    	--          The State is then OUT.
    returns Boolean from Standard;
    
    
    State(me)  returns State  from TopAbs;
    	---Purpose: Returns the result of the classification.
    
    IsOnAFace(me) returns Boolean from Standard;
    	---Purpose: Returns True when the point is a point of a face.
    
    Face(me) 
    	---Purpose: Returns the face used to determine the 
    	--          classification. When the state is ON, this is the 
    	--          face containing the point. 
    	--          
    	--          When Rejected() returns True, Face() has no signification.
    returns Face from TopoDS;
    	    
fields

    myFace         : Face       from TopoDS;
    myState        : Integer    from Standard;  -- 1: Rejected     2: IsOnFace  3: In  4: Out
    
end SolidClassifier;
