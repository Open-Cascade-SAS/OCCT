-- Created on: 2009-01-26
-- Created by: Pavel TELKOV
-- Copyright (c) 2009-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PairOfPolygon from BRepMesh 

	---Purpose: 

uses
    PolygonOnTriangulation from Poly

is
    Create
    ---Purpose: Create empty pair with null fileds
    returns PairOfPolygon from BRepMesh;

    Clear(me: out);
    ---Purpose: Clear pair handles
    
    Prepend (me: out; thePoly: PolygonOnTriangulation from Poly);
    --- Initialise first polygon on triangulation
    
    Append (me: out; thePoly: PolygonOnTriangulation from Poly);
    --- Initialise first or last polygon on triangulation
    
    First(me)
    ---Purpose: Returns first polygon on triangulation
    ---C++: return const &
    ---C++: inline
    returns PolygonOnTriangulation from Poly;

    Last(me)
    ---Purpose: Returns last polygon on triangulation
    ---C++: return const &
    ---C++: inline
    returns PolygonOnTriangulation from Poly;

fields
    myFirst : PolygonOnTriangulation from Poly;
    myLast  : PolygonOnTriangulation from Poly;
     
end PairOfPolygon;
