-- Created on: 1995-02-24
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



generic class SurfProps from Contap 
    (TheSurface     as any;
     TheSurfaceTool as any) -- as SurfaceTool from Contap

	---Purpose: Internal tool used  to compute the  normal and its
	--          derivatives. 

uses Pnt from gp,
     Vec from gp

is

    Normale(myclass; S: TheSurface; U,V: Real from Standard;
                     P: out Pnt from gp;
		     N: out Vec from gp);

	---Purpose: Computes  the point <P>, and  normal vector <N> on
	--          <S> at parameters U,V.



    DerivAndNorm(myclass; S: TheSurface; U,V: Real from Standard;
                          P      : out Pnt from gp;
			  d1u,d1v: out Vec from gp;
		          N      : out Vec from gp);

	---Purpose: Computes  the point <P>, and  normal vector <N> on
	--          <S> at parameters U,V.



    NormAndDn(myclass; S: TheSurface; U,V: Real from Standard;
                       P        : out Pnt from gp;
		       N,Dnu,Dnv: out Vec from gp);

	---Purpose: Computes the point <P>, normal vector <N>, and its
	--          derivatives <Dnu> and <Dnv> on <S> at parameters U,V.


end SurfProps;
