-- Created on: 1996-01-26
-- Created by: Christian CAILLET
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SignValidity  from IFSelect  inherits Signature

    ---Purpose : This Signature returns the Validity Status of an entity, as
    --           deducted from data in the model : it can be
    --           "OK" "Unknown" "Unloaded" "Syntactic Fail"(but loaded)
    --           "Syntactic Warning" "Semantic Fail" "Semantic Warning"


uses CString, Transient, InterfaceModel

is

    Create returns SignValidity;
    ---Purpose : Returns a SignValidity

    CVal  (myclass; ent : any Transient; model : InterfaceModel) returns CString;
    ---Purpose : Returns the Signature for a Transient object, as a validity
    --           deducted from data (reports) stored in the model.
    --           Class method, can be called by any one

    Value (me; ent : any Transient; model : InterfaceModel) returns CString;
    ---Purpose : Returns the Signature for a Transient object, as a validity
    --           deducted from data (reports) stored in the model
    --           Calls the class method CVal

end SignValidity;
