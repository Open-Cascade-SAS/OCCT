-- Created on: 1995-05-29
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PntFace from LocOpe

	---Purpose: 

uses Pnt         from gp,
     Face        from TopoDS,
     Orientation from TopAbs
     

is

    Create
	---Purpose: Empty constructor. Useful only for the list.
    	returns PntFace from LocOpe;


    Create (P: Pnt from gp; F: Face from TopoDS;
            Or: Orientation from TopAbs; Param,UPar,VPar: Real from Standard) 
	    
    	returns PntFace from LocOpe;
	---C++: inline

    Pnt(me)
    
    	returns Pnt from gp
	---C++: return const&
	---C++: inline
	is static;


    Face(me)
    
    	returns Face from TopoDS
	---C++: return const&
	---C++: inline
	is static;

    Orientation(me)
    
    	returns Orientation from TopAbs
	---C++: inline
	is static;


    ChangeOrientation(me: in out)
    
    	returns Orientation from TopAbs
	---C++: return &
	---C++: inline
	is static;


    Parameter(me)
    
    	returns Real from Standard
	---C++: inline
	is static;


    UParameter(me)
    
    	returns Real from Standard
	---C++: inline
	is static;


    VParameter(me)
    
    	returns Real from Standard
	---C++: inline
	is static;


fields

    myPnt  : Pnt         from gp;
    myFace : Face        from TopoDS;
    myOri  : Orientation from TopAbs;
    myPar  : Real        from Standard;
    myUPar : Real        from Standard;
    myVPar : Real        from Standard;

end PntFace;
