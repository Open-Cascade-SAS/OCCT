-- Created on: 1998-03-12
-- Created by: Roman LYGIN
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SplitCurve3d from ShapeUpgrade inherits SplitCurve from ShapeUpgrade 

    ---Purpose: Splits a 3d curve with a criterion.
    
uses     
    Curve          from Geom,
    HArray1OfCurve from TColGeom
   
is 
 
    Create returns SplitCurve3d from ShapeUpgrade;
    	---Purpose: Empty constructor.

    Init (me: mutable; C: Curve from  Geom);
       	---Purpose: Initializes with curve with its first and last parameters.
	
    Init (me: mutable; C          : Curve from  Geom;
    	    	       First, Last: Real);
       	---Purpose: Initializes with curve with its parameters.
	
    Build (me: mutable; Segment: Boolean) is redefined;
       ---Purpose: If Segment is True, the result is composed with
       --  segments of the curve bounded by the SplitValues.  If
       --  Segment is False, the result is composed with trimmed
       --  Curves all based on the same complete curve.
       --  
    
    GetCurves(me) returns  HArray1OfCurve  from  TColGeom;
       ---C++: return const &

fields 
 
    myCurve          : Curve  from  Geom is protected;
    myResultingCurves: HArray1OfCurve  from TColGeom is protected;
    
end;
    
