-- Created on: 1997-04-21
-- Created by: Denis PASCAL
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class Dimension from DrawDim inherits Drawable3D from Draw

	---Purpose: 

uses 
    Real       from Standard,
    Pnt        from gp,
    Color      from Draw,
    Display    from Draw

is

    Initialize;

    SetValue (me : mutable; avalue : Real from Standard);
    
    GetValue (me)
    returns Real from Standard;
    
    IsValued (me)
    returns Boolean from Standard;
    
    TextColor(me : mutable; C : Color from Draw);
    
    TextColor(me) returns Color from Draw;
    
    DrawText(me; Pos : Pnt from gp; D : in out Display from Draw);
    
fields

    is_valued     : Boolean from Standard is protected;
    myValue       : Real    from Standard is protected;
    myTextColor   : Color   from Draw     is protected;
    
end Dimension;
