-- Created on: 1991-02-27
-- Created by: Jean Claude Vauthier
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class UniformDeflection from CPnts 
 
        ---Purpose : This class defines an algorithm to create a set of points
        -- (with a given chordal deviation) at the
        --  positions of constant deflection of a given parametrized curve or a trimmed
        --  circle.
        --  The continuity of the curve must be at least C2.
        --
        --  the usage of the is the following.
        --          
        --  class myUniformDFeflection instantiates
        --                     UniformDeflection(Curve, Tool);
        --
        --      
        -- Curve C; // Curve inherits from Curve or Curve2d from Adaptor2d
        -- myUniformDeflection Iter1;
        -- DefPntOfmyUniformDeflection P;
        --        
        -- for(Iter1.Initialize(C, Deflection, EPSILON, True); 
        --     Iter1.More();
        --     Iter1.Next()) {
        --   P = Iter1.Value();
        --   ... make something with P
        -- }
        -- if(!Iter1.IsAllDone()) {
        --    ... something wrong happened 
        -- }
uses
    Curve   from Adaptor3d,
    Curve2d from Adaptor2d,
    Pnt     from gp

raises DomainError from Standard, 
       NotDone     from StdFail, 
       OutOfRange  from Standard

is


        --        
  
  Create 
  ---Purpose: creation of a indefinite UniformDeflection
  returns UniformDeflection;

  Create(C : Curve from Adaptor3d; Deflection,  Resolution  : Real; 
                                 WithControl : Boolean )
        --- Purpose :  Computes a uniform deflection distribution of points
        --  on the curve <C>.
        --  <Deflection> defines the constant deflection value.
        --  The algorithm computes the number of points and the points.
        --  The curve <C> must be at least C2 else the computation can fail.
        --  If just some parts of the curve is C2 it is better to give the 
        --  parameters bounds and to use the below constructor .
        --  if <WithControl> is True, the algorithm controls the estimate 
        --  deflection
        --  when the curve is singular at the point P(u),the algorithm 
        --  computes the next point as  
        --  P(u + Max(CurrentStep,Abs(LastParameter-FirstParameter)))
        --  if the singularity is at the first point ,the next point
        --  calculated is the P(LastParameter)   
     returns UniformDeflection;

  Create(C : Curve2d from Adaptor2d; Deflection,  Resolution  : Real; 
                                   WithControl : Boolean )
	---Purpose: As above with 2d curve
     returns UniformDeflection;

  Create(C : Curve from Adaptor3d; Deflection, U1, U2, Resolution : Real; 
                    WithControl : Boolean)
        --- Purpose :
        --  Computes an uniform deflection distribution of points on a part of
        --  the curve <C>. Deflection defines the step between the points.
        --  <U1> and <U2> define the distribution span. 
        --  <U1> and <U2> must be in the parametric range of the curve.
     returns UniformDeflection
     raises DomainError;
        --  raised if U1 and U2 are not in the parametric bounds of the curve.

  Create(C : Curve2d from Adaptor2d; Deflection, U1, U2, Resolution : Real; 
                    WithControl : Boolean)
        --- Purpose : As above with 2d curve
     returns UniformDeflection
     raises DomainError;
        --  raised if U1 and U2 are not in the parametric bounds of the curve.

    Initialize(me : in out; C : Curve from Adaptor3d; 
                            Deflection, Resolution : Real; 
                            WithControl : Boolean)
    	---Purpose: Initialize the algoritms with <C>, <Deflection>, <UStep>,
    	--          <Resolution> and <WithControl>
        is static;
     
    Initialize(me : in out; C : Curve2d from Adaptor2d; 
                            Deflection, Resolution : Real; 
                            WithControl : Boolean)
    	---Purpose: Initialize the algoritms with <C>, <Deflection>, <UStep>,
    	--          <Resolution> and <WithControl>
        is static;
     
    Initialize(me : in out; C : Curve from Adaptor3d; 
                            Deflection, U1, U2, Resolution : Real; 
                            WithControl : Boolean)
    	---Purpose: Initialize the algoritms with <C>, <Deflection>, <UStep>,
    	--          <U1>, <U2> and <WithControl>
     	raises DomainError
	is static;
  
    Initialize(me : in out; C : Curve2d from Adaptor2d; 
                            Deflection, U1, U2, Resolution : Real; 
                            WithControl : Boolean)
    	---Purpose: Initialize the algoritms with <C>, <Deflection>, <UStep>,
    	--          <U1>, <U2> and <WithControl>
     	raises DomainError
	is static;
  
    IsAllDone (me)
        --- Purpose : To know if all the calculus were done successfully
        --  (ie all the points have been computed). The calculus can fail if
        --  the Curve is not C1 in the considered domain.
        --  Returns True if the calculus was successful.
        ---C++: inline
        returns Boolean
     	is static;

    Next(me : in out)
        ---Purpose: go to the next Point.
        ---C++: inline
    	raises OutOfRange
    	is static;  

    More(me : in out)
        ---Purpose: returns True if it exists a next Point.
    	returns Boolean
      	is static;
  
    Value(me) returns Real
        ---Purpose : return the computed parameter
        ---C++: inline
    	is static;


    Point(me) returns Pnt from gp
        ---Purpose : return the computed parameter
        ---C++: inline
    	is static;
	
    Perform (me : in out)  
        ---Purpose: algorithm 
    	is static private;
	
fields

    myDone       : Boolean;
    my3d         : Boolean;
    myCurve      : Address from Standard;
    myFinish     : Boolean;
    myTolCur     : Real;
    myControl    : Boolean;
    myIPoint     : Integer;
    myNbPoints   : Integer;
    myParams     : Real[3];
    myPoints     : Pnt from gp [3] ;
    myDwmax      : Real;
    myDeflection : Real;
    myFirstParam : Real;
    myLastParam  : Real;
    myDu         : Real;
    
end UniformDeflection;





