-- Created on: 2002-10-29
-- Created by: Michael SAZONOV
-- Copyright (c) 2002-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


deferred class ADriver from BinMDF inherits TShared from MMgt

        ---Purpose: Attribute Storage/Retrieval Driver.

uses
    ExtendedString   from TCollection,
    MessageDriver    from CDM,
    AsciiString      from TCollection,
    Attribute        from TDF,
    RRelocationTable from BinObjMgt,
    SRelocationTable from BinObjMgt,
    Persistent       from BinObjMgt

is
    Initialize (theMsgDriver: MessageDriver from CDM;
                theName     : CString from Standard = NULL);

    NewEmpty    (me)
        returns mutable Attribute from TDF
        is deferred;
        ---Purpose: Creates a new attribute from TDF.

    SourceType  (me) returns Type from Standard;
        ---C++: return const &
	---C++: inline
        ---Purpose: Returns the type of source object,
        --          inheriting from Attribute from TDF.

    TypeName    (me)
        returns AsciiString from TCollection
        is static;
        ---C++: return const &
	---C++: inline
        ---Purpose: Returns the type name of the attribute object

    Paste       (me; aSource     : Persistent from BinObjMgt;
                     aTarget     : mutable Attribute from TDF;
                     aRelocTable : out RRelocationTable from BinObjMgt)
        returns Boolean from Standard is deferred;
        ---Purpose: Translate the contents of <aSource> and put it
        --          into <aTarget>, using the relocation table
        --          <aRelocTable> to keep the sharings.

    Paste       (me; aSource     : Attribute from TDF;
                     aTarget     : in out Persistent from BinObjMgt;
                     aRelocTable : out SRelocationTable from BinObjMgt)
        is deferred;
        ---Purpose: Translate the contents of <aSource> and put it
        --          into <aTarget>, using the relocation table
        --          <aRelocTable> to keep the sharings.

    WriteMessage (me; theMessage : ExtendedString from TCollection);
        ---Purpose: Send message to Application (usually when error occurres)

fields

    myMessageDriver : MessageDriver from CDM;
    myTypeName      : AsciiString   from TCollection is protected;

end ADriver;
